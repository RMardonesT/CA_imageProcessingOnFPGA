`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/10/2022 12:12:04 PM
// Design Name: 
// Module Name: GRID_SCRIPT
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module GRID_SCRIPT
    #(parameter M = 3, N = 3)

    (


    input logic clk, reset,
    
    input logic [2:0] operation,       
    
    input logic [0:0] data_in,
    
    
    
    output logic [0:0] gen [M*N -1 :0] ,
    output logic [7:0] data_out    
        
    );/******************* CELL 0 ***************/  

	CELDA   #(.ic(0), .top_row(1), .load_cell(1))

		cell0 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[96]),
			.N(gen[95]),
			.NE(gen[96]),

			.O(data_in),
			.E(gen[1]),

			.SO(gen[96]),
			.S(gen[95]),
			.SE(gen[96]),

			.SELF(gen[0]),
			.cell_state(gen[0])
		); 

/******************* CELL 1 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell1 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[95]),
			.N(gen[96]),
			.NE(gen[97]),

			.O(gen[0]),
			.E(gen[2]),

			.SO(gen[95]),
			.S(gen[96]),
			.SE(gen[97]),

			.SELF(gen[1]),
			.cell_state(gen[1])
		); 

/******************* CELL 2 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell2 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[96]),
			.N(gen[97]),
			.NE(gen[98]),

			.O(gen[1]),
			.E(gen[3]),

			.SO(gen[96]),
			.S(gen[97]),
			.SE(gen[98]),

			.SELF(gen[2]),
			.cell_state(gen[2])
		); 

/******************* CELL 3 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell3 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[97]),
			.N(gen[98]),
			.NE(gen[99]),

			.O(gen[2]),
			.E(gen[4]),

			.SO(gen[97]),
			.S(gen[98]),
			.SE(gen[99]),

			.SELF(gen[3]),
			.cell_state(gen[3])
		); 

/******************* CELL 4 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell4 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[98]),
			.N(gen[99]),
			.NE(gen[100]),

			.O(gen[3]),
			.E(gen[5]),

			.SO(gen[98]),
			.S(gen[99]),
			.SE(gen[100]),

			.SELF(gen[4]),
			.cell_state(gen[4])
		); 

/******************* CELL 5 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell5 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[99]),
			.N(gen[100]),
			.NE(gen[101]),

			.O(gen[4]),
			.E(gen[6]),

			.SO(gen[99]),
			.S(gen[100]),
			.SE(gen[101]),

			.SELF(gen[5]),
			.cell_state(gen[5])
		); 

/******************* CELL 6 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell6 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[100]),
			.N(gen[101]),
			.NE(gen[102]),

			.O(gen[5]),
			.E(gen[7]),

			.SO(gen[100]),
			.S(gen[101]),
			.SE(gen[102]),

			.SELF(gen[6]),
			.cell_state(gen[6])
		); 

/******************* CELL 7 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell7 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[101]),
			.N(gen[102]),
			.NE(gen[103]),

			.O(gen[6]),
			.E(gen[8]),

			.SO(gen[101]),
			.S(gen[102]),
			.SE(gen[103]),

			.SELF(gen[7]),
			.cell_state(gen[7])
		); 

/******************* CELL 8 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell8 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[102]),
			.N(gen[103]),
			.NE(gen[104]),

			.O(gen[7]),
			.E(gen[9]),

			.SO(gen[102]),
			.S(gen[103]),
			.SE(gen[104]),

			.SELF(gen[8]),
			.cell_state(gen[8])
		); 

/******************* CELL 9 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell9 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[103]),
			.N(gen[104]),
			.NE(gen[105]),

			.O(gen[8]),
			.E(gen[10]),

			.SO(gen[103]),
			.S(gen[104]),
			.SE(gen[105]),

			.SELF(gen[9]),
			.cell_state(gen[9])
		); 

/******************* CELL 10 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell10 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[104]),
			.N(gen[105]),
			.NE(gen[106]),

			.O(gen[9]),
			.E(gen[11]),

			.SO(gen[104]),
			.S(gen[105]),
			.SE(gen[106]),

			.SELF(gen[10]),
			.cell_state(gen[10])
		); 

/******************* CELL 11 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell11 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[105]),
			.N(gen[106]),
			.NE(gen[107]),

			.O(gen[10]),
			.E(gen[12]),

			.SO(gen[105]),
			.S(gen[106]),
			.SE(gen[107]),

			.SELF(gen[11]),
			.cell_state(gen[11])
		); 

/******************* CELL 12 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell12 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[106]),
			.N(gen[107]),
			.NE(gen[108]),

			.O(gen[11]),
			.E(gen[13]),

			.SO(gen[106]),
			.S(gen[107]),
			.SE(gen[108]),

			.SELF(gen[12]),
			.cell_state(gen[12])
		); 

/******************* CELL 13 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell13 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[107]),
			.N(gen[108]),
			.NE(gen[109]),

			.O(gen[12]),
			.E(gen[14]),

			.SO(gen[107]),
			.S(gen[108]),
			.SE(gen[109]),

			.SELF(gen[13]),
			.cell_state(gen[13])
		); 

/******************* CELL 14 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell14 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[108]),
			.N(gen[109]),
			.NE(gen[110]),

			.O(gen[13]),
			.E(gen[15]),

			.SO(gen[108]),
			.S(gen[109]),
			.SE(gen[110]),

			.SELF(gen[14]),
			.cell_state(gen[14])
		); 

/******************* CELL 15 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell15 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[109]),
			.N(gen[110]),
			.NE(gen[111]),

			.O(gen[14]),
			.E(gen[16]),

			.SO(gen[109]),
			.S(gen[110]),
			.SE(gen[111]),

			.SELF(gen[15]),
			.cell_state(gen[15])
		); 

/******************* CELL 16 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell16 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[110]),
			.N(gen[111]),
			.NE(gen[112]),

			.O(gen[15]),
			.E(gen[17]),

			.SO(gen[110]),
			.S(gen[111]),
			.SE(gen[112]),

			.SELF(gen[16]),
			.cell_state(gen[16])
		); 

/******************* CELL 17 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell17 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[111]),
			.N(gen[112]),
			.NE(gen[113]),

			.O(gen[16]),
			.E(gen[18]),

			.SO(gen[111]),
			.S(gen[112]),
			.SE(gen[113]),

			.SELF(gen[17]),
			.cell_state(gen[17])
		); 

/******************* CELL 18 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell18 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[112]),
			.N(gen[113]),
			.NE(gen[114]),

			.O(gen[17]),
			.E(gen[19]),

			.SO(gen[112]),
			.S(gen[113]),
			.SE(gen[114]),

			.SELF(gen[18]),
			.cell_state(gen[18])
		); 

/******************* CELL 19 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell19 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[113]),
			.N(gen[114]),
			.NE(gen[115]),

			.O(gen[18]),
			.E(gen[20]),

			.SO(gen[113]),
			.S(gen[114]),
			.SE(gen[115]),

			.SELF(gen[19]),
			.cell_state(gen[19])
		); 

/******************* CELL 20 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell20 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[114]),
			.N(gen[115]),
			.NE(gen[116]),

			.O(gen[19]),
			.E(gen[21]),

			.SO(gen[114]),
			.S(gen[115]),
			.SE(gen[116]),

			.SELF(gen[20]),
			.cell_state(gen[20])
		); 

/******************* CELL 21 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell21 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[115]),
			.N(gen[116]),
			.NE(gen[117]),

			.O(gen[20]),
			.E(gen[22]),

			.SO(gen[115]),
			.S(gen[116]),
			.SE(gen[117]),

			.SELF(gen[21]),
			.cell_state(gen[21])
		); 

/******************* CELL 22 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell22 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[116]),
			.N(gen[117]),
			.NE(gen[118]),

			.O(gen[21]),
			.E(gen[23]),

			.SO(gen[116]),
			.S(gen[117]),
			.SE(gen[118]),

			.SELF(gen[22]),
			.cell_state(gen[22])
		); 

/******************* CELL 23 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell23 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[117]),
			.N(gen[118]),
			.NE(gen[119]),

			.O(gen[22]),
			.E(gen[24]),

			.SO(gen[117]),
			.S(gen[118]),
			.SE(gen[119]),

			.SELF(gen[23]),
			.cell_state(gen[23])
		); 

/******************* CELL 24 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell24 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[118]),
			.N(gen[119]),
			.NE(gen[120]),

			.O(gen[23]),
			.E(gen[25]),

			.SO(gen[118]),
			.S(gen[119]),
			.SE(gen[120]),

			.SELF(gen[24]),
			.cell_state(gen[24])
		); 

/******************* CELL 25 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell25 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[119]),
			.N(gen[120]),
			.NE(gen[121]),

			.O(gen[24]),
			.E(gen[26]),

			.SO(gen[119]),
			.S(gen[120]),
			.SE(gen[121]),

			.SELF(gen[25]),
			.cell_state(gen[25])
		); 

/******************* CELL 26 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell26 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[120]),
			.N(gen[121]),
			.NE(gen[122]),

			.O(gen[25]),
			.E(gen[27]),

			.SO(gen[120]),
			.S(gen[121]),
			.SE(gen[122]),

			.SELF(gen[26]),
			.cell_state(gen[26])
		); 

/******************* CELL 27 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell27 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[121]),
			.N(gen[122]),
			.NE(gen[123]),

			.O(gen[26]),
			.E(gen[28]),

			.SO(gen[121]),
			.S(gen[122]),
			.SE(gen[123]),

			.SELF(gen[27]),
			.cell_state(gen[27])
		); 

/******************* CELL 28 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell28 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[122]),
			.N(gen[123]),
			.NE(gen[124]),

			.O(gen[27]),
			.E(gen[29]),

			.SO(gen[122]),
			.S(gen[123]),
			.SE(gen[124]),

			.SELF(gen[28]),
			.cell_state(gen[28])
		); 

/******************* CELL 29 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell29 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[123]),
			.N(gen[124]),
			.NE(gen[125]),

			.O(gen[28]),
			.E(gen[30]),

			.SO(gen[123]),
			.S(gen[124]),
			.SE(gen[125]),

			.SELF(gen[29]),
			.cell_state(gen[29])
		); 

/******************* CELL 30 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell30 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[124]),
			.N(gen[125]),
			.NE(gen[126]),

			.O(gen[29]),
			.E(gen[31]),

			.SO(gen[124]),
			.S(gen[125]),
			.SE(gen[126]),

			.SELF(gen[30]),
			.cell_state(gen[30])
		); 

/******************* CELL 31 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell31 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[125]),
			.N(gen[126]),
			.NE(gen[127]),

			.O(gen[30]),
			.E(gen[32]),

			.SO(gen[125]),
			.S(gen[126]),
			.SE(gen[127]),

			.SELF(gen[31]),
			.cell_state(gen[31])
		); 

/******************* CELL 32 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell32 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[126]),
			.N(gen[127]),
			.NE(gen[128]),

			.O(gen[31]),
			.E(gen[33]),

			.SO(gen[126]),
			.S(gen[127]),
			.SE(gen[128]),

			.SELF(gen[32]),
			.cell_state(gen[32])
		); 

/******************* CELL 33 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell33 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[127]),
			.N(gen[128]),
			.NE(gen[129]),

			.O(gen[32]),
			.E(gen[34]),

			.SO(gen[127]),
			.S(gen[128]),
			.SE(gen[129]),

			.SELF(gen[33]),
			.cell_state(gen[33])
		); 

/******************* CELL 34 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell34 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[128]),
			.N(gen[129]),
			.NE(gen[130]),

			.O(gen[33]),
			.E(gen[35]),

			.SO(gen[128]),
			.S(gen[129]),
			.SE(gen[130]),

			.SELF(gen[34]),
			.cell_state(gen[34])
		); 

/******************* CELL 35 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell35 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[129]),
			.N(gen[130]),
			.NE(gen[131]),

			.O(gen[34]),
			.E(gen[36]),

			.SO(gen[129]),
			.S(gen[130]),
			.SE(gen[131]),

			.SELF(gen[35]),
			.cell_state(gen[35])
		); 

/******************* CELL 36 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell36 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[130]),
			.N(gen[131]),
			.NE(gen[132]),

			.O(gen[35]),
			.E(gen[37]),

			.SO(gen[130]),
			.S(gen[131]),
			.SE(gen[132]),

			.SELF(gen[36]),
			.cell_state(gen[36])
		); 

/******************* CELL 37 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell37 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[131]),
			.N(gen[132]),
			.NE(gen[133]),

			.O(gen[36]),
			.E(gen[38]),

			.SO(gen[131]),
			.S(gen[132]),
			.SE(gen[133]),

			.SELF(gen[37]),
			.cell_state(gen[37])
		); 

/******************* CELL 38 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell38 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[132]),
			.N(gen[133]),
			.NE(gen[134]),

			.O(gen[37]),
			.E(gen[39]),

			.SO(gen[132]),
			.S(gen[133]),
			.SE(gen[134]),

			.SELF(gen[38]),
			.cell_state(gen[38])
		); 

/******************* CELL 39 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell39 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[133]),
			.N(gen[134]),
			.NE(gen[135]),

			.O(gen[38]),
			.E(gen[40]),

			.SO(gen[133]),
			.S(gen[134]),
			.SE(gen[135]),

			.SELF(gen[39]),
			.cell_state(gen[39])
		); 

/******************* CELL 40 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell40 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[134]),
			.N(gen[135]),
			.NE(gen[136]),

			.O(gen[39]),
			.E(gen[41]),

			.SO(gen[134]),
			.S(gen[135]),
			.SE(gen[136]),

			.SELF(gen[40]),
			.cell_state(gen[40])
		); 

/******************* CELL 41 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell41 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[135]),
			.N(gen[136]),
			.NE(gen[137]),

			.O(gen[40]),
			.E(gen[42]),

			.SO(gen[135]),
			.S(gen[136]),
			.SE(gen[137]),

			.SELF(gen[41]),
			.cell_state(gen[41])
		); 

/******************* CELL 42 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell42 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[136]),
			.N(gen[137]),
			.NE(gen[138]),

			.O(gen[41]),
			.E(gen[43]),

			.SO(gen[136]),
			.S(gen[137]),
			.SE(gen[138]),

			.SELF(gen[42]),
			.cell_state(gen[42])
		); 

/******************* CELL 43 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell43 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[137]),
			.N(gen[138]),
			.NE(gen[139]),

			.O(gen[42]),
			.E(gen[44]),

			.SO(gen[137]),
			.S(gen[138]),
			.SE(gen[139]),

			.SELF(gen[43]),
			.cell_state(gen[43])
		); 

/******************* CELL 44 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell44 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[138]),
			.N(gen[139]),
			.NE(gen[140]),

			.O(gen[43]),
			.E(gen[45]),

			.SO(gen[138]),
			.S(gen[139]),
			.SE(gen[140]),

			.SELF(gen[44]),
			.cell_state(gen[44])
		); 

/******************* CELL 45 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell45 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[139]),
			.N(gen[140]),
			.NE(gen[141]),

			.O(gen[44]),
			.E(gen[46]),

			.SO(gen[139]),
			.S(gen[140]),
			.SE(gen[141]),

			.SELF(gen[45]),
			.cell_state(gen[45])
		); 

/******************* CELL 46 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell46 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[140]),
			.N(gen[141]),
			.NE(gen[142]),

			.O(gen[45]),
			.E(gen[47]),

			.SO(gen[140]),
			.S(gen[141]),
			.SE(gen[142]),

			.SELF(gen[46]),
			.cell_state(gen[46])
		); 

/******************* CELL 47 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell47 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[141]),
			.N(gen[142]),
			.NE(gen[143]),

			.O(gen[46]),
			.E(gen[48]),

			.SO(gen[141]),
			.S(gen[142]),
			.SE(gen[143]),

			.SELF(gen[47]),
			.cell_state(gen[47])
		); 

/******************* CELL 48 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell48 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[142]),
			.N(gen[143]),
			.NE(gen[144]),

			.O(gen[47]),
			.E(gen[49]),

			.SO(gen[142]),
			.S(gen[143]),
			.SE(gen[144]),

			.SELF(gen[48]),
			.cell_state(gen[48])
		); 

/******************* CELL 49 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell49 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[143]),
			.N(gen[144]),
			.NE(gen[145]),

			.O(gen[48]),
			.E(gen[50]),

			.SO(gen[143]),
			.S(gen[144]),
			.SE(gen[145]),

			.SELF(gen[49]),
			.cell_state(gen[49])
		); 

/******************* CELL 50 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell50 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[144]),
			.N(gen[145]),
			.NE(gen[146]),

			.O(gen[49]),
			.E(gen[51]),

			.SO(gen[144]),
			.S(gen[145]),
			.SE(gen[146]),

			.SELF(gen[50]),
			.cell_state(gen[50])
		); 

/******************* CELL 51 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell51 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[145]),
			.N(gen[146]),
			.NE(gen[147]),

			.O(gen[50]),
			.E(gen[52]),

			.SO(gen[145]),
			.S(gen[146]),
			.SE(gen[147]),

			.SELF(gen[51]),
			.cell_state(gen[51])
		); 

/******************* CELL 52 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell52 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[146]),
			.N(gen[147]),
			.NE(gen[148]),

			.O(gen[51]),
			.E(gen[53]),

			.SO(gen[146]),
			.S(gen[147]),
			.SE(gen[148]),

			.SELF(gen[52]),
			.cell_state(gen[52])
		); 

/******************* CELL 53 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell53 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[147]),
			.N(gen[148]),
			.NE(gen[149]),

			.O(gen[52]),
			.E(gen[54]),

			.SO(gen[147]),
			.S(gen[148]),
			.SE(gen[149]),

			.SELF(gen[53]),
			.cell_state(gen[53])
		); 

/******************* CELL 54 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell54 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[148]),
			.N(gen[149]),
			.NE(gen[150]),

			.O(gen[53]),
			.E(gen[55]),

			.SO(gen[148]),
			.S(gen[149]),
			.SE(gen[150]),

			.SELF(gen[54]),
			.cell_state(gen[54])
		); 

/******************* CELL 55 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell55 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[149]),
			.N(gen[150]),
			.NE(gen[151]),

			.O(gen[54]),
			.E(gen[56]),

			.SO(gen[149]),
			.S(gen[150]),
			.SE(gen[151]),

			.SELF(gen[55]),
			.cell_state(gen[55])
		); 

/******************* CELL 56 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell56 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[150]),
			.N(gen[151]),
			.NE(gen[152]),

			.O(gen[55]),
			.E(gen[57]),

			.SO(gen[150]),
			.S(gen[151]),
			.SE(gen[152]),

			.SELF(gen[56]),
			.cell_state(gen[56])
		); 

/******************* CELL 57 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell57 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[151]),
			.N(gen[152]),
			.NE(gen[153]),

			.O(gen[56]),
			.E(gen[58]),

			.SO(gen[151]),
			.S(gen[152]),
			.SE(gen[153]),

			.SELF(gen[57]),
			.cell_state(gen[57])
		); 

/******************* CELL 58 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell58 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[152]),
			.N(gen[153]),
			.NE(gen[154]),

			.O(gen[57]),
			.E(gen[59]),

			.SO(gen[152]),
			.S(gen[153]),
			.SE(gen[154]),

			.SELF(gen[58]),
			.cell_state(gen[58])
		); 

/******************* CELL 59 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell59 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[153]),
			.N(gen[154]),
			.NE(gen[155]),

			.O(gen[58]),
			.E(gen[60]),

			.SO(gen[153]),
			.S(gen[154]),
			.SE(gen[155]),

			.SELF(gen[59]),
			.cell_state(gen[59])
		); 

/******************* CELL 60 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell60 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[154]),
			.N(gen[155]),
			.NE(gen[156]),

			.O(gen[59]),
			.E(gen[61]),

			.SO(gen[154]),
			.S(gen[155]),
			.SE(gen[156]),

			.SELF(gen[60]),
			.cell_state(gen[60])
		); 

/******************* CELL 61 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell61 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[155]),
			.N(gen[156]),
			.NE(gen[157]),

			.O(gen[60]),
			.E(gen[62]),

			.SO(gen[155]),
			.S(gen[156]),
			.SE(gen[157]),

			.SELF(gen[61]),
			.cell_state(gen[61])
		); 

/******************* CELL 62 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell62 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[156]),
			.N(gen[157]),
			.NE(gen[158]),

			.O(gen[61]),
			.E(gen[63]),

			.SO(gen[156]),
			.S(gen[157]),
			.SE(gen[158]),

			.SELF(gen[62]),
			.cell_state(gen[62])
		); 

/******************* CELL 63 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell63 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[157]),
			.N(gen[158]),
			.NE(gen[159]),

			.O(gen[62]),
			.E(gen[64]),

			.SO(gen[157]),
			.S(gen[158]),
			.SE(gen[159]),

			.SELF(gen[63]),
			.cell_state(gen[63])
		); 

/******************* CELL 64 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell64 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[158]),
			.N(gen[159]),
			.NE(gen[160]),

			.O(gen[63]),
			.E(gen[65]),

			.SO(gen[158]),
			.S(gen[159]),
			.SE(gen[160]),

			.SELF(gen[64]),
			.cell_state(gen[64])
		); 

/******************* CELL 65 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell65 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[159]),
			.N(gen[160]),
			.NE(gen[161]),

			.O(gen[64]),
			.E(gen[66]),

			.SO(gen[159]),
			.S(gen[160]),
			.SE(gen[161]),

			.SELF(gen[65]),
			.cell_state(gen[65])
		); 

/******************* CELL 66 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell66 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[160]),
			.N(gen[161]),
			.NE(gen[162]),

			.O(gen[65]),
			.E(gen[67]),

			.SO(gen[160]),
			.S(gen[161]),
			.SE(gen[162]),

			.SELF(gen[66]),
			.cell_state(gen[66])
		); 

/******************* CELL 67 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell67 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[161]),
			.N(gen[162]),
			.NE(gen[163]),

			.O(gen[66]),
			.E(gen[68]),

			.SO(gen[161]),
			.S(gen[162]),
			.SE(gen[163]),

			.SELF(gen[67]),
			.cell_state(gen[67])
		); 

/******************* CELL 68 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell68 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[162]),
			.N(gen[163]),
			.NE(gen[164]),

			.O(gen[67]),
			.E(gen[69]),

			.SO(gen[162]),
			.S(gen[163]),
			.SE(gen[164]),

			.SELF(gen[68]),
			.cell_state(gen[68])
		); 

/******************* CELL 69 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell69 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[163]),
			.N(gen[164]),
			.NE(gen[165]),

			.O(gen[68]),
			.E(gen[70]),

			.SO(gen[163]),
			.S(gen[164]),
			.SE(gen[165]),

			.SELF(gen[69]),
			.cell_state(gen[69])
		); 

/******************* CELL 70 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell70 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[164]),
			.N(gen[165]),
			.NE(gen[166]),

			.O(gen[69]),
			.E(gen[71]),

			.SO(gen[164]),
			.S(gen[165]),
			.SE(gen[166]),

			.SELF(gen[70]),
			.cell_state(gen[70])
		); 

/******************* CELL 71 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell71 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[165]),
			.N(gen[166]),
			.NE(gen[167]),

			.O(gen[70]),
			.E(gen[72]),

			.SO(gen[165]),
			.S(gen[166]),
			.SE(gen[167]),

			.SELF(gen[71]),
			.cell_state(gen[71])
		); 

/******************* CELL 72 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell72 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[166]),
			.N(gen[167]),
			.NE(gen[168]),

			.O(gen[71]),
			.E(gen[73]),

			.SO(gen[166]),
			.S(gen[167]),
			.SE(gen[168]),

			.SELF(gen[72]),
			.cell_state(gen[72])
		); 

/******************* CELL 73 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell73 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[167]),
			.N(gen[168]),
			.NE(gen[169]),

			.O(gen[72]),
			.E(gen[74]),

			.SO(gen[167]),
			.S(gen[168]),
			.SE(gen[169]),

			.SELF(gen[73]),
			.cell_state(gen[73])
		); 

/******************* CELL 74 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell74 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[168]),
			.N(gen[169]),
			.NE(gen[170]),

			.O(gen[73]),
			.E(gen[75]),

			.SO(gen[168]),
			.S(gen[169]),
			.SE(gen[170]),

			.SELF(gen[74]),
			.cell_state(gen[74])
		); 

/******************* CELL 75 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell75 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[169]),
			.N(gen[170]),
			.NE(gen[171]),

			.O(gen[74]),
			.E(gen[76]),

			.SO(gen[169]),
			.S(gen[170]),
			.SE(gen[171]),

			.SELF(gen[75]),
			.cell_state(gen[75])
		); 

/******************* CELL 76 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell76 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[170]),
			.N(gen[171]),
			.NE(gen[172]),

			.O(gen[75]),
			.E(gen[77]),

			.SO(gen[170]),
			.S(gen[171]),
			.SE(gen[172]),

			.SELF(gen[76]),
			.cell_state(gen[76])
		); 

/******************* CELL 77 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell77 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[171]),
			.N(gen[172]),
			.NE(gen[173]),

			.O(gen[76]),
			.E(gen[78]),

			.SO(gen[171]),
			.S(gen[172]),
			.SE(gen[173]),

			.SELF(gen[77]),
			.cell_state(gen[77])
		); 

/******************* CELL 78 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell78 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[172]),
			.N(gen[173]),
			.NE(gen[174]),

			.O(gen[77]),
			.E(gen[79]),

			.SO(gen[172]),
			.S(gen[173]),
			.SE(gen[174]),

			.SELF(gen[78]),
			.cell_state(gen[78])
		); 

/******************* CELL 79 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell79 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[173]),
			.N(gen[174]),
			.NE(gen[175]),

			.O(gen[78]),
			.E(gen[80]),

			.SO(gen[173]),
			.S(gen[174]),
			.SE(gen[175]),

			.SELF(gen[79]),
			.cell_state(gen[79])
		); 

/******************* CELL 80 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell80 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[174]),
			.N(gen[175]),
			.NE(gen[176]),

			.O(gen[79]),
			.E(gen[81]),

			.SO(gen[174]),
			.S(gen[175]),
			.SE(gen[176]),

			.SELF(gen[80]),
			.cell_state(gen[80])
		); 

/******************* CELL 81 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell81 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[175]),
			.N(gen[176]),
			.NE(gen[177]),

			.O(gen[80]),
			.E(gen[82]),

			.SO(gen[175]),
			.S(gen[176]),
			.SE(gen[177]),

			.SELF(gen[81]),
			.cell_state(gen[81])
		); 

/******************* CELL 82 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell82 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[176]),
			.N(gen[177]),
			.NE(gen[178]),

			.O(gen[81]),
			.E(gen[83]),

			.SO(gen[176]),
			.S(gen[177]),
			.SE(gen[178]),

			.SELF(gen[82]),
			.cell_state(gen[82])
		); 

/******************* CELL 83 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell83 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[177]),
			.N(gen[178]),
			.NE(gen[179]),

			.O(gen[82]),
			.E(gen[84]),

			.SO(gen[177]),
			.S(gen[178]),
			.SE(gen[179]),

			.SELF(gen[83]),
			.cell_state(gen[83])
		); 

/******************* CELL 84 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell84 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[178]),
			.N(gen[179]),
			.NE(gen[180]),

			.O(gen[83]),
			.E(gen[85]),

			.SO(gen[178]),
			.S(gen[179]),
			.SE(gen[180]),

			.SELF(gen[84]),
			.cell_state(gen[84])
		); 

/******************* CELL 85 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell85 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[179]),
			.N(gen[180]),
			.NE(gen[181]),

			.O(gen[84]),
			.E(gen[86]),

			.SO(gen[179]),
			.S(gen[180]),
			.SE(gen[181]),

			.SELF(gen[85]),
			.cell_state(gen[85])
		); 

/******************* CELL 86 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell86 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[180]),
			.N(gen[181]),
			.NE(gen[182]),

			.O(gen[85]),
			.E(gen[87]),

			.SO(gen[180]),
			.S(gen[181]),
			.SE(gen[182]),

			.SELF(gen[86]),
			.cell_state(gen[86])
		); 

/******************* CELL 87 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell87 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[181]),
			.N(gen[182]),
			.NE(gen[183]),

			.O(gen[86]),
			.E(gen[88]),

			.SO(gen[181]),
			.S(gen[182]),
			.SE(gen[183]),

			.SELF(gen[87]),
			.cell_state(gen[87])
		); 

/******************* CELL 88 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell88 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[182]),
			.N(gen[183]),
			.NE(gen[184]),

			.O(gen[87]),
			.E(gen[89]),

			.SO(gen[182]),
			.S(gen[183]),
			.SE(gen[184]),

			.SELF(gen[88]),
			.cell_state(gen[88])
		); 

/******************* CELL 89 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell89 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[183]),
			.N(gen[184]),
			.NE(gen[185]),

			.O(gen[88]),
			.E(gen[90]),

			.SO(gen[183]),
			.S(gen[184]),
			.SE(gen[185]),

			.SELF(gen[89]),
			.cell_state(gen[89])
		); 

/******************* CELL 90 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell90 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[184]),
			.N(gen[185]),
			.NE(gen[186]),

			.O(gen[89]),
			.E(gen[91]),

			.SO(gen[184]),
			.S(gen[185]),
			.SE(gen[186]),

			.SELF(gen[90]),
			.cell_state(gen[90])
		); 

/******************* CELL 91 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell91 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[185]),
			.N(gen[186]),
			.NE(gen[187]),

			.O(gen[90]),
			.E(gen[92]),

			.SO(gen[185]),
			.S(gen[186]),
			.SE(gen[187]),

			.SELF(gen[91]),
			.cell_state(gen[91])
		); 

/******************* CELL 92 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell92 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[186]),
			.N(gen[187]),
			.NE(gen[188]),

			.O(gen[91]),
			.E(gen[93]),

			.SO(gen[186]),
			.S(gen[187]),
			.SE(gen[188]),

			.SELF(gen[92]),
			.cell_state(gen[92])
		); 

/******************* CELL 93 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell93 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[187]),
			.N(gen[188]),
			.NE(gen[189]),

			.O(gen[92]),
			.E(gen[94]),

			.SO(gen[187]),
			.S(gen[188]),
			.SE(gen[189]),

			.SELF(gen[93]),
			.cell_state(gen[93])
		); 

/******************* CELL 94 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell94 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[188]),
			.N(gen[189]),
			.NE(gen[188]),

			.O(gen[93]),
			.E(gen[93]),

			.SO(gen[188]),
			.S(gen[189]),
			.SE(gen[188]),

			.SELF(gen[94]),
			.cell_state(gen[94])
		); 

/******************* CELL 95 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell95 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1]),
			.N(gen[0]),
			.NE(gen[1]),

			.O(gen[96]),
			.E(gen[96]),

			.SO(gen[191]),
			.S(gen[190]),
			.SE(gen[191]),

			.SELF(gen[95]),
			.cell_state(gen[95])
		); 

/******************* CELL 96 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell96 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[0]),
			.N(gen[1]),
			.NE(gen[2]),

			.O(gen[95]),
			.E(gen[97]),

			.SO(gen[190]),
			.S(gen[191]),
			.SE(gen[192]),

			.SELF(gen[96]),
			.cell_state(gen[96])
		); 

/******************* CELL 97 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell97 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1]),
			.N(gen[2]),
			.NE(gen[3]),

			.O(gen[96]),
			.E(gen[98]),

			.SO(gen[191]),
			.S(gen[192]),
			.SE(gen[193]),

			.SELF(gen[97]),
			.cell_state(gen[97])
		); 

/******************* CELL 98 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell98 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2]),
			.N(gen[3]),
			.NE(gen[4]),

			.O(gen[97]),
			.E(gen[99]),

			.SO(gen[192]),
			.S(gen[193]),
			.SE(gen[194]),

			.SELF(gen[98]),
			.cell_state(gen[98])
		); 

/******************* CELL 99 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell99 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3]),
			.N(gen[4]),
			.NE(gen[5]),

			.O(gen[98]),
			.E(gen[100]),

			.SO(gen[193]),
			.S(gen[194]),
			.SE(gen[195]),

			.SELF(gen[99]),
			.cell_state(gen[99])
		); 

/******************* CELL 100 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell100 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4]),
			.N(gen[5]),
			.NE(gen[6]),

			.O(gen[99]),
			.E(gen[101]),

			.SO(gen[194]),
			.S(gen[195]),
			.SE(gen[196]),

			.SELF(gen[100]),
			.cell_state(gen[100])
		); 

/******************* CELL 101 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell101 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5]),
			.N(gen[6]),
			.NE(gen[7]),

			.O(gen[100]),
			.E(gen[102]),

			.SO(gen[195]),
			.S(gen[196]),
			.SE(gen[197]),

			.SELF(gen[101]),
			.cell_state(gen[101])
		); 

/******************* CELL 102 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell102 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6]),
			.N(gen[7]),
			.NE(gen[8]),

			.O(gen[101]),
			.E(gen[103]),

			.SO(gen[196]),
			.S(gen[197]),
			.SE(gen[198]),

			.SELF(gen[102]),
			.cell_state(gen[102])
		); 

/******************* CELL 103 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell103 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7]),
			.N(gen[8]),
			.NE(gen[9]),

			.O(gen[102]),
			.E(gen[104]),

			.SO(gen[197]),
			.S(gen[198]),
			.SE(gen[199]),

			.SELF(gen[103]),
			.cell_state(gen[103])
		); 

/******************* CELL 104 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell104 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8]),
			.N(gen[9]),
			.NE(gen[10]),

			.O(gen[103]),
			.E(gen[105]),

			.SO(gen[198]),
			.S(gen[199]),
			.SE(gen[200]),

			.SELF(gen[104]),
			.cell_state(gen[104])
		); 

/******************* CELL 105 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell105 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[9]),
			.N(gen[10]),
			.NE(gen[11]),

			.O(gen[104]),
			.E(gen[106]),

			.SO(gen[199]),
			.S(gen[200]),
			.SE(gen[201]),

			.SELF(gen[105]),
			.cell_state(gen[105])
		); 

/******************* CELL 106 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell106 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[10]),
			.N(gen[11]),
			.NE(gen[12]),

			.O(gen[105]),
			.E(gen[107]),

			.SO(gen[200]),
			.S(gen[201]),
			.SE(gen[202]),

			.SELF(gen[106]),
			.cell_state(gen[106])
		); 

/******************* CELL 107 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell107 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[11]),
			.N(gen[12]),
			.NE(gen[13]),

			.O(gen[106]),
			.E(gen[108]),

			.SO(gen[201]),
			.S(gen[202]),
			.SE(gen[203]),

			.SELF(gen[107]),
			.cell_state(gen[107])
		); 

/******************* CELL 108 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell108 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[12]),
			.N(gen[13]),
			.NE(gen[14]),

			.O(gen[107]),
			.E(gen[109]),

			.SO(gen[202]),
			.S(gen[203]),
			.SE(gen[204]),

			.SELF(gen[108]),
			.cell_state(gen[108])
		); 

/******************* CELL 109 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell109 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[13]),
			.N(gen[14]),
			.NE(gen[15]),

			.O(gen[108]),
			.E(gen[110]),

			.SO(gen[203]),
			.S(gen[204]),
			.SE(gen[205]),

			.SELF(gen[109]),
			.cell_state(gen[109])
		); 

/******************* CELL 110 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell110 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[14]),
			.N(gen[15]),
			.NE(gen[16]),

			.O(gen[109]),
			.E(gen[111]),

			.SO(gen[204]),
			.S(gen[205]),
			.SE(gen[206]),

			.SELF(gen[110]),
			.cell_state(gen[110])
		); 

/******************* CELL 111 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell111 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[15]),
			.N(gen[16]),
			.NE(gen[17]),

			.O(gen[110]),
			.E(gen[112]),

			.SO(gen[205]),
			.S(gen[206]),
			.SE(gen[207]),

			.SELF(gen[111]),
			.cell_state(gen[111])
		); 

/******************* CELL 112 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell112 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[16]),
			.N(gen[17]),
			.NE(gen[18]),

			.O(gen[111]),
			.E(gen[113]),

			.SO(gen[206]),
			.S(gen[207]),
			.SE(gen[208]),

			.SELF(gen[112]),
			.cell_state(gen[112])
		); 

/******************* CELL 113 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell113 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[17]),
			.N(gen[18]),
			.NE(gen[19]),

			.O(gen[112]),
			.E(gen[114]),

			.SO(gen[207]),
			.S(gen[208]),
			.SE(gen[209]),

			.SELF(gen[113]),
			.cell_state(gen[113])
		); 

/******************* CELL 114 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell114 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[18]),
			.N(gen[19]),
			.NE(gen[20]),

			.O(gen[113]),
			.E(gen[115]),

			.SO(gen[208]),
			.S(gen[209]),
			.SE(gen[210]),

			.SELF(gen[114]),
			.cell_state(gen[114])
		); 

/******************* CELL 115 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell115 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[19]),
			.N(gen[20]),
			.NE(gen[21]),

			.O(gen[114]),
			.E(gen[116]),

			.SO(gen[209]),
			.S(gen[210]),
			.SE(gen[211]),

			.SELF(gen[115]),
			.cell_state(gen[115])
		); 

/******************* CELL 116 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell116 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[20]),
			.N(gen[21]),
			.NE(gen[22]),

			.O(gen[115]),
			.E(gen[117]),

			.SO(gen[210]),
			.S(gen[211]),
			.SE(gen[212]),

			.SELF(gen[116]),
			.cell_state(gen[116])
		); 

/******************* CELL 117 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell117 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[21]),
			.N(gen[22]),
			.NE(gen[23]),

			.O(gen[116]),
			.E(gen[118]),

			.SO(gen[211]),
			.S(gen[212]),
			.SE(gen[213]),

			.SELF(gen[117]),
			.cell_state(gen[117])
		); 

/******************* CELL 118 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell118 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[22]),
			.N(gen[23]),
			.NE(gen[24]),

			.O(gen[117]),
			.E(gen[119]),

			.SO(gen[212]),
			.S(gen[213]),
			.SE(gen[214]),

			.SELF(gen[118]),
			.cell_state(gen[118])
		); 

/******************* CELL 119 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell119 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[23]),
			.N(gen[24]),
			.NE(gen[25]),

			.O(gen[118]),
			.E(gen[120]),

			.SO(gen[213]),
			.S(gen[214]),
			.SE(gen[215]),

			.SELF(gen[119]),
			.cell_state(gen[119])
		); 

/******************* CELL 120 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell120 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[24]),
			.N(gen[25]),
			.NE(gen[26]),

			.O(gen[119]),
			.E(gen[121]),

			.SO(gen[214]),
			.S(gen[215]),
			.SE(gen[216]),

			.SELF(gen[120]),
			.cell_state(gen[120])
		); 

/******************* CELL 121 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell121 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[25]),
			.N(gen[26]),
			.NE(gen[27]),

			.O(gen[120]),
			.E(gen[122]),

			.SO(gen[215]),
			.S(gen[216]),
			.SE(gen[217]),

			.SELF(gen[121]),
			.cell_state(gen[121])
		); 

/******************* CELL 122 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell122 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[26]),
			.N(gen[27]),
			.NE(gen[28]),

			.O(gen[121]),
			.E(gen[123]),

			.SO(gen[216]),
			.S(gen[217]),
			.SE(gen[218]),

			.SELF(gen[122]),
			.cell_state(gen[122])
		); 

/******************* CELL 123 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell123 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[27]),
			.N(gen[28]),
			.NE(gen[29]),

			.O(gen[122]),
			.E(gen[124]),

			.SO(gen[217]),
			.S(gen[218]),
			.SE(gen[219]),

			.SELF(gen[123]),
			.cell_state(gen[123])
		); 

/******************* CELL 124 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell124 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[28]),
			.N(gen[29]),
			.NE(gen[30]),

			.O(gen[123]),
			.E(gen[125]),

			.SO(gen[218]),
			.S(gen[219]),
			.SE(gen[220]),

			.SELF(gen[124]),
			.cell_state(gen[124])
		); 

/******************* CELL 125 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell125 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[29]),
			.N(gen[30]),
			.NE(gen[31]),

			.O(gen[124]),
			.E(gen[126]),

			.SO(gen[219]),
			.S(gen[220]),
			.SE(gen[221]),

			.SELF(gen[125]),
			.cell_state(gen[125])
		); 

/******************* CELL 126 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell126 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[30]),
			.N(gen[31]),
			.NE(gen[32]),

			.O(gen[125]),
			.E(gen[127]),

			.SO(gen[220]),
			.S(gen[221]),
			.SE(gen[222]),

			.SELF(gen[126]),
			.cell_state(gen[126])
		); 

/******************* CELL 127 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell127 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[31]),
			.N(gen[32]),
			.NE(gen[33]),

			.O(gen[126]),
			.E(gen[128]),

			.SO(gen[221]),
			.S(gen[222]),
			.SE(gen[223]),

			.SELF(gen[127]),
			.cell_state(gen[127])
		); 

/******************* CELL 128 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell128 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[32]),
			.N(gen[33]),
			.NE(gen[34]),

			.O(gen[127]),
			.E(gen[129]),

			.SO(gen[222]),
			.S(gen[223]),
			.SE(gen[224]),

			.SELF(gen[128]),
			.cell_state(gen[128])
		); 

/******************* CELL 129 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell129 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[33]),
			.N(gen[34]),
			.NE(gen[35]),

			.O(gen[128]),
			.E(gen[130]),

			.SO(gen[223]),
			.S(gen[224]),
			.SE(gen[225]),

			.SELF(gen[129]),
			.cell_state(gen[129])
		); 

/******************* CELL 130 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell130 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[34]),
			.N(gen[35]),
			.NE(gen[36]),

			.O(gen[129]),
			.E(gen[131]),

			.SO(gen[224]),
			.S(gen[225]),
			.SE(gen[226]),

			.SELF(gen[130]),
			.cell_state(gen[130])
		); 

/******************* CELL 131 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell131 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[35]),
			.N(gen[36]),
			.NE(gen[37]),

			.O(gen[130]),
			.E(gen[132]),

			.SO(gen[225]),
			.S(gen[226]),
			.SE(gen[227]),

			.SELF(gen[131]),
			.cell_state(gen[131])
		); 

/******************* CELL 132 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell132 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[36]),
			.N(gen[37]),
			.NE(gen[38]),

			.O(gen[131]),
			.E(gen[133]),

			.SO(gen[226]),
			.S(gen[227]),
			.SE(gen[228]),

			.SELF(gen[132]),
			.cell_state(gen[132])
		); 

/******************* CELL 133 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell133 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[37]),
			.N(gen[38]),
			.NE(gen[39]),

			.O(gen[132]),
			.E(gen[134]),

			.SO(gen[227]),
			.S(gen[228]),
			.SE(gen[229]),

			.SELF(gen[133]),
			.cell_state(gen[133])
		); 

/******************* CELL 134 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell134 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[38]),
			.N(gen[39]),
			.NE(gen[40]),

			.O(gen[133]),
			.E(gen[135]),

			.SO(gen[228]),
			.S(gen[229]),
			.SE(gen[230]),

			.SELF(gen[134]),
			.cell_state(gen[134])
		); 

/******************* CELL 135 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell135 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[39]),
			.N(gen[40]),
			.NE(gen[41]),

			.O(gen[134]),
			.E(gen[136]),

			.SO(gen[229]),
			.S(gen[230]),
			.SE(gen[231]),

			.SELF(gen[135]),
			.cell_state(gen[135])
		); 

/******************* CELL 136 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell136 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[40]),
			.N(gen[41]),
			.NE(gen[42]),

			.O(gen[135]),
			.E(gen[137]),

			.SO(gen[230]),
			.S(gen[231]),
			.SE(gen[232]),

			.SELF(gen[136]),
			.cell_state(gen[136])
		); 

/******************* CELL 137 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell137 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[41]),
			.N(gen[42]),
			.NE(gen[43]),

			.O(gen[136]),
			.E(gen[138]),

			.SO(gen[231]),
			.S(gen[232]),
			.SE(gen[233]),

			.SELF(gen[137]),
			.cell_state(gen[137])
		); 

/******************* CELL 138 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell138 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[42]),
			.N(gen[43]),
			.NE(gen[44]),

			.O(gen[137]),
			.E(gen[139]),

			.SO(gen[232]),
			.S(gen[233]),
			.SE(gen[234]),

			.SELF(gen[138]),
			.cell_state(gen[138])
		); 

/******************* CELL 139 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell139 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[43]),
			.N(gen[44]),
			.NE(gen[45]),

			.O(gen[138]),
			.E(gen[140]),

			.SO(gen[233]),
			.S(gen[234]),
			.SE(gen[235]),

			.SELF(gen[139]),
			.cell_state(gen[139])
		); 

/******************* CELL 140 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell140 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[44]),
			.N(gen[45]),
			.NE(gen[46]),

			.O(gen[139]),
			.E(gen[141]),

			.SO(gen[234]),
			.S(gen[235]),
			.SE(gen[236]),

			.SELF(gen[140]),
			.cell_state(gen[140])
		); 

/******************* CELL 141 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell141 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[45]),
			.N(gen[46]),
			.NE(gen[47]),

			.O(gen[140]),
			.E(gen[142]),

			.SO(gen[235]),
			.S(gen[236]),
			.SE(gen[237]),

			.SELF(gen[141]),
			.cell_state(gen[141])
		); 

/******************* CELL 142 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell142 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[46]),
			.N(gen[47]),
			.NE(gen[48]),

			.O(gen[141]),
			.E(gen[143]),

			.SO(gen[236]),
			.S(gen[237]),
			.SE(gen[238]),

			.SELF(gen[142]),
			.cell_state(gen[142])
		); 

/******************* CELL 143 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell143 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[47]),
			.N(gen[48]),
			.NE(gen[49]),

			.O(gen[142]),
			.E(gen[144]),

			.SO(gen[237]),
			.S(gen[238]),
			.SE(gen[239]),

			.SELF(gen[143]),
			.cell_state(gen[143])
		); 

/******************* CELL 144 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell144 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[48]),
			.N(gen[49]),
			.NE(gen[50]),

			.O(gen[143]),
			.E(gen[145]),

			.SO(gen[238]),
			.S(gen[239]),
			.SE(gen[240]),

			.SELF(gen[144]),
			.cell_state(gen[144])
		); 

/******************* CELL 145 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell145 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[49]),
			.N(gen[50]),
			.NE(gen[51]),

			.O(gen[144]),
			.E(gen[146]),

			.SO(gen[239]),
			.S(gen[240]),
			.SE(gen[241]),

			.SELF(gen[145]),
			.cell_state(gen[145])
		); 

/******************* CELL 146 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell146 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[50]),
			.N(gen[51]),
			.NE(gen[52]),

			.O(gen[145]),
			.E(gen[147]),

			.SO(gen[240]),
			.S(gen[241]),
			.SE(gen[242]),

			.SELF(gen[146]),
			.cell_state(gen[146])
		); 

/******************* CELL 147 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell147 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[51]),
			.N(gen[52]),
			.NE(gen[53]),

			.O(gen[146]),
			.E(gen[148]),

			.SO(gen[241]),
			.S(gen[242]),
			.SE(gen[243]),

			.SELF(gen[147]),
			.cell_state(gen[147])
		); 

/******************* CELL 148 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell148 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[52]),
			.N(gen[53]),
			.NE(gen[54]),

			.O(gen[147]),
			.E(gen[149]),

			.SO(gen[242]),
			.S(gen[243]),
			.SE(gen[244]),

			.SELF(gen[148]),
			.cell_state(gen[148])
		); 

/******************* CELL 149 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell149 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[53]),
			.N(gen[54]),
			.NE(gen[55]),

			.O(gen[148]),
			.E(gen[150]),

			.SO(gen[243]),
			.S(gen[244]),
			.SE(gen[245]),

			.SELF(gen[149]),
			.cell_state(gen[149])
		); 

/******************* CELL 150 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell150 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[54]),
			.N(gen[55]),
			.NE(gen[56]),

			.O(gen[149]),
			.E(gen[151]),

			.SO(gen[244]),
			.S(gen[245]),
			.SE(gen[246]),

			.SELF(gen[150]),
			.cell_state(gen[150])
		); 

/******************* CELL 151 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell151 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[55]),
			.N(gen[56]),
			.NE(gen[57]),

			.O(gen[150]),
			.E(gen[152]),

			.SO(gen[245]),
			.S(gen[246]),
			.SE(gen[247]),

			.SELF(gen[151]),
			.cell_state(gen[151])
		); 

/******************* CELL 152 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell152 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[56]),
			.N(gen[57]),
			.NE(gen[58]),

			.O(gen[151]),
			.E(gen[153]),

			.SO(gen[246]),
			.S(gen[247]),
			.SE(gen[248]),

			.SELF(gen[152]),
			.cell_state(gen[152])
		); 

/******************* CELL 153 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell153 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[57]),
			.N(gen[58]),
			.NE(gen[59]),

			.O(gen[152]),
			.E(gen[154]),

			.SO(gen[247]),
			.S(gen[248]),
			.SE(gen[249]),

			.SELF(gen[153]),
			.cell_state(gen[153])
		); 

/******************* CELL 154 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell154 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[58]),
			.N(gen[59]),
			.NE(gen[60]),

			.O(gen[153]),
			.E(gen[155]),

			.SO(gen[248]),
			.S(gen[249]),
			.SE(gen[250]),

			.SELF(gen[154]),
			.cell_state(gen[154])
		); 

/******************* CELL 155 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell155 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[59]),
			.N(gen[60]),
			.NE(gen[61]),

			.O(gen[154]),
			.E(gen[156]),

			.SO(gen[249]),
			.S(gen[250]),
			.SE(gen[251]),

			.SELF(gen[155]),
			.cell_state(gen[155])
		); 

/******************* CELL 156 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell156 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[60]),
			.N(gen[61]),
			.NE(gen[62]),

			.O(gen[155]),
			.E(gen[157]),

			.SO(gen[250]),
			.S(gen[251]),
			.SE(gen[252]),

			.SELF(gen[156]),
			.cell_state(gen[156])
		); 

/******************* CELL 157 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell157 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[61]),
			.N(gen[62]),
			.NE(gen[63]),

			.O(gen[156]),
			.E(gen[158]),

			.SO(gen[251]),
			.S(gen[252]),
			.SE(gen[253]),

			.SELF(gen[157]),
			.cell_state(gen[157])
		); 

/******************* CELL 158 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell158 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[62]),
			.N(gen[63]),
			.NE(gen[64]),

			.O(gen[157]),
			.E(gen[159]),

			.SO(gen[252]),
			.S(gen[253]),
			.SE(gen[254]),

			.SELF(gen[158]),
			.cell_state(gen[158])
		); 

/******************* CELL 159 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell159 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[63]),
			.N(gen[64]),
			.NE(gen[65]),

			.O(gen[158]),
			.E(gen[160]),

			.SO(gen[253]),
			.S(gen[254]),
			.SE(gen[255]),

			.SELF(gen[159]),
			.cell_state(gen[159])
		); 

/******************* CELL 160 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell160 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[64]),
			.N(gen[65]),
			.NE(gen[66]),

			.O(gen[159]),
			.E(gen[161]),

			.SO(gen[254]),
			.S(gen[255]),
			.SE(gen[256]),

			.SELF(gen[160]),
			.cell_state(gen[160])
		); 

/******************* CELL 161 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell161 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[65]),
			.N(gen[66]),
			.NE(gen[67]),

			.O(gen[160]),
			.E(gen[162]),

			.SO(gen[255]),
			.S(gen[256]),
			.SE(gen[257]),

			.SELF(gen[161]),
			.cell_state(gen[161])
		); 

/******************* CELL 162 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell162 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[66]),
			.N(gen[67]),
			.NE(gen[68]),

			.O(gen[161]),
			.E(gen[163]),

			.SO(gen[256]),
			.S(gen[257]),
			.SE(gen[258]),

			.SELF(gen[162]),
			.cell_state(gen[162])
		); 

/******************* CELL 163 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell163 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[67]),
			.N(gen[68]),
			.NE(gen[69]),

			.O(gen[162]),
			.E(gen[164]),

			.SO(gen[257]),
			.S(gen[258]),
			.SE(gen[259]),

			.SELF(gen[163]),
			.cell_state(gen[163])
		); 

/******************* CELL 164 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell164 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[68]),
			.N(gen[69]),
			.NE(gen[70]),

			.O(gen[163]),
			.E(gen[165]),

			.SO(gen[258]),
			.S(gen[259]),
			.SE(gen[260]),

			.SELF(gen[164]),
			.cell_state(gen[164])
		); 

/******************* CELL 165 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell165 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[69]),
			.N(gen[70]),
			.NE(gen[71]),

			.O(gen[164]),
			.E(gen[166]),

			.SO(gen[259]),
			.S(gen[260]),
			.SE(gen[261]),

			.SELF(gen[165]),
			.cell_state(gen[165])
		); 

/******************* CELL 166 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell166 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[70]),
			.N(gen[71]),
			.NE(gen[72]),

			.O(gen[165]),
			.E(gen[167]),

			.SO(gen[260]),
			.S(gen[261]),
			.SE(gen[262]),

			.SELF(gen[166]),
			.cell_state(gen[166])
		); 

/******************* CELL 167 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell167 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[71]),
			.N(gen[72]),
			.NE(gen[73]),

			.O(gen[166]),
			.E(gen[168]),

			.SO(gen[261]),
			.S(gen[262]),
			.SE(gen[263]),

			.SELF(gen[167]),
			.cell_state(gen[167])
		); 

/******************* CELL 168 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell168 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[72]),
			.N(gen[73]),
			.NE(gen[74]),

			.O(gen[167]),
			.E(gen[169]),

			.SO(gen[262]),
			.S(gen[263]),
			.SE(gen[264]),

			.SELF(gen[168]),
			.cell_state(gen[168])
		); 

/******************* CELL 169 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell169 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[73]),
			.N(gen[74]),
			.NE(gen[75]),

			.O(gen[168]),
			.E(gen[170]),

			.SO(gen[263]),
			.S(gen[264]),
			.SE(gen[265]),

			.SELF(gen[169]),
			.cell_state(gen[169])
		); 

/******************* CELL 170 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell170 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[74]),
			.N(gen[75]),
			.NE(gen[76]),

			.O(gen[169]),
			.E(gen[171]),

			.SO(gen[264]),
			.S(gen[265]),
			.SE(gen[266]),

			.SELF(gen[170]),
			.cell_state(gen[170])
		); 

/******************* CELL 171 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell171 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[75]),
			.N(gen[76]),
			.NE(gen[77]),

			.O(gen[170]),
			.E(gen[172]),

			.SO(gen[265]),
			.S(gen[266]),
			.SE(gen[267]),

			.SELF(gen[171]),
			.cell_state(gen[171])
		); 

/******************* CELL 172 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell172 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[76]),
			.N(gen[77]),
			.NE(gen[78]),

			.O(gen[171]),
			.E(gen[173]),

			.SO(gen[266]),
			.S(gen[267]),
			.SE(gen[268]),

			.SELF(gen[172]),
			.cell_state(gen[172])
		); 

/******************* CELL 173 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell173 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[77]),
			.N(gen[78]),
			.NE(gen[79]),

			.O(gen[172]),
			.E(gen[174]),

			.SO(gen[267]),
			.S(gen[268]),
			.SE(gen[269]),

			.SELF(gen[173]),
			.cell_state(gen[173])
		); 

/******************* CELL 174 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell174 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[78]),
			.N(gen[79]),
			.NE(gen[80]),

			.O(gen[173]),
			.E(gen[175]),

			.SO(gen[268]),
			.S(gen[269]),
			.SE(gen[270]),

			.SELF(gen[174]),
			.cell_state(gen[174])
		); 

/******************* CELL 175 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell175 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[79]),
			.N(gen[80]),
			.NE(gen[81]),

			.O(gen[174]),
			.E(gen[176]),

			.SO(gen[269]),
			.S(gen[270]),
			.SE(gen[271]),

			.SELF(gen[175]),
			.cell_state(gen[175])
		); 

/******************* CELL 176 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell176 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[80]),
			.N(gen[81]),
			.NE(gen[82]),

			.O(gen[175]),
			.E(gen[177]),

			.SO(gen[270]),
			.S(gen[271]),
			.SE(gen[272]),

			.SELF(gen[176]),
			.cell_state(gen[176])
		); 

/******************* CELL 177 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell177 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[81]),
			.N(gen[82]),
			.NE(gen[83]),

			.O(gen[176]),
			.E(gen[178]),

			.SO(gen[271]),
			.S(gen[272]),
			.SE(gen[273]),

			.SELF(gen[177]),
			.cell_state(gen[177])
		); 

/******************* CELL 178 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell178 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[82]),
			.N(gen[83]),
			.NE(gen[84]),

			.O(gen[177]),
			.E(gen[179]),

			.SO(gen[272]),
			.S(gen[273]),
			.SE(gen[274]),

			.SELF(gen[178]),
			.cell_state(gen[178])
		); 

/******************* CELL 179 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell179 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[83]),
			.N(gen[84]),
			.NE(gen[85]),

			.O(gen[178]),
			.E(gen[180]),

			.SO(gen[273]),
			.S(gen[274]),
			.SE(gen[275]),

			.SELF(gen[179]),
			.cell_state(gen[179])
		); 

/******************* CELL 180 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell180 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[84]),
			.N(gen[85]),
			.NE(gen[86]),

			.O(gen[179]),
			.E(gen[181]),

			.SO(gen[274]),
			.S(gen[275]),
			.SE(gen[276]),

			.SELF(gen[180]),
			.cell_state(gen[180])
		); 

/******************* CELL 181 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell181 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[85]),
			.N(gen[86]),
			.NE(gen[87]),

			.O(gen[180]),
			.E(gen[182]),

			.SO(gen[275]),
			.S(gen[276]),
			.SE(gen[277]),

			.SELF(gen[181]),
			.cell_state(gen[181])
		); 

/******************* CELL 182 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell182 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[86]),
			.N(gen[87]),
			.NE(gen[88]),

			.O(gen[181]),
			.E(gen[183]),

			.SO(gen[276]),
			.S(gen[277]),
			.SE(gen[278]),

			.SELF(gen[182]),
			.cell_state(gen[182])
		); 

/******************* CELL 183 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell183 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[87]),
			.N(gen[88]),
			.NE(gen[89]),

			.O(gen[182]),
			.E(gen[184]),

			.SO(gen[277]),
			.S(gen[278]),
			.SE(gen[279]),

			.SELF(gen[183]),
			.cell_state(gen[183])
		); 

/******************* CELL 184 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell184 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[88]),
			.N(gen[89]),
			.NE(gen[90]),

			.O(gen[183]),
			.E(gen[185]),

			.SO(gen[278]),
			.S(gen[279]),
			.SE(gen[280]),

			.SELF(gen[184]),
			.cell_state(gen[184])
		); 

/******************* CELL 185 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell185 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[89]),
			.N(gen[90]),
			.NE(gen[91]),

			.O(gen[184]),
			.E(gen[186]),

			.SO(gen[279]),
			.S(gen[280]),
			.SE(gen[281]),

			.SELF(gen[185]),
			.cell_state(gen[185])
		); 

/******************* CELL 186 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell186 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[90]),
			.N(gen[91]),
			.NE(gen[92]),

			.O(gen[185]),
			.E(gen[187]),

			.SO(gen[280]),
			.S(gen[281]),
			.SE(gen[282]),

			.SELF(gen[186]),
			.cell_state(gen[186])
		); 

/******************* CELL 187 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell187 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[91]),
			.N(gen[92]),
			.NE(gen[93]),

			.O(gen[186]),
			.E(gen[188]),

			.SO(gen[281]),
			.S(gen[282]),
			.SE(gen[283]),

			.SELF(gen[187]),
			.cell_state(gen[187])
		); 

/******************* CELL 188 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell188 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[92]),
			.N(gen[93]),
			.NE(gen[94]),

			.O(gen[187]),
			.E(gen[189]),

			.SO(gen[282]),
			.S(gen[283]),
			.SE(gen[284]),

			.SELF(gen[188]),
			.cell_state(gen[188])
		); 

/******************* CELL 189 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell189 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[93]),
			.N(gen[94]),
			.NE(gen[93]),

			.O(gen[188]),
			.E(gen[188]),

			.SO(gen[283]),
			.S(gen[284]),
			.SE(gen[283]),

			.SELF(gen[189]),
			.cell_state(gen[189])
		); 

/******************* CELL 190 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell190 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[96]),
			.N(gen[95]),
			.NE(gen[96]),

			.O(gen[191]),
			.E(gen[191]),

			.SO(gen[286]),
			.S(gen[285]),
			.SE(gen[286]),

			.SELF(gen[190]),
			.cell_state(gen[190])
		); 

/******************* CELL 191 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell191 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[95]),
			.N(gen[96]),
			.NE(gen[97]),

			.O(gen[190]),
			.E(gen[192]),

			.SO(gen[285]),
			.S(gen[286]),
			.SE(gen[287]),

			.SELF(gen[191]),
			.cell_state(gen[191])
		); 

/******************* CELL 192 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell192 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[96]),
			.N(gen[97]),
			.NE(gen[98]),

			.O(gen[191]),
			.E(gen[193]),

			.SO(gen[286]),
			.S(gen[287]),
			.SE(gen[288]),

			.SELF(gen[192]),
			.cell_state(gen[192])
		); 

/******************* CELL 193 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell193 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[97]),
			.N(gen[98]),
			.NE(gen[99]),

			.O(gen[192]),
			.E(gen[194]),

			.SO(gen[287]),
			.S(gen[288]),
			.SE(gen[289]),

			.SELF(gen[193]),
			.cell_state(gen[193])
		); 

/******************* CELL 194 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell194 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[98]),
			.N(gen[99]),
			.NE(gen[100]),

			.O(gen[193]),
			.E(gen[195]),

			.SO(gen[288]),
			.S(gen[289]),
			.SE(gen[290]),

			.SELF(gen[194]),
			.cell_state(gen[194])
		); 

/******************* CELL 195 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell195 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[99]),
			.N(gen[100]),
			.NE(gen[101]),

			.O(gen[194]),
			.E(gen[196]),

			.SO(gen[289]),
			.S(gen[290]),
			.SE(gen[291]),

			.SELF(gen[195]),
			.cell_state(gen[195])
		); 

/******************* CELL 196 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell196 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[100]),
			.N(gen[101]),
			.NE(gen[102]),

			.O(gen[195]),
			.E(gen[197]),

			.SO(gen[290]),
			.S(gen[291]),
			.SE(gen[292]),

			.SELF(gen[196]),
			.cell_state(gen[196])
		); 

/******************* CELL 197 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell197 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[101]),
			.N(gen[102]),
			.NE(gen[103]),

			.O(gen[196]),
			.E(gen[198]),

			.SO(gen[291]),
			.S(gen[292]),
			.SE(gen[293]),

			.SELF(gen[197]),
			.cell_state(gen[197])
		); 

/******************* CELL 198 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell198 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[102]),
			.N(gen[103]),
			.NE(gen[104]),

			.O(gen[197]),
			.E(gen[199]),

			.SO(gen[292]),
			.S(gen[293]),
			.SE(gen[294]),

			.SELF(gen[198]),
			.cell_state(gen[198])
		); 

/******************* CELL 199 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell199 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[103]),
			.N(gen[104]),
			.NE(gen[105]),

			.O(gen[198]),
			.E(gen[200]),

			.SO(gen[293]),
			.S(gen[294]),
			.SE(gen[295]),

			.SELF(gen[199]),
			.cell_state(gen[199])
		); 

/******************* CELL 200 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell200 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[104]),
			.N(gen[105]),
			.NE(gen[106]),

			.O(gen[199]),
			.E(gen[201]),

			.SO(gen[294]),
			.S(gen[295]),
			.SE(gen[296]),

			.SELF(gen[200]),
			.cell_state(gen[200])
		); 

/******************* CELL 201 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell201 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[105]),
			.N(gen[106]),
			.NE(gen[107]),

			.O(gen[200]),
			.E(gen[202]),

			.SO(gen[295]),
			.S(gen[296]),
			.SE(gen[297]),

			.SELF(gen[201]),
			.cell_state(gen[201])
		); 

/******************* CELL 202 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell202 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[106]),
			.N(gen[107]),
			.NE(gen[108]),

			.O(gen[201]),
			.E(gen[203]),

			.SO(gen[296]),
			.S(gen[297]),
			.SE(gen[298]),

			.SELF(gen[202]),
			.cell_state(gen[202])
		); 

/******************* CELL 203 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell203 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[107]),
			.N(gen[108]),
			.NE(gen[109]),

			.O(gen[202]),
			.E(gen[204]),

			.SO(gen[297]),
			.S(gen[298]),
			.SE(gen[299]),

			.SELF(gen[203]),
			.cell_state(gen[203])
		); 

/******************* CELL 204 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell204 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[108]),
			.N(gen[109]),
			.NE(gen[110]),

			.O(gen[203]),
			.E(gen[205]),

			.SO(gen[298]),
			.S(gen[299]),
			.SE(gen[300]),

			.SELF(gen[204]),
			.cell_state(gen[204])
		); 

/******************* CELL 205 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell205 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[109]),
			.N(gen[110]),
			.NE(gen[111]),

			.O(gen[204]),
			.E(gen[206]),

			.SO(gen[299]),
			.S(gen[300]),
			.SE(gen[301]),

			.SELF(gen[205]),
			.cell_state(gen[205])
		); 

/******************* CELL 206 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell206 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[110]),
			.N(gen[111]),
			.NE(gen[112]),

			.O(gen[205]),
			.E(gen[207]),

			.SO(gen[300]),
			.S(gen[301]),
			.SE(gen[302]),

			.SELF(gen[206]),
			.cell_state(gen[206])
		); 

/******************* CELL 207 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell207 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[111]),
			.N(gen[112]),
			.NE(gen[113]),

			.O(gen[206]),
			.E(gen[208]),

			.SO(gen[301]),
			.S(gen[302]),
			.SE(gen[303]),

			.SELF(gen[207]),
			.cell_state(gen[207])
		); 

/******************* CELL 208 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell208 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[112]),
			.N(gen[113]),
			.NE(gen[114]),

			.O(gen[207]),
			.E(gen[209]),

			.SO(gen[302]),
			.S(gen[303]),
			.SE(gen[304]),

			.SELF(gen[208]),
			.cell_state(gen[208])
		); 

/******************* CELL 209 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell209 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[113]),
			.N(gen[114]),
			.NE(gen[115]),

			.O(gen[208]),
			.E(gen[210]),

			.SO(gen[303]),
			.S(gen[304]),
			.SE(gen[305]),

			.SELF(gen[209]),
			.cell_state(gen[209])
		); 

/******************* CELL 210 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell210 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[114]),
			.N(gen[115]),
			.NE(gen[116]),

			.O(gen[209]),
			.E(gen[211]),

			.SO(gen[304]),
			.S(gen[305]),
			.SE(gen[306]),

			.SELF(gen[210]),
			.cell_state(gen[210])
		); 

/******************* CELL 211 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell211 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[115]),
			.N(gen[116]),
			.NE(gen[117]),

			.O(gen[210]),
			.E(gen[212]),

			.SO(gen[305]),
			.S(gen[306]),
			.SE(gen[307]),

			.SELF(gen[211]),
			.cell_state(gen[211])
		); 

/******************* CELL 212 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell212 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[116]),
			.N(gen[117]),
			.NE(gen[118]),

			.O(gen[211]),
			.E(gen[213]),

			.SO(gen[306]),
			.S(gen[307]),
			.SE(gen[308]),

			.SELF(gen[212]),
			.cell_state(gen[212])
		); 

/******************* CELL 213 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell213 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[117]),
			.N(gen[118]),
			.NE(gen[119]),

			.O(gen[212]),
			.E(gen[214]),

			.SO(gen[307]),
			.S(gen[308]),
			.SE(gen[309]),

			.SELF(gen[213]),
			.cell_state(gen[213])
		); 

/******************* CELL 214 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell214 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[118]),
			.N(gen[119]),
			.NE(gen[120]),

			.O(gen[213]),
			.E(gen[215]),

			.SO(gen[308]),
			.S(gen[309]),
			.SE(gen[310]),

			.SELF(gen[214]),
			.cell_state(gen[214])
		); 

/******************* CELL 215 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell215 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[119]),
			.N(gen[120]),
			.NE(gen[121]),

			.O(gen[214]),
			.E(gen[216]),

			.SO(gen[309]),
			.S(gen[310]),
			.SE(gen[311]),

			.SELF(gen[215]),
			.cell_state(gen[215])
		); 

/******************* CELL 216 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell216 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[120]),
			.N(gen[121]),
			.NE(gen[122]),

			.O(gen[215]),
			.E(gen[217]),

			.SO(gen[310]),
			.S(gen[311]),
			.SE(gen[312]),

			.SELF(gen[216]),
			.cell_state(gen[216])
		); 

/******************* CELL 217 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell217 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[121]),
			.N(gen[122]),
			.NE(gen[123]),

			.O(gen[216]),
			.E(gen[218]),

			.SO(gen[311]),
			.S(gen[312]),
			.SE(gen[313]),

			.SELF(gen[217]),
			.cell_state(gen[217])
		); 

/******************* CELL 218 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell218 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[122]),
			.N(gen[123]),
			.NE(gen[124]),

			.O(gen[217]),
			.E(gen[219]),

			.SO(gen[312]),
			.S(gen[313]),
			.SE(gen[314]),

			.SELF(gen[218]),
			.cell_state(gen[218])
		); 

/******************* CELL 219 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell219 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[123]),
			.N(gen[124]),
			.NE(gen[125]),

			.O(gen[218]),
			.E(gen[220]),

			.SO(gen[313]),
			.S(gen[314]),
			.SE(gen[315]),

			.SELF(gen[219]),
			.cell_state(gen[219])
		); 

/******************* CELL 220 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell220 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[124]),
			.N(gen[125]),
			.NE(gen[126]),

			.O(gen[219]),
			.E(gen[221]),

			.SO(gen[314]),
			.S(gen[315]),
			.SE(gen[316]),

			.SELF(gen[220]),
			.cell_state(gen[220])
		); 

/******************* CELL 221 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell221 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[125]),
			.N(gen[126]),
			.NE(gen[127]),

			.O(gen[220]),
			.E(gen[222]),

			.SO(gen[315]),
			.S(gen[316]),
			.SE(gen[317]),

			.SELF(gen[221]),
			.cell_state(gen[221])
		); 

/******************* CELL 222 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell222 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[126]),
			.N(gen[127]),
			.NE(gen[128]),

			.O(gen[221]),
			.E(gen[223]),

			.SO(gen[316]),
			.S(gen[317]),
			.SE(gen[318]),

			.SELF(gen[222]),
			.cell_state(gen[222])
		); 

/******************* CELL 223 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell223 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[127]),
			.N(gen[128]),
			.NE(gen[129]),

			.O(gen[222]),
			.E(gen[224]),

			.SO(gen[317]),
			.S(gen[318]),
			.SE(gen[319]),

			.SELF(gen[223]),
			.cell_state(gen[223])
		); 

/******************* CELL 224 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell224 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[128]),
			.N(gen[129]),
			.NE(gen[130]),

			.O(gen[223]),
			.E(gen[225]),

			.SO(gen[318]),
			.S(gen[319]),
			.SE(gen[320]),

			.SELF(gen[224]),
			.cell_state(gen[224])
		); 

/******************* CELL 225 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell225 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[129]),
			.N(gen[130]),
			.NE(gen[131]),

			.O(gen[224]),
			.E(gen[226]),

			.SO(gen[319]),
			.S(gen[320]),
			.SE(gen[321]),

			.SELF(gen[225]),
			.cell_state(gen[225])
		); 

/******************* CELL 226 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell226 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[130]),
			.N(gen[131]),
			.NE(gen[132]),

			.O(gen[225]),
			.E(gen[227]),

			.SO(gen[320]),
			.S(gen[321]),
			.SE(gen[322]),

			.SELF(gen[226]),
			.cell_state(gen[226])
		); 

/******************* CELL 227 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell227 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[131]),
			.N(gen[132]),
			.NE(gen[133]),

			.O(gen[226]),
			.E(gen[228]),

			.SO(gen[321]),
			.S(gen[322]),
			.SE(gen[323]),

			.SELF(gen[227]),
			.cell_state(gen[227])
		); 

/******************* CELL 228 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell228 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[132]),
			.N(gen[133]),
			.NE(gen[134]),

			.O(gen[227]),
			.E(gen[229]),

			.SO(gen[322]),
			.S(gen[323]),
			.SE(gen[324]),

			.SELF(gen[228]),
			.cell_state(gen[228])
		); 

/******************* CELL 229 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell229 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[133]),
			.N(gen[134]),
			.NE(gen[135]),

			.O(gen[228]),
			.E(gen[230]),

			.SO(gen[323]),
			.S(gen[324]),
			.SE(gen[325]),

			.SELF(gen[229]),
			.cell_state(gen[229])
		); 

/******************* CELL 230 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell230 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[134]),
			.N(gen[135]),
			.NE(gen[136]),

			.O(gen[229]),
			.E(gen[231]),

			.SO(gen[324]),
			.S(gen[325]),
			.SE(gen[326]),

			.SELF(gen[230]),
			.cell_state(gen[230])
		); 

/******************* CELL 231 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell231 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[135]),
			.N(gen[136]),
			.NE(gen[137]),

			.O(gen[230]),
			.E(gen[232]),

			.SO(gen[325]),
			.S(gen[326]),
			.SE(gen[327]),

			.SELF(gen[231]),
			.cell_state(gen[231])
		); 

/******************* CELL 232 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell232 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[136]),
			.N(gen[137]),
			.NE(gen[138]),

			.O(gen[231]),
			.E(gen[233]),

			.SO(gen[326]),
			.S(gen[327]),
			.SE(gen[328]),

			.SELF(gen[232]),
			.cell_state(gen[232])
		); 

/******************* CELL 233 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell233 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[137]),
			.N(gen[138]),
			.NE(gen[139]),

			.O(gen[232]),
			.E(gen[234]),

			.SO(gen[327]),
			.S(gen[328]),
			.SE(gen[329]),

			.SELF(gen[233]),
			.cell_state(gen[233])
		); 

/******************* CELL 234 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell234 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[138]),
			.N(gen[139]),
			.NE(gen[140]),

			.O(gen[233]),
			.E(gen[235]),

			.SO(gen[328]),
			.S(gen[329]),
			.SE(gen[330]),

			.SELF(gen[234]),
			.cell_state(gen[234])
		); 

/******************* CELL 235 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell235 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[139]),
			.N(gen[140]),
			.NE(gen[141]),

			.O(gen[234]),
			.E(gen[236]),

			.SO(gen[329]),
			.S(gen[330]),
			.SE(gen[331]),

			.SELF(gen[235]),
			.cell_state(gen[235])
		); 

/******************* CELL 236 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell236 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[140]),
			.N(gen[141]),
			.NE(gen[142]),

			.O(gen[235]),
			.E(gen[237]),

			.SO(gen[330]),
			.S(gen[331]),
			.SE(gen[332]),

			.SELF(gen[236]),
			.cell_state(gen[236])
		); 

/******************* CELL 237 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell237 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[141]),
			.N(gen[142]),
			.NE(gen[143]),

			.O(gen[236]),
			.E(gen[238]),

			.SO(gen[331]),
			.S(gen[332]),
			.SE(gen[333]),

			.SELF(gen[237]),
			.cell_state(gen[237])
		); 

/******************* CELL 238 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell238 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[142]),
			.N(gen[143]),
			.NE(gen[144]),

			.O(gen[237]),
			.E(gen[239]),

			.SO(gen[332]),
			.S(gen[333]),
			.SE(gen[334]),

			.SELF(gen[238]),
			.cell_state(gen[238])
		); 

/******************* CELL 239 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell239 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[143]),
			.N(gen[144]),
			.NE(gen[145]),

			.O(gen[238]),
			.E(gen[240]),

			.SO(gen[333]),
			.S(gen[334]),
			.SE(gen[335]),

			.SELF(gen[239]),
			.cell_state(gen[239])
		); 

/******************* CELL 240 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell240 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[144]),
			.N(gen[145]),
			.NE(gen[146]),

			.O(gen[239]),
			.E(gen[241]),

			.SO(gen[334]),
			.S(gen[335]),
			.SE(gen[336]),

			.SELF(gen[240]),
			.cell_state(gen[240])
		); 

/******************* CELL 241 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell241 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[145]),
			.N(gen[146]),
			.NE(gen[147]),

			.O(gen[240]),
			.E(gen[242]),

			.SO(gen[335]),
			.S(gen[336]),
			.SE(gen[337]),

			.SELF(gen[241]),
			.cell_state(gen[241])
		); 

/******************* CELL 242 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell242 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[146]),
			.N(gen[147]),
			.NE(gen[148]),

			.O(gen[241]),
			.E(gen[243]),

			.SO(gen[336]),
			.S(gen[337]),
			.SE(gen[338]),

			.SELF(gen[242]),
			.cell_state(gen[242])
		); 

/******************* CELL 243 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell243 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[147]),
			.N(gen[148]),
			.NE(gen[149]),

			.O(gen[242]),
			.E(gen[244]),

			.SO(gen[337]),
			.S(gen[338]),
			.SE(gen[339]),

			.SELF(gen[243]),
			.cell_state(gen[243])
		); 

/******************* CELL 244 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell244 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[148]),
			.N(gen[149]),
			.NE(gen[150]),

			.O(gen[243]),
			.E(gen[245]),

			.SO(gen[338]),
			.S(gen[339]),
			.SE(gen[340]),

			.SELF(gen[244]),
			.cell_state(gen[244])
		); 

/******************* CELL 245 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell245 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[149]),
			.N(gen[150]),
			.NE(gen[151]),

			.O(gen[244]),
			.E(gen[246]),

			.SO(gen[339]),
			.S(gen[340]),
			.SE(gen[341]),

			.SELF(gen[245]),
			.cell_state(gen[245])
		); 

/******************* CELL 246 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell246 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[150]),
			.N(gen[151]),
			.NE(gen[152]),

			.O(gen[245]),
			.E(gen[247]),

			.SO(gen[340]),
			.S(gen[341]),
			.SE(gen[342]),

			.SELF(gen[246]),
			.cell_state(gen[246])
		); 

/******************* CELL 247 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell247 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[151]),
			.N(gen[152]),
			.NE(gen[153]),

			.O(gen[246]),
			.E(gen[248]),

			.SO(gen[341]),
			.S(gen[342]),
			.SE(gen[343]),

			.SELF(gen[247]),
			.cell_state(gen[247])
		); 

/******************* CELL 248 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell248 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[152]),
			.N(gen[153]),
			.NE(gen[154]),

			.O(gen[247]),
			.E(gen[249]),

			.SO(gen[342]),
			.S(gen[343]),
			.SE(gen[344]),

			.SELF(gen[248]),
			.cell_state(gen[248])
		); 

/******************* CELL 249 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell249 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[153]),
			.N(gen[154]),
			.NE(gen[155]),

			.O(gen[248]),
			.E(gen[250]),

			.SO(gen[343]),
			.S(gen[344]),
			.SE(gen[345]),

			.SELF(gen[249]),
			.cell_state(gen[249])
		); 

/******************* CELL 250 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell250 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[154]),
			.N(gen[155]),
			.NE(gen[156]),

			.O(gen[249]),
			.E(gen[251]),

			.SO(gen[344]),
			.S(gen[345]),
			.SE(gen[346]),

			.SELF(gen[250]),
			.cell_state(gen[250])
		); 

/******************* CELL 251 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell251 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[155]),
			.N(gen[156]),
			.NE(gen[157]),

			.O(gen[250]),
			.E(gen[252]),

			.SO(gen[345]),
			.S(gen[346]),
			.SE(gen[347]),

			.SELF(gen[251]),
			.cell_state(gen[251])
		); 

/******************* CELL 252 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell252 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[156]),
			.N(gen[157]),
			.NE(gen[158]),

			.O(gen[251]),
			.E(gen[253]),

			.SO(gen[346]),
			.S(gen[347]),
			.SE(gen[348]),

			.SELF(gen[252]),
			.cell_state(gen[252])
		); 

/******************* CELL 253 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell253 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[157]),
			.N(gen[158]),
			.NE(gen[159]),

			.O(gen[252]),
			.E(gen[254]),

			.SO(gen[347]),
			.S(gen[348]),
			.SE(gen[349]),

			.SELF(gen[253]),
			.cell_state(gen[253])
		); 

/******************* CELL 254 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell254 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[158]),
			.N(gen[159]),
			.NE(gen[160]),

			.O(gen[253]),
			.E(gen[255]),

			.SO(gen[348]),
			.S(gen[349]),
			.SE(gen[350]),

			.SELF(gen[254]),
			.cell_state(gen[254])
		); 

/******************* CELL 255 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell255 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[159]),
			.N(gen[160]),
			.NE(gen[161]),

			.O(gen[254]),
			.E(gen[256]),

			.SO(gen[349]),
			.S(gen[350]),
			.SE(gen[351]),

			.SELF(gen[255]),
			.cell_state(gen[255])
		); 

/******************* CELL 256 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell256 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[160]),
			.N(gen[161]),
			.NE(gen[162]),

			.O(gen[255]),
			.E(gen[257]),

			.SO(gen[350]),
			.S(gen[351]),
			.SE(gen[352]),

			.SELF(gen[256]),
			.cell_state(gen[256])
		); 

/******************* CELL 257 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell257 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[161]),
			.N(gen[162]),
			.NE(gen[163]),

			.O(gen[256]),
			.E(gen[258]),

			.SO(gen[351]),
			.S(gen[352]),
			.SE(gen[353]),

			.SELF(gen[257]),
			.cell_state(gen[257])
		); 

/******************* CELL 258 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell258 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[162]),
			.N(gen[163]),
			.NE(gen[164]),

			.O(gen[257]),
			.E(gen[259]),

			.SO(gen[352]),
			.S(gen[353]),
			.SE(gen[354]),

			.SELF(gen[258]),
			.cell_state(gen[258])
		); 

/******************* CELL 259 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell259 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[163]),
			.N(gen[164]),
			.NE(gen[165]),

			.O(gen[258]),
			.E(gen[260]),

			.SO(gen[353]),
			.S(gen[354]),
			.SE(gen[355]),

			.SELF(gen[259]),
			.cell_state(gen[259])
		); 

/******************* CELL 260 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell260 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[164]),
			.N(gen[165]),
			.NE(gen[166]),

			.O(gen[259]),
			.E(gen[261]),

			.SO(gen[354]),
			.S(gen[355]),
			.SE(gen[356]),

			.SELF(gen[260]),
			.cell_state(gen[260])
		); 

/******************* CELL 261 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell261 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[165]),
			.N(gen[166]),
			.NE(gen[167]),

			.O(gen[260]),
			.E(gen[262]),

			.SO(gen[355]),
			.S(gen[356]),
			.SE(gen[357]),

			.SELF(gen[261]),
			.cell_state(gen[261])
		); 

/******************* CELL 262 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell262 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[166]),
			.N(gen[167]),
			.NE(gen[168]),

			.O(gen[261]),
			.E(gen[263]),

			.SO(gen[356]),
			.S(gen[357]),
			.SE(gen[358]),

			.SELF(gen[262]),
			.cell_state(gen[262])
		); 

/******************* CELL 263 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell263 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[167]),
			.N(gen[168]),
			.NE(gen[169]),

			.O(gen[262]),
			.E(gen[264]),

			.SO(gen[357]),
			.S(gen[358]),
			.SE(gen[359]),

			.SELF(gen[263]),
			.cell_state(gen[263])
		); 

/******************* CELL 264 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell264 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[168]),
			.N(gen[169]),
			.NE(gen[170]),

			.O(gen[263]),
			.E(gen[265]),

			.SO(gen[358]),
			.S(gen[359]),
			.SE(gen[360]),

			.SELF(gen[264]),
			.cell_state(gen[264])
		); 

/******************* CELL 265 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell265 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[169]),
			.N(gen[170]),
			.NE(gen[171]),

			.O(gen[264]),
			.E(gen[266]),

			.SO(gen[359]),
			.S(gen[360]),
			.SE(gen[361]),

			.SELF(gen[265]),
			.cell_state(gen[265])
		); 

/******************* CELL 266 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell266 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[170]),
			.N(gen[171]),
			.NE(gen[172]),

			.O(gen[265]),
			.E(gen[267]),

			.SO(gen[360]),
			.S(gen[361]),
			.SE(gen[362]),

			.SELF(gen[266]),
			.cell_state(gen[266])
		); 

/******************* CELL 267 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell267 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[171]),
			.N(gen[172]),
			.NE(gen[173]),

			.O(gen[266]),
			.E(gen[268]),

			.SO(gen[361]),
			.S(gen[362]),
			.SE(gen[363]),

			.SELF(gen[267]),
			.cell_state(gen[267])
		); 

/******************* CELL 268 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell268 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[172]),
			.N(gen[173]),
			.NE(gen[174]),

			.O(gen[267]),
			.E(gen[269]),

			.SO(gen[362]),
			.S(gen[363]),
			.SE(gen[364]),

			.SELF(gen[268]),
			.cell_state(gen[268])
		); 

/******************* CELL 269 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell269 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[173]),
			.N(gen[174]),
			.NE(gen[175]),

			.O(gen[268]),
			.E(gen[270]),

			.SO(gen[363]),
			.S(gen[364]),
			.SE(gen[365]),

			.SELF(gen[269]),
			.cell_state(gen[269])
		); 

/******************* CELL 270 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell270 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[174]),
			.N(gen[175]),
			.NE(gen[176]),

			.O(gen[269]),
			.E(gen[271]),

			.SO(gen[364]),
			.S(gen[365]),
			.SE(gen[366]),

			.SELF(gen[270]),
			.cell_state(gen[270])
		); 

/******************* CELL 271 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell271 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[175]),
			.N(gen[176]),
			.NE(gen[177]),

			.O(gen[270]),
			.E(gen[272]),

			.SO(gen[365]),
			.S(gen[366]),
			.SE(gen[367]),

			.SELF(gen[271]),
			.cell_state(gen[271])
		); 

/******************* CELL 272 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell272 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[176]),
			.N(gen[177]),
			.NE(gen[178]),

			.O(gen[271]),
			.E(gen[273]),

			.SO(gen[366]),
			.S(gen[367]),
			.SE(gen[368]),

			.SELF(gen[272]),
			.cell_state(gen[272])
		); 

/******************* CELL 273 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell273 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[177]),
			.N(gen[178]),
			.NE(gen[179]),

			.O(gen[272]),
			.E(gen[274]),

			.SO(gen[367]),
			.S(gen[368]),
			.SE(gen[369]),

			.SELF(gen[273]),
			.cell_state(gen[273])
		); 

/******************* CELL 274 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell274 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[178]),
			.N(gen[179]),
			.NE(gen[180]),

			.O(gen[273]),
			.E(gen[275]),

			.SO(gen[368]),
			.S(gen[369]),
			.SE(gen[370]),

			.SELF(gen[274]),
			.cell_state(gen[274])
		); 

/******************* CELL 275 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell275 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[179]),
			.N(gen[180]),
			.NE(gen[181]),

			.O(gen[274]),
			.E(gen[276]),

			.SO(gen[369]),
			.S(gen[370]),
			.SE(gen[371]),

			.SELF(gen[275]),
			.cell_state(gen[275])
		); 

/******************* CELL 276 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell276 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[180]),
			.N(gen[181]),
			.NE(gen[182]),

			.O(gen[275]),
			.E(gen[277]),

			.SO(gen[370]),
			.S(gen[371]),
			.SE(gen[372]),

			.SELF(gen[276]),
			.cell_state(gen[276])
		); 

/******************* CELL 277 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell277 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[181]),
			.N(gen[182]),
			.NE(gen[183]),

			.O(gen[276]),
			.E(gen[278]),

			.SO(gen[371]),
			.S(gen[372]),
			.SE(gen[373]),

			.SELF(gen[277]),
			.cell_state(gen[277])
		); 

/******************* CELL 278 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell278 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[182]),
			.N(gen[183]),
			.NE(gen[184]),

			.O(gen[277]),
			.E(gen[279]),

			.SO(gen[372]),
			.S(gen[373]),
			.SE(gen[374]),

			.SELF(gen[278]),
			.cell_state(gen[278])
		); 

/******************* CELL 279 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell279 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[183]),
			.N(gen[184]),
			.NE(gen[185]),

			.O(gen[278]),
			.E(gen[280]),

			.SO(gen[373]),
			.S(gen[374]),
			.SE(gen[375]),

			.SELF(gen[279]),
			.cell_state(gen[279])
		); 

/******************* CELL 280 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell280 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[184]),
			.N(gen[185]),
			.NE(gen[186]),

			.O(gen[279]),
			.E(gen[281]),

			.SO(gen[374]),
			.S(gen[375]),
			.SE(gen[376]),

			.SELF(gen[280]),
			.cell_state(gen[280])
		); 

/******************* CELL 281 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell281 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[185]),
			.N(gen[186]),
			.NE(gen[187]),

			.O(gen[280]),
			.E(gen[282]),

			.SO(gen[375]),
			.S(gen[376]),
			.SE(gen[377]),

			.SELF(gen[281]),
			.cell_state(gen[281])
		); 

/******************* CELL 282 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell282 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[186]),
			.N(gen[187]),
			.NE(gen[188]),

			.O(gen[281]),
			.E(gen[283]),

			.SO(gen[376]),
			.S(gen[377]),
			.SE(gen[378]),

			.SELF(gen[282]),
			.cell_state(gen[282])
		); 

/******************* CELL 283 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell283 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[187]),
			.N(gen[188]),
			.NE(gen[189]),

			.O(gen[282]),
			.E(gen[284]),

			.SO(gen[377]),
			.S(gen[378]),
			.SE(gen[379]),

			.SELF(gen[283]),
			.cell_state(gen[283])
		); 

/******************* CELL 284 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell284 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[188]),
			.N(gen[189]),
			.NE(gen[188]),

			.O(gen[283]),
			.E(gen[283]),

			.SO(gen[378]),
			.S(gen[379]),
			.SE(gen[378]),

			.SELF(gen[284]),
			.cell_state(gen[284])
		); 

/******************* CELL 285 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell285 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[191]),
			.N(gen[190]),
			.NE(gen[191]),

			.O(gen[286]),
			.E(gen[286]),

			.SO(gen[381]),
			.S(gen[380]),
			.SE(gen[381]),

			.SELF(gen[285]),
			.cell_state(gen[285])
		); 

/******************* CELL 286 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell286 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[190]),
			.N(gen[191]),
			.NE(gen[192]),

			.O(gen[285]),
			.E(gen[287]),

			.SO(gen[380]),
			.S(gen[381]),
			.SE(gen[382]),

			.SELF(gen[286]),
			.cell_state(gen[286])
		); 

/******************* CELL 287 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell287 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[191]),
			.N(gen[192]),
			.NE(gen[193]),

			.O(gen[286]),
			.E(gen[288]),

			.SO(gen[381]),
			.S(gen[382]),
			.SE(gen[383]),

			.SELF(gen[287]),
			.cell_state(gen[287])
		); 

/******************* CELL 288 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell288 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[192]),
			.N(gen[193]),
			.NE(gen[194]),

			.O(gen[287]),
			.E(gen[289]),

			.SO(gen[382]),
			.S(gen[383]),
			.SE(gen[384]),

			.SELF(gen[288]),
			.cell_state(gen[288])
		); 

/******************* CELL 289 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell289 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[193]),
			.N(gen[194]),
			.NE(gen[195]),

			.O(gen[288]),
			.E(gen[290]),

			.SO(gen[383]),
			.S(gen[384]),
			.SE(gen[385]),

			.SELF(gen[289]),
			.cell_state(gen[289])
		); 

/******************* CELL 290 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell290 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[194]),
			.N(gen[195]),
			.NE(gen[196]),

			.O(gen[289]),
			.E(gen[291]),

			.SO(gen[384]),
			.S(gen[385]),
			.SE(gen[386]),

			.SELF(gen[290]),
			.cell_state(gen[290])
		); 

/******************* CELL 291 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell291 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[195]),
			.N(gen[196]),
			.NE(gen[197]),

			.O(gen[290]),
			.E(gen[292]),

			.SO(gen[385]),
			.S(gen[386]),
			.SE(gen[387]),

			.SELF(gen[291]),
			.cell_state(gen[291])
		); 

/******************* CELL 292 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell292 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[196]),
			.N(gen[197]),
			.NE(gen[198]),

			.O(gen[291]),
			.E(gen[293]),

			.SO(gen[386]),
			.S(gen[387]),
			.SE(gen[388]),

			.SELF(gen[292]),
			.cell_state(gen[292])
		); 

/******************* CELL 293 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell293 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[197]),
			.N(gen[198]),
			.NE(gen[199]),

			.O(gen[292]),
			.E(gen[294]),

			.SO(gen[387]),
			.S(gen[388]),
			.SE(gen[389]),

			.SELF(gen[293]),
			.cell_state(gen[293])
		); 

/******************* CELL 294 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell294 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[198]),
			.N(gen[199]),
			.NE(gen[200]),

			.O(gen[293]),
			.E(gen[295]),

			.SO(gen[388]),
			.S(gen[389]),
			.SE(gen[390]),

			.SELF(gen[294]),
			.cell_state(gen[294])
		); 

/******************* CELL 295 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell295 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[199]),
			.N(gen[200]),
			.NE(gen[201]),

			.O(gen[294]),
			.E(gen[296]),

			.SO(gen[389]),
			.S(gen[390]),
			.SE(gen[391]),

			.SELF(gen[295]),
			.cell_state(gen[295])
		); 

/******************* CELL 296 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell296 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[200]),
			.N(gen[201]),
			.NE(gen[202]),

			.O(gen[295]),
			.E(gen[297]),

			.SO(gen[390]),
			.S(gen[391]),
			.SE(gen[392]),

			.SELF(gen[296]),
			.cell_state(gen[296])
		); 

/******************* CELL 297 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell297 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[201]),
			.N(gen[202]),
			.NE(gen[203]),

			.O(gen[296]),
			.E(gen[298]),

			.SO(gen[391]),
			.S(gen[392]),
			.SE(gen[393]),

			.SELF(gen[297]),
			.cell_state(gen[297])
		); 

/******************* CELL 298 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell298 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[202]),
			.N(gen[203]),
			.NE(gen[204]),

			.O(gen[297]),
			.E(gen[299]),

			.SO(gen[392]),
			.S(gen[393]),
			.SE(gen[394]),

			.SELF(gen[298]),
			.cell_state(gen[298])
		); 

/******************* CELL 299 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell299 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[203]),
			.N(gen[204]),
			.NE(gen[205]),

			.O(gen[298]),
			.E(gen[300]),

			.SO(gen[393]),
			.S(gen[394]),
			.SE(gen[395]),

			.SELF(gen[299]),
			.cell_state(gen[299])
		); 

/******************* CELL 300 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell300 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[204]),
			.N(gen[205]),
			.NE(gen[206]),

			.O(gen[299]),
			.E(gen[301]),

			.SO(gen[394]),
			.S(gen[395]),
			.SE(gen[396]),

			.SELF(gen[300]),
			.cell_state(gen[300])
		); 

/******************* CELL 301 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell301 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[205]),
			.N(gen[206]),
			.NE(gen[207]),

			.O(gen[300]),
			.E(gen[302]),

			.SO(gen[395]),
			.S(gen[396]),
			.SE(gen[397]),

			.SELF(gen[301]),
			.cell_state(gen[301])
		); 

/******************* CELL 302 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell302 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[206]),
			.N(gen[207]),
			.NE(gen[208]),

			.O(gen[301]),
			.E(gen[303]),

			.SO(gen[396]),
			.S(gen[397]),
			.SE(gen[398]),

			.SELF(gen[302]),
			.cell_state(gen[302])
		); 

/******************* CELL 303 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell303 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[207]),
			.N(gen[208]),
			.NE(gen[209]),

			.O(gen[302]),
			.E(gen[304]),

			.SO(gen[397]),
			.S(gen[398]),
			.SE(gen[399]),

			.SELF(gen[303]),
			.cell_state(gen[303])
		); 

/******************* CELL 304 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell304 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[208]),
			.N(gen[209]),
			.NE(gen[210]),

			.O(gen[303]),
			.E(gen[305]),

			.SO(gen[398]),
			.S(gen[399]),
			.SE(gen[400]),

			.SELF(gen[304]),
			.cell_state(gen[304])
		); 

/******************* CELL 305 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell305 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[209]),
			.N(gen[210]),
			.NE(gen[211]),

			.O(gen[304]),
			.E(gen[306]),

			.SO(gen[399]),
			.S(gen[400]),
			.SE(gen[401]),

			.SELF(gen[305]),
			.cell_state(gen[305])
		); 

/******************* CELL 306 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell306 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[210]),
			.N(gen[211]),
			.NE(gen[212]),

			.O(gen[305]),
			.E(gen[307]),

			.SO(gen[400]),
			.S(gen[401]),
			.SE(gen[402]),

			.SELF(gen[306]),
			.cell_state(gen[306])
		); 

/******************* CELL 307 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell307 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[211]),
			.N(gen[212]),
			.NE(gen[213]),

			.O(gen[306]),
			.E(gen[308]),

			.SO(gen[401]),
			.S(gen[402]),
			.SE(gen[403]),

			.SELF(gen[307]),
			.cell_state(gen[307])
		); 

/******************* CELL 308 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell308 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[212]),
			.N(gen[213]),
			.NE(gen[214]),

			.O(gen[307]),
			.E(gen[309]),

			.SO(gen[402]),
			.S(gen[403]),
			.SE(gen[404]),

			.SELF(gen[308]),
			.cell_state(gen[308])
		); 

/******************* CELL 309 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell309 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[213]),
			.N(gen[214]),
			.NE(gen[215]),

			.O(gen[308]),
			.E(gen[310]),

			.SO(gen[403]),
			.S(gen[404]),
			.SE(gen[405]),

			.SELF(gen[309]),
			.cell_state(gen[309])
		); 

/******************* CELL 310 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell310 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[214]),
			.N(gen[215]),
			.NE(gen[216]),

			.O(gen[309]),
			.E(gen[311]),

			.SO(gen[404]),
			.S(gen[405]),
			.SE(gen[406]),

			.SELF(gen[310]),
			.cell_state(gen[310])
		); 

/******************* CELL 311 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell311 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[215]),
			.N(gen[216]),
			.NE(gen[217]),

			.O(gen[310]),
			.E(gen[312]),

			.SO(gen[405]),
			.S(gen[406]),
			.SE(gen[407]),

			.SELF(gen[311]),
			.cell_state(gen[311])
		); 

/******************* CELL 312 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell312 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[216]),
			.N(gen[217]),
			.NE(gen[218]),

			.O(gen[311]),
			.E(gen[313]),

			.SO(gen[406]),
			.S(gen[407]),
			.SE(gen[408]),

			.SELF(gen[312]),
			.cell_state(gen[312])
		); 

/******************* CELL 313 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell313 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[217]),
			.N(gen[218]),
			.NE(gen[219]),

			.O(gen[312]),
			.E(gen[314]),

			.SO(gen[407]),
			.S(gen[408]),
			.SE(gen[409]),

			.SELF(gen[313]),
			.cell_state(gen[313])
		); 

/******************* CELL 314 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell314 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[218]),
			.N(gen[219]),
			.NE(gen[220]),

			.O(gen[313]),
			.E(gen[315]),

			.SO(gen[408]),
			.S(gen[409]),
			.SE(gen[410]),

			.SELF(gen[314]),
			.cell_state(gen[314])
		); 

/******************* CELL 315 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell315 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[219]),
			.N(gen[220]),
			.NE(gen[221]),

			.O(gen[314]),
			.E(gen[316]),

			.SO(gen[409]),
			.S(gen[410]),
			.SE(gen[411]),

			.SELF(gen[315]),
			.cell_state(gen[315])
		); 

/******************* CELL 316 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell316 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[220]),
			.N(gen[221]),
			.NE(gen[222]),

			.O(gen[315]),
			.E(gen[317]),

			.SO(gen[410]),
			.S(gen[411]),
			.SE(gen[412]),

			.SELF(gen[316]),
			.cell_state(gen[316])
		); 

/******************* CELL 317 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell317 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[221]),
			.N(gen[222]),
			.NE(gen[223]),

			.O(gen[316]),
			.E(gen[318]),

			.SO(gen[411]),
			.S(gen[412]),
			.SE(gen[413]),

			.SELF(gen[317]),
			.cell_state(gen[317])
		); 

/******************* CELL 318 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell318 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[222]),
			.N(gen[223]),
			.NE(gen[224]),

			.O(gen[317]),
			.E(gen[319]),

			.SO(gen[412]),
			.S(gen[413]),
			.SE(gen[414]),

			.SELF(gen[318]),
			.cell_state(gen[318])
		); 

/******************* CELL 319 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell319 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[223]),
			.N(gen[224]),
			.NE(gen[225]),

			.O(gen[318]),
			.E(gen[320]),

			.SO(gen[413]),
			.S(gen[414]),
			.SE(gen[415]),

			.SELF(gen[319]),
			.cell_state(gen[319])
		); 

/******************* CELL 320 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell320 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[224]),
			.N(gen[225]),
			.NE(gen[226]),

			.O(gen[319]),
			.E(gen[321]),

			.SO(gen[414]),
			.S(gen[415]),
			.SE(gen[416]),

			.SELF(gen[320]),
			.cell_state(gen[320])
		); 

/******************* CELL 321 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell321 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[225]),
			.N(gen[226]),
			.NE(gen[227]),

			.O(gen[320]),
			.E(gen[322]),

			.SO(gen[415]),
			.S(gen[416]),
			.SE(gen[417]),

			.SELF(gen[321]),
			.cell_state(gen[321])
		); 

/******************* CELL 322 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell322 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[226]),
			.N(gen[227]),
			.NE(gen[228]),

			.O(gen[321]),
			.E(gen[323]),

			.SO(gen[416]),
			.S(gen[417]),
			.SE(gen[418]),

			.SELF(gen[322]),
			.cell_state(gen[322])
		); 

/******************* CELL 323 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell323 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[227]),
			.N(gen[228]),
			.NE(gen[229]),

			.O(gen[322]),
			.E(gen[324]),

			.SO(gen[417]),
			.S(gen[418]),
			.SE(gen[419]),

			.SELF(gen[323]),
			.cell_state(gen[323])
		); 

/******************* CELL 324 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell324 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[228]),
			.N(gen[229]),
			.NE(gen[230]),

			.O(gen[323]),
			.E(gen[325]),

			.SO(gen[418]),
			.S(gen[419]),
			.SE(gen[420]),

			.SELF(gen[324]),
			.cell_state(gen[324])
		); 

/******************* CELL 325 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell325 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[229]),
			.N(gen[230]),
			.NE(gen[231]),

			.O(gen[324]),
			.E(gen[326]),

			.SO(gen[419]),
			.S(gen[420]),
			.SE(gen[421]),

			.SELF(gen[325]),
			.cell_state(gen[325])
		); 

/******************* CELL 326 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell326 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[230]),
			.N(gen[231]),
			.NE(gen[232]),

			.O(gen[325]),
			.E(gen[327]),

			.SO(gen[420]),
			.S(gen[421]),
			.SE(gen[422]),

			.SELF(gen[326]),
			.cell_state(gen[326])
		); 

/******************* CELL 327 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell327 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[231]),
			.N(gen[232]),
			.NE(gen[233]),

			.O(gen[326]),
			.E(gen[328]),

			.SO(gen[421]),
			.S(gen[422]),
			.SE(gen[423]),

			.SELF(gen[327]),
			.cell_state(gen[327])
		); 

/******************* CELL 328 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell328 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[232]),
			.N(gen[233]),
			.NE(gen[234]),

			.O(gen[327]),
			.E(gen[329]),

			.SO(gen[422]),
			.S(gen[423]),
			.SE(gen[424]),

			.SELF(gen[328]),
			.cell_state(gen[328])
		); 

/******************* CELL 329 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell329 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[233]),
			.N(gen[234]),
			.NE(gen[235]),

			.O(gen[328]),
			.E(gen[330]),

			.SO(gen[423]),
			.S(gen[424]),
			.SE(gen[425]),

			.SELF(gen[329]),
			.cell_state(gen[329])
		); 

/******************* CELL 330 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell330 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[234]),
			.N(gen[235]),
			.NE(gen[236]),

			.O(gen[329]),
			.E(gen[331]),

			.SO(gen[424]),
			.S(gen[425]),
			.SE(gen[426]),

			.SELF(gen[330]),
			.cell_state(gen[330])
		); 

/******************* CELL 331 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell331 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[235]),
			.N(gen[236]),
			.NE(gen[237]),

			.O(gen[330]),
			.E(gen[332]),

			.SO(gen[425]),
			.S(gen[426]),
			.SE(gen[427]),

			.SELF(gen[331]),
			.cell_state(gen[331])
		); 

/******************* CELL 332 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell332 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[236]),
			.N(gen[237]),
			.NE(gen[238]),

			.O(gen[331]),
			.E(gen[333]),

			.SO(gen[426]),
			.S(gen[427]),
			.SE(gen[428]),

			.SELF(gen[332]),
			.cell_state(gen[332])
		); 

/******************* CELL 333 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell333 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[237]),
			.N(gen[238]),
			.NE(gen[239]),

			.O(gen[332]),
			.E(gen[334]),

			.SO(gen[427]),
			.S(gen[428]),
			.SE(gen[429]),

			.SELF(gen[333]),
			.cell_state(gen[333])
		); 

/******************* CELL 334 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell334 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[238]),
			.N(gen[239]),
			.NE(gen[240]),

			.O(gen[333]),
			.E(gen[335]),

			.SO(gen[428]),
			.S(gen[429]),
			.SE(gen[430]),

			.SELF(gen[334]),
			.cell_state(gen[334])
		); 

/******************* CELL 335 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell335 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[239]),
			.N(gen[240]),
			.NE(gen[241]),

			.O(gen[334]),
			.E(gen[336]),

			.SO(gen[429]),
			.S(gen[430]),
			.SE(gen[431]),

			.SELF(gen[335]),
			.cell_state(gen[335])
		); 

/******************* CELL 336 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell336 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[240]),
			.N(gen[241]),
			.NE(gen[242]),

			.O(gen[335]),
			.E(gen[337]),

			.SO(gen[430]),
			.S(gen[431]),
			.SE(gen[432]),

			.SELF(gen[336]),
			.cell_state(gen[336])
		); 

/******************* CELL 337 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell337 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[241]),
			.N(gen[242]),
			.NE(gen[243]),

			.O(gen[336]),
			.E(gen[338]),

			.SO(gen[431]),
			.S(gen[432]),
			.SE(gen[433]),

			.SELF(gen[337]),
			.cell_state(gen[337])
		); 

/******************* CELL 338 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell338 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[242]),
			.N(gen[243]),
			.NE(gen[244]),

			.O(gen[337]),
			.E(gen[339]),

			.SO(gen[432]),
			.S(gen[433]),
			.SE(gen[434]),

			.SELF(gen[338]),
			.cell_state(gen[338])
		); 

/******************* CELL 339 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell339 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[243]),
			.N(gen[244]),
			.NE(gen[245]),

			.O(gen[338]),
			.E(gen[340]),

			.SO(gen[433]),
			.S(gen[434]),
			.SE(gen[435]),

			.SELF(gen[339]),
			.cell_state(gen[339])
		); 

/******************* CELL 340 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell340 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[244]),
			.N(gen[245]),
			.NE(gen[246]),

			.O(gen[339]),
			.E(gen[341]),

			.SO(gen[434]),
			.S(gen[435]),
			.SE(gen[436]),

			.SELF(gen[340]),
			.cell_state(gen[340])
		); 

/******************* CELL 341 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell341 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[245]),
			.N(gen[246]),
			.NE(gen[247]),

			.O(gen[340]),
			.E(gen[342]),

			.SO(gen[435]),
			.S(gen[436]),
			.SE(gen[437]),

			.SELF(gen[341]),
			.cell_state(gen[341])
		); 

/******************* CELL 342 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell342 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[246]),
			.N(gen[247]),
			.NE(gen[248]),

			.O(gen[341]),
			.E(gen[343]),

			.SO(gen[436]),
			.S(gen[437]),
			.SE(gen[438]),

			.SELF(gen[342]),
			.cell_state(gen[342])
		); 

/******************* CELL 343 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell343 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[247]),
			.N(gen[248]),
			.NE(gen[249]),

			.O(gen[342]),
			.E(gen[344]),

			.SO(gen[437]),
			.S(gen[438]),
			.SE(gen[439]),

			.SELF(gen[343]),
			.cell_state(gen[343])
		); 

/******************* CELL 344 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell344 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[248]),
			.N(gen[249]),
			.NE(gen[250]),

			.O(gen[343]),
			.E(gen[345]),

			.SO(gen[438]),
			.S(gen[439]),
			.SE(gen[440]),

			.SELF(gen[344]),
			.cell_state(gen[344])
		); 

/******************* CELL 345 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell345 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[249]),
			.N(gen[250]),
			.NE(gen[251]),

			.O(gen[344]),
			.E(gen[346]),

			.SO(gen[439]),
			.S(gen[440]),
			.SE(gen[441]),

			.SELF(gen[345]),
			.cell_state(gen[345])
		); 

/******************* CELL 346 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell346 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[250]),
			.N(gen[251]),
			.NE(gen[252]),

			.O(gen[345]),
			.E(gen[347]),

			.SO(gen[440]),
			.S(gen[441]),
			.SE(gen[442]),

			.SELF(gen[346]),
			.cell_state(gen[346])
		); 

/******************* CELL 347 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell347 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[251]),
			.N(gen[252]),
			.NE(gen[253]),

			.O(gen[346]),
			.E(gen[348]),

			.SO(gen[441]),
			.S(gen[442]),
			.SE(gen[443]),

			.SELF(gen[347]),
			.cell_state(gen[347])
		); 

/******************* CELL 348 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell348 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[252]),
			.N(gen[253]),
			.NE(gen[254]),

			.O(gen[347]),
			.E(gen[349]),

			.SO(gen[442]),
			.S(gen[443]),
			.SE(gen[444]),

			.SELF(gen[348]),
			.cell_state(gen[348])
		); 

/******************* CELL 349 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell349 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[253]),
			.N(gen[254]),
			.NE(gen[255]),

			.O(gen[348]),
			.E(gen[350]),

			.SO(gen[443]),
			.S(gen[444]),
			.SE(gen[445]),

			.SELF(gen[349]),
			.cell_state(gen[349])
		); 

/******************* CELL 350 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell350 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[254]),
			.N(gen[255]),
			.NE(gen[256]),

			.O(gen[349]),
			.E(gen[351]),

			.SO(gen[444]),
			.S(gen[445]),
			.SE(gen[446]),

			.SELF(gen[350]),
			.cell_state(gen[350])
		); 

/******************* CELL 351 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell351 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[255]),
			.N(gen[256]),
			.NE(gen[257]),

			.O(gen[350]),
			.E(gen[352]),

			.SO(gen[445]),
			.S(gen[446]),
			.SE(gen[447]),

			.SELF(gen[351]),
			.cell_state(gen[351])
		); 

/******************* CELL 352 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell352 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[256]),
			.N(gen[257]),
			.NE(gen[258]),

			.O(gen[351]),
			.E(gen[353]),

			.SO(gen[446]),
			.S(gen[447]),
			.SE(gen[448]),

			.SELF(gen[352]),
			.cell_state(gen[352])
		); 

/******************* CELL 353 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell353 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[257]),
			.N(gen[258]),
			.NE(gen[259]),

			.O(gen[352]),
			.E(gen[354]),

			.SO(gen[447]),
			.S(gen[448]),
			.SE(gen[449]),

			.SELF(gen[353]),
			.cell_state(gen[353])
		); 

/******************* CELL 354 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell354 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[258]),
			.N(gen[259]),
			.NE(gen[260]),

			.O(gen[353]),
			.E(gen[355]),

			.SO(gen[448]),
			.S(gen[449]),
			.SE(gen[450]),

			.SELF(gen[354]),
			.cell_state(gen[354])
		); 

/******************* CELL 355 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell355 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[259]),
			.N(gen[260]),
			.NE(gen[261]),

			.O(gen[354]),
			.E(gen[356]),

			.SO(gen[449]),
			.S(gen[450]),
			.SE(gen[451]),

			.SELF(gen[355]),
			.cell_state(gen[355])
		); 

/******************* CELL 356 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell356 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[260]),
			.N(gen[261]),
			.NE(gen[262]),

			.O(gen[355]),
			.E(gen[357]),

			.SO(gen[450]),
			.S(gen[451]),
			.SE(gen[452]),

			.SELF(gen[356]),
			.cell_state(gen[356])
		); 

/******************* CELL 357 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell357 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[261]),
			.N(gen[262]),
			.NE(gen[263]),

			.O(gen[356]),
			.E(gen[358]),

			.SO(gen[451]),
			.S(gen[452]),
			.SE(gen[453]),

			.SELF(gen[357]),
			.cell_state(gen[357])
		); 

/******************* CELL 358 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell358 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[262]),
			.N(gen[263]),
			.NE(gen[264]),

			.O(gen[357]),
			.E(gen[359]),

			.SO(gen[452]),
			.S(gen[453]),
			.SE(gen[454]),

			.SELF(gen[358]),
			.cell_state(gen[358])
		); 

/******************* CELL 359 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell359 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[263]),
			.N(gen[264]),
			.NE(gen[265]),

			.O(gen[358]),
			.E(gen[360]),

			.SO(gen[453]),
			.S(gen[454]),
			.SE(gen[455]),

			.SELF(gen[359]),
			.cell_state(gen[359])
		); 

/******************* CELL 360 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell360 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[264]),
			.N(gen[265]),
			.NE(gen[266]),

			.O(gen[359]),
			.E(gen[361]),

			.SO(gen[454]),
			.S(gen[455]),
			.SE(gen[456]),

			.SELF(gen[360]),
			.cell_state(gen[360])
		); 

/******************* CELL 361 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell361 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[265]),
			.N(gen[266]),
			.NE(gen[267]),

			.O(gen[360]),
			.E(gen[362]),

			.SO(gen[455]),
			.S(gen[456]),
			.SE(gen[457]),

			.SELF(gen[361]),
			.cell_state(gen[361])
		); 

/******************* CELL 362 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell362 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[266]),
			.N(gen[267]),
			.NE(gen[268]),

			.O(gen[361]),
			.E(gen[363]),

			.SO(gen[456]),
			.S(gen[457]),
			.SE(gen[458]),

			.SELF(gen[362]),
			.cell_state(gen[362])
		); 

/******************* CELL 363 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell363 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[267]),
			.N(gen[268]),
			.NE(gen[269]),

			.O(gen[362]),
			.E(gen[364]),

			.SO(gen[457]),
			.S(gen[458]),
			.SE(gen[459]),

			.SELF(gen[363]),
			.cell_state(gen[363])
		); 

/******************* CELL 364 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell364 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[268]),
			.N(gen[269]),
			.NE(gen[270]),

			.O(gen[363]),
			.E(gen[365]),

			.SO(gen[458]),
			.S(gen[459]),
			.SE(gen[460]),

			.SELF(gen[364]),
			.cell_state(gen[364])
		); 

/******************* CELL 365 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell365 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[269]),
			.N(gen[270]),
			.NE(gen[271]),

			.O(gen[364]),
			.E(gen[366]),

			.SO(gen[459]),
			.S(gen[460]),
			.SE(gen[461]),

			.SELF(gen[365]),
			.cell_state(gen[365])
		); 

/******************* CELL 366 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell366 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[270]),
			.N(gen[271]),
			.NE(gen[272]),

			.O(gen[365]),
			.E(gen[367]),

			.SO(gen[460]),
			.S(gen[461]),
			.SE(gen[462]),

			.SELF(gen[366]),
			.cell_state(gen[366])
		); 

/******************* CELL 367 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell367 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[271]),
			.N(gen[272]),
			.NE(gen[273]),

			.O(gen[366]),
			.E(gen[368]),

			.SO(gen[461]),
			.S(gen[462]),
			.SE(gen[463]),

			.SELF(gen[367]),
			.cell_state(gen[367])
		); 

/******************* CELL 368 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell368 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[272]),
			.N(gen[273]),
			.NE(gen[274]),

			.O(gen[367]),
			.E(gen[369]),

			.SO(gen[462]),
			.S(gen[463]),
			.SE(gen[464]),

			.SELF(gen[368]),
			.cell_state(gen[368])
		); 

/******************* CELL 369 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell369 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[273]),
			.N(gen[274]),
			.NE(gen[275]),

			.O(gen[368]),
			.E(gen[370]),

			.SO(gen[463]),
			.S(gen[464]),
			.SE(gen[465]),

			.SELF(gen[369]),
			.cell_state(gen[369])
		); 

/******************* CELL 370 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell370 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[274]),
			.N(gen[275]),
			.NE(gen[276]),

			.O(gen[369]),
			.E(gen[371]),

			.SO(gen[464]),
			.S(gen[465]),
			.SE(gen[466]),

			.SELF(gen[370]),
			.cell_state(gen[370])
		); 

/******************* CELL 371 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell371 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[275]),
			.N(gen[276]),
			.NE(gen[277]),

			.O(gen[370]),
			.E(gen[372]),

			.SO(gen[465]),
			.S(gen[466]),
			.SE(gen[467]),

			.SELF(gen[371]),
			.cell_state(gen[371])
		); 

/******************* CELL 372 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell372 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[276]),
			.N(gen[277]),
			.NE(gen[278]),

			.O(gen[371]),
			.E(gen[373]),

			.SO(gen[466]),
			.S(gen[467]),
			.SE(gen[468]),

			.SELF(gen[372]),
			.cell_state(gen[372])
		); 

/******************* CELL 373 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell373 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[277]),
			.N(gen[278]),
			.NE(gen[279]),

			.O(gen[372]),
			.E(gen[374]),

			.SO(gen[467]),
			.S(gen[468]),
			.SE(gen[469]),

			.SELF(gen[373]),
			.cell_state(gen[373])
		); 

/******************* CELL 374 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell374 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[278]),
			.N(gen[279]),
			.NE(gen[280]),

			.O(gen[373]),
			.E(gen[375]),

			.SO(gen[468]),
			.S(gen[469]),
			.SE(gen[470]),

			.SELF(gen[374]),
			.cell_state(gen[374])
		); 

/******************* CELL 375 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell375 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[279]),
			.N(gen[280]),
			.NE(gen[281]),

			.O(gen[374]),
			.E(gen[376]),

			.SO(gen[469]),
			.S(gen[470]),
			.SE(gen[471]),

			.SELF(gen[375]),
			.cell_state(gen[375])
		); 

/******************* CELL 376 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell376 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[280]),
			.N(gen[281]),
			.NE(gen[282]),

			.O(gen[375]),
			.E(gen[377]),

			.SO(gen[470]),
			.S(gen[471]),
			.SE(gen[472]),

			.SELF(gen[376]),
			.cell_state(gen[376])
		); 

/******************* CELL 377 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell377 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[281]),
			.N(gen[282]),
			.NE(gen[283]),

			.O(gen[376]),
			.E(gen[378]),

			.SO(gen[471]),
			.S(gen[472]),
			.SE(gen[473]),

			.SELF(gen[377]),
			.cell_state(gen[377])
		); 

/******************* CELL 378 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell378 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[282]),
			.N(gen[283]),
			.NE(gen[284]),

			.O(gen[377]),
			.E(gen[379]),

			.SO(gen[472]),
			.S(gen[473]),
			.SE(gen[474]),

			.SELF(gen[378]),
			.cell_state(gen[378])
		); 

/******************* CELL 379 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell379 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[283]),
			.N(gen[284]),
			.NE(gen[283]),

			.O(gen[378]),
			.E(gen[378]),

			.SO(gen[473]),
			.S(gen[474]),
			.SE(gen[473]),

			.SELF(gen[379]),
			.cell_state(gen[379])
		); 

/******************* CELL 380 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell380 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[286]),
			.N(gen[285]),
			.NE(gen[286]),

			.O(gen[381]),
			.E(gen[381]),

			.SO(gen[476]),
			.S(gen[475]),
			.SE(gen[476]),

			.SELF(gen[380]),
			.cell_state(gen[380])
		); 

/******************* CELL 381 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell381 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[285]),
			.N(gen[286]),
			.NE(gen[287]),

			.O(gen[380]),
			.E(gen[382]),

			.SO(gen[475]),
			.S(gen[476]),
			.SE(gen[477]),

			.SELF(gen[381]),
			.cell_state(gen[381])
		); 

/******************* CELL 382 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell382 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[286]),
			.N(gen[287]),
			.NE(gen[288]),

			.O(gen[381]),
			.E(gen[383]),

			.SO(gen[476]),
			.S(gen[477]),
			.SE(gen[478]),

			.SELF(gen[382]),
			.cell_state(gen[382])
		); 

/******************* CELL 383 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell383 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[287]),
			.N(gen[288]),
			.NE(gen[289]),

			.O(gen[382]),
			.E(gen[384]),

			.SO(gen[477]),
			.S(gen[478]),
			.SE(gen[479]),

			.SELF(gen[383]),
			.cell_state(gen[383])
		); 

/******************* CELL 384 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell384 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[288]),
			.N(gen[289]),
			.NE(gen[290]),

			.O(gen[383]),
			.E(gen[385]),

			.SO(gen[478]),
			.S(gen[479]),
			.SE(gen[480]),

			.SELF(gen[384]),
			.cell_state(gen[384])
		); 

/******************* CELL 385 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell385 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[289]),
			.N(gen[290]),
			.NE(gen[291]),

			.O(gen[384]),
			.E(gen[386]),

			.SO(gen[479]),
			.S(gen[480]),
			.SE(gen[481]),

			.SELF(gen[385]),
			.cell_state(gen[385])
		); 

/******************* CELL 386 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell386 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[290]),
			.N(gen[291]),
			.NE(gen[292]),

			.O(gen[385]),
			.E(gen[387]),

			.SO(gen[480]),
			.S(gen[481]),
			.SE(gen[482]),

			.SELF(gen[386]),
			.cell_state(gen[386])
		); 

/******************* CELL 387 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell387 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[291]),
			.N(gen[292]),
			.NE(gen[293]),

			.O(gen[386]),
			.E(gen[388]),

			.SO(gen[481]),
			.S(gen[482]),
			.SE(gen[483]),

			.SELF(gen[387]),
			.cell_state(gen[387])
		); 

/******************* CELL 388 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell388 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[292]),
			.N(gen[293]),
			.NE(gen[294]),

			.O(gen[387]),
			.E(gen[389]),

			.SO(gen[482]),
			.S(gen[483]),
			.SE(gen[484]),

			.SELF(gen[388]),
			.cell_state(gen[388])
		); 

/******************* CELL 389 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell389 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[293]),
			.N(gen[294]),
			.NE(gen[295]),

			.O(gen[388]),
			.E(gen[390]),

			.SO(gen[483]),
			.S(gen[484]),
			.SE(gen[485]),

			.SELF(gen[389]),
			.cell_state(gen[389])
		); 

/******************* CELL 390 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell390 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[294]),
			.N(gen[295]),
			.NE(gen[296]),

			.O(gen[389]),
			.E(gen[391]),

			.SO(gen[484]),
			.S(gen[485]),
			.SE(gen[486]),

			.SELF(gen[390]),
			.cell_state(gen[390])
		); 

/******************* CELL 391 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell391 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[295]),
			.N(gen[296]),
			.NE(gen[297]),

			.O(gen[390]),
			.E(gen[392]),

			.SO(gen[485]),
			.S(gen[486]),
			.SE(gen[487]),

			.SELF(gen[391]),
			.cell_state(gen[391])
		); 

/******************* CELL 392 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell392 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[296]),
			.N(gen[297]),
			.NE(gen[298]),

			.O(gen[391]),
			.E(gen[393]),

			.SO(gen[486]),
			.S(gen[487]),
			.SE(gen[488]),

			.SELF(gen[392]),
			.cell_state(gen[392])
		); 

/******************* CELL 393 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell393 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[297]),
			.N(gen[298]),
			.NE(gen[299]),

			.O(gen[392]),
			.E(gen[394]),

			.SO(gen[487]),
			.S(gen[488]),
			.SE(gen[489]),

			.SELF(gen[393]),
			.cell_state(gen[393])
		); 

/******************* CELL 394 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell394 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[298]),
			.N(gen[299]),
			.NE(gen[300]),

			.O(gen[393]),
			.E(gen[395]),

			.SO(gen[488]),
			.S(gen[489]),
			.SE(gen[490]),

			.SELF(gen[394]),
			.cell_state(gen[394])
		); 

/******************* CELL 395 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell395 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[299]),
			.N(gen[300]),
			.NE(gen[301]),

			.O(gen[394]),
			.E(gen[396]),

			.SO(gen[489]),
			.S(gen[490]),
			.SE(gen[491]),

			.SELF(gen[395]),
			.cell_state(gen[395])
		); 

/******************* CELL 396 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell396 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[300]),
			.N(gen[301]),
			.NE(gen[302]),

			.O(gen[395]),
			.E(gen[397]),

			.SO(gen[490]),
			.S(gen[491]),
			.SE(gen[492]),

			.SELF(gen[396]),
			.cell_state(gen[396])
		); 

/******************* CELL 397 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell397 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[301]),
			.N(gen[302]),
			.NE(gen[303]),

			.O(gen[396]),
			.E(gen[398]),

			.SO(gen[491]),
			.S(gen[492]),
			.SE(gen[493]),

			.SELF(gen[397]),
			.cell_state(gen[397])
		); 

/******************* CELL 398 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell398 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[302]),
			.N(gen[303]),
			.NE(gen[304]),

			.O(gen[397]),
			.E(gen[399]),

			.SO(gen[492]),
			.S(gen[493]),
			.SE(gen[494]),

			.SELF(gen[398]),
			.cell_state(gen[398])
		); 

/******************* CELL 399 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell399 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[303]),
			.N(gen[304]),
			.NE(gen[305]),

			.O(gen[398]),
			.E(gen[400]),

			.SO(gen[493]),
			.S(gen[494]),
			.SE(gen[495]),

			.SELF(gen[399]),
			.cell_state(gen[399])
		); 

/******************* CELL 400 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell400 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[304]),
			.N(gen[305]),
			.NE(gen[306]),

			.O(gen[399]),
			.E(gen[401]),

			.SO(gen[494]),
			.S(gen[495]),
			.SE(gen[496]),

			.SELF(gen[400]),
			.cell_state(gen[400])
		); 

/******************* CELL 401 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell401 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[305]),
			.N(gen[306]),
			.NE(gen[307]),

			.O(gen[400]),
			.E(gen[402]),

			.SO(gen[495]),
			.S(gen[496]),
			.SE(gen[497]),

			.SELF(gen[401]),
			.cell_state(gen[401])
		); 

/******************* CELL 402 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell402 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[306]),
			.N(gen[307]),
			.NE(gen[308]),

			.O(gen[401]),
			.E(gen[403]),

			.SO(gen[496]),
			.S(gen[497]),
			.SE(gen[498]),

			.SELF(gen[402]),
			.cell_state(gen[402])
		); 

/******************* CELL 403 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell403 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[307]),
			.N(gen[308]),
			.NE(gen[309]),

			.O(gen[402]),
			.E(gen[404]),

			.SO(gen[497]),
			.S(gen[498]),
			.SE(gen[499]),

			.SELF(gen[403]),
			.cell_state(gen[403])
		); 

/******************* CELL 404 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell404 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[308]),
			.N(gen[309]),
			.NE(gen[310]),

			.O(gen[403]),
			.E(gen[405]),

			.SO(gen[498]),
			.S(gen[499]),
			.SE(gen[500]),

			.SELF(gen[404]),
			.cell_state(gen[404])
		); 

/******************* CELL 405 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell405 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[309]),
			.N(gen[310]),
			.NE(gen[311]),

			.O(gen[404]),
			.E(gen[406]),

			.SO(gen[499]),
			.S(gen[500]),
			.SE(gen[501]),

			.SELF(gen[405]),
			.cell_state(gen[405])
		); 

/******************* CELL 406 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell406 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[310]),
			.N(gen[311]),
			.NE(gen[312]),

			.O(gen[405]),
			.E(gen[407]),

			.SO(gen[500]),
			.S(gen[501]),
			.SE(gen[502]),

			.SELF(gen[406]),
			.cell_state(gen[406])
		); 

/******************* CELL 407 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell407 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[311]),
			.N(gen[312]),
			.NE(gen[313]),

			.O(gen[406]),
			.E(gen[408]),

			.SO(gen[501]),
			.S(gen[502]),
			.SE(gen[503]),

			.SELF(gen[407]),
			.cell_state(gen[407])
		); 

/******************* CELL 408 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell408 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[312]),
			.N(gen[313]),
			.NE(gen[314]),

			.O(gen[407]),
			.E(gen[409]),

			.SO(gen[502]),
			.S(gen[503]),
			.SE(gen[504]),

			.SELF(gen[408]),
			.cell_state(gen[408])
		); 

/******************* CELL 409 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell409 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[313]),
			.N(gen[314]),
			.NE(gen[315]),

			.O(gen[408]),
			.E(gen[410]),

			.SO(gen[503]),
			.S(gen[504]),
			.SE(gen[505]),

			.SELF(gen[409]),
			.cell_state(gen[409])
		); 

/******************* CELL 410 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell410 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[314]),
			.N(gen[315]),
			.NE(gen[316]),

			.O(gen[409]),
			.E(gen[411]),

			.SO(gen[504]),
			.S(gen[505]),
			.SE(gen[506]),

			.SELF(gen[410]),
			.cell_state(gen[410])
		); 

/******************* CELL 411 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell411 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[315]),
			.N(gen[316]),
			.NE(gen[317]),

			.O(gen[410]),
			.E(gen[412]),

			.SO(gen[505]),
			.S(gen[506]),
			.SE(gen[507]),

			.SELF(gen[411]),
			.cell_state(gen[411])
		); 

/******************* CELL 412 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell412 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[316]),
			.N(gen[317]),
			.NE(gen[318]),

			.O(gen[411]),
			.E(gen[413]),

			.SO(gen[506]),
			.S(gen[507]),
			.SE(gen[508]),

			.SELF(gen[412]),
			.cell_state(gen[412])
		); 

/******************* CELL 413 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell413 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[317]),
			.N(gen[318]),
			.NE(gen[319]),

			.O(gen[412]),
			.E(gen[414]),

			.SO(gen[507]),
			.S(gen[508]),
			.SE(gen[509]),

			.SELF(gen[413]),
			.cell_state(gen[413])
		); 

/******************* CELL 414 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell414 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[318]),
			.N(gen[319]),
			.NE(gen[320]),

			.O(gen[413]),
			.E(gen[415]),

			.SO(gen[508]),
			.S(gen[509]),
			.SE(gen[510]),

			.SELF(gen[414]),
			.cell_state(gen[414])
		); 

/******************* CELL 415 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell415 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[319]),
			.N(gen[320]),
			.NE(gen[321]),

			.O(gen[414]),
			.E(gen[416]),

			.SO(gen[509]),
			.S(gen[510]),
			.SE(gen[511]),

			.SELF(gen[415]),
			.cell_state(gen[415])
		); 

/******************* CELL 416 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell416 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[320]),
			.N(gen[321]),
			.NE(gen[322]),

			.O(gen[415]),
			.E(gen[417]),

			.SO(gen[510]),
			.S(gen[511]),
			.SE(gen[512]),

			.SELF(gen[416]),
			.cell_state(gen[416])
		); 

/******************* CELL 417 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell417 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[321]),
			.N(gen[322]),
			.NE(gen[323]),

			.O(gen[416]),
			.E(gen[418]),

			.SO(gen[511]),
			.S(gen[512]),
			.SE(gen[513]),

			.SELF(gen[417]),
			.cell_state(gen[417])
		); 

/******************* CELL 418 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell418 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[322]),
			.N(gen[323]),
			.NE(gen[324]),

			.O(gen[417]),
			.E(gen[419]),

			.SO(gen[512]),
			.S(gen[513]),
			.SE(gen[514]),

			.SELF(gen[418]),
			.cell_state(gen[418])
		); 

/******************* CELL 419 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell419 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[323]),
			.N(gen[324]),
			.NE(gen[325]),

			.O(gen[418]),
			.E(gen[420]),

			.SO(gen[513]),
			.S(gen[514]),
			.SE(gen[515]),

			.SELF(gen[419]),
			.cell_state(gen[419])
		); 

/******************* CELL 420 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell420 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[324]),
			.N(gen[325]),
			.NE(gen[326]),

			.O(gen[419]),
			.E(gen[421]),

			.SO(gen[514]),
			.S(gen[515]),
			.SE(gen[516]),

			.SELF(gen[420]),
			.cell_state(gen[420])
		); 

/******************* CELL 421 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell421 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[325]),
			.N(gen[326]),
			.NE(gen[327]),

			.O(gen[420]),
			.E(gen[422]),

			.SO(gen[515]),
			.S(gen[516]),
			.SE(gen[517]),

			.SELF(gen[421]),
			.cell_state(gen[421])
		); 

/******************* CELL 422 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell422 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[326]),
			.N(gen[327]),
			.NE(gen[328]),

			.O(gen[421]),
			.E(gen[423]),

			.SO(gen[516]),
			.S(gen[517]),
			.SE(gen[518]),

			.SELF(gen[422]),
			.cell_state(gen[422])
		); 

/******************* CELL 423 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell423 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[327]),
			.N(gen[328]),
			.NE(gen[329]),

			.O(gen[422]),
			.E(gen[424]),

			.SO(gen[517]),
			.S(gen[518]),
			.SE(gen[519]),

			.SELF(gen[423]),
			.cell_state(gen[423])
		); 

/******************* CELL 424 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell424 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[328]),
			.N(gen[329]),
			.NE(gen[330]),

			.O(gen[423]),
			.E(gen[425]),

			.SO(gen[518]),
			.S(gen[519]),
			.SE(gen[520]),

			.SELF(gen[424]),
			.cell_state(gen[424])
		); 

/******************* CELL 425 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell425 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[329]),
			.N(gen[330]),
			.NE(gen[331]),

			.O(gen[424]),
			.E(gen[426]),

			.SO(gen[519]),
			.S(gen[520]),
			.SE(gen[521]),

			.SELF(gen[425]),
			.cell_state(gen[425])
		); 

/******************* CELL 426 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell426 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[330]),
			.N(gen[331]),
			.NE(gen[332]),

			.O(gen[425]),
			.E(gen[427]),

			.SO(gen[520]),
			.S(gen[521]),
			.SE(gen[522]),

			.SELF(gen[426]),
			.cell_state(gen[426])
		); 

/******************* CELL 427 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell427 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[331]),
			.N(gen[332]),
			.NE(gen[333]),

			.O(gen[426]),
			.E(gen[428]),

			.SO(gen[521]),
			.S(gen[522]),
			.SE(gen[523]),

			.SELF(gen[427]),
			.cell_state(gen[427])
		); 

/******************* CELL 428 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell428 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[332]),
			.N(gen[333]),
			.NE(gen[334]),

			.O(gen[427]),
			.E(gen[429]),

			.SO(gen[522]),
			.S(gen[523]),
			.SE(gen[524]),

			.SELF(gen[428]),
			.cell_state(gen[428])
		); 

/******************* CELL 429 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell429 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[333]),
			.N(gen[334]),
			.NE(gen[335]),

			.O(gen[428]),
			.E(gen[430]),

			.SO(gen[523]),
			.S(gen[524]),
			.SE(gen[525]),

			.SELF(gen[429]),
			.cell_state(gen[429])
		); 

/******************* CELL 430 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell430 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[334]),
			.N(gen[335]),
			.NE(gen[336]),

			.O(gen[429]),
			.E(gen[431]),

			.SO(gen[524]),
			.S(gen[525]),
			.SE(gen[526]),

			.SELF(gen[430]),
			.cell_state(gen[430])
		); 

/******************* CELL 431 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell431 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[335]),
			.N(gen[336]),
			.NE(gen[337]),

			.O(gen[430]),
			.E(gen[432]),

			.SO(gen[525]),
			.S(gen[526]),
			.SE(gen[527]),

			.SELF(gen[431]),
			.cell_state(gen[431])
		); 

/******************* CELL 432 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell432 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[336]),
			.N(gen[337]),
			.NE(gen[338]),

			.O(gen[431]),
			.E(gen[433]),

			.SO(gen[526]),
			.S(gen[527]),
			.SE(gen[528]),

			.SELF(gen[432]),
			.cell_state(gen[432])
		); 

/******************* CELL 433 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell433 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[337]),
			.N(gen[338]),
			.NE(gen[339]),

			.O(gen[432]),
			.E(gen[434]),

			.SO(gen[527]),
			.S(gen[528]),
			.SE(gen[529]),

			.SELF(gen[433]),
			.cell_state(gen[433])
		); 

/******************* CELL 434 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell434 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[338]),
			.N(gen[339]),
			.NE(gen[340]),

			.O(gen[433]),
			.E(gen[435]),

			.SO(gen[528]),
			.S(gen[529]),
			.SE(gen[530]),

			.SELF(gen[434]),
			.cell_state(gen[434])
		); 

/******************* CELL 435 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell435 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[339]),
			.N(gen[340]),
			.NE(gen[341]),

			.O(gen[434]),
			.E(gen[436]),

			.SO(gen[529]),
			.S(gen[530]),
			.SE(gen[531]),

			.SELF(gen[435]),
			.cell_state(gen[435])
		); 

/******************* CELL 436 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell436 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[340]),
			.N(gen[341]),
			.NE(gen[342]),

			.O(gen[435]),
			.E(gen[437]),

			.SO(gen[530]),
			.S(gen[531]),
			.SE(gen[532]),

			.SELF(gen[436]),
			.cell_state(gen[436])
		); 

/******************* CELL 437 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell437 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[341]),
			.N(gen[342]),
			.NE(gen[343]),

			.O(gen[436]),
			.E(gen[438]),

			.SO(gen[531]),
			.S(gen[532]),
			.SE(gen[533]),

			.SELF(gen[437]),
			.cell_state(gen[437])
		); 

/******************* CELL 438 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell438 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[342]),
			.N(gen[343]),
			.NE(gen[344]),

			.O(gen[437]),
			.E(gen[439]),

			.SO(gen[532]),
			.S(gen[533]),
			.SE(gen[534]),

			.SELF(gen[438]),
			.cell_state(gen[438])
		); 

/******************* CELL 439 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell439 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[343]),
			.N(gen[344]),
			.NE(gen[345]),

			.O(gen[438]),
			.E(gen[440]),

			.SO(gen[533]),
			.S(gen[534]),
			.SE(gen[535]),

			.SELF(gen[439]),
			.cell_state(gen[439])
		); 

/******************* CELL 440 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell440 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[344]),
			.N(gen[345]),
			.NE(gen[346]),

			.O(gen[439]),
			.E(gen[441]),

			.SO(gen[534]),
			.S(gen[535]),
			.SE(gen[536]),

			.SELF(gen[440]),
			.cell_state(gen[440])
		); 

/******************* CELL 441 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell441 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[345]),
			.N(gen[346]),
			.NE(gen[347]),

			.O(gen[440]),
			.E(gen[442]),

			.SO(gen[535]),
			.S(gen[536]),
			.SE(gen[537]),

			.SELF(gen[441]),
			.cell_state(gen[441])
		); 

/******************* CELL 442 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell442 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[346]),
			.N(gen[347]),
			.NE(gen[348]),

			.O(gen[441]),
			.E(gen[443]),

			.SO(gen[536]),
			.S(gen[537]),
			.SE(gen[538]),

			.SELF(gen[442]),
			.cell_state(gen[442])
		); 

/******************* CELL 443 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell443 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[347]),
			.N(gen[348]),
			.NE(gen[349]),

			.O(gen[442]),
			.E(gen[444]),

			.SO(gen[537]),
			.S(gen[538]),
			.SE(gen[539]),

			.SELF(gen[443]),
			.cell_state(gen[443])
		); 

/******************* CELL 444 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell444 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[348]),
			.N(gen[349]),
			.NE(gen[350]),

			.O(gen[443]),
			.E(gen[445]),

			.SO(gen[538]),
			.S(gen[539]),
			.SE(gen[540]),

			.SELF(gen[444]),
			.cell_state(gen[444])
		); 

/******************* CELL 445 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell445 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[349]),
			.N(gen[350]),
			.NE(gen[351]),

			.O(gen[444]),
			.E(gen[446]),

			.SO(gen[539]),
			.S(gen[540]),
			.SE(gen[541]),

			.SELF(gen[445]),
			.cell_state(gen[445])
		); 

/******************* CELL 446 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell446 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[350]),
			.N(gen[351]),
			.NE(gen[352]),

			.O(gen[445]),
			.E(gen[447]),

			.SO(gen[540]),
			.S(gen[541]),
			.SE(gen[542]),

			.SELF(gen[446]),
			.cell_state(gen[446])
		); 

/******************* CELL 447 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell447 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[351]),
			.N(gen[352]),
			.NE(gen[353]),

			.O(gen[446]),
			.E(gen[448]),

			.SO(gen[541]),
			.S(gen[542]),
			.SE(gen[543]),

			.SELF(gen[447]),
			.cell_state(gen[447])
		); 

/******************* CELL 448 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell448 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[352]),
			.N(gen[353]),
			.NE(gen[354]),

			.O(gen[447]),
			.E(gen[449]),

			.SO(gen[542]),
			.S(gen[543]),
			.SE(gen[544]),

			.SELF(gen[448]),
			.cell_state(gen[448])
		); 

/******************* CELL 449 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell449 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[353]),
			.N(gen[354]),
			.NE(gen[355]),

			.O(gen[448]),
			.E(gen[450]),

			.SO(gen[543]),
			.S(gen[544]),
			.SE(gen[545]),

			.SELF(gen[449]),
			.cell_state(gen[449])
		); 

/******************* CELL 450 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell450 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[354]),
			.N(gen[355]),
			.NE(gen[356]),

			.O(gen[449]),
			.E(gen[451]),

			.SO(gen[544]),
			.S(gen[545]),
			.SE(gen[546]),

			.SELF(gen[450]),
			.cell_state(gen[450])
		); 

/******************* CELL 451 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell451 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[355]),
			.N(gen[356]),
			.NE(gen[357]),

			.O(gen[450]),
			.E(gen[452]),

			.SO(gen[545]),
			.S(gen[546]),
			.SE(gen[547]),

			.SELF(gen[451]),
			.cell_state(gen[451])
		); 

/******************* CELL 452 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell452 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[356]),
			.N(gen[357]),
			.NE(gen[358]),

			.O(gen[451]),
			.E(gen[453]),

			.SO(gen[546]),
			.S(gen[547]),
			.SE(gen[548]),

			.SELF(gen[452]),
			.cell_state(gen[452])
		); 

/******************* CELL 453 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell453 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[357]),
			.N(gen[358]),
			.NE(gen[359]),

			.O(gen[452]),
			.E(gen[454]),

			.SO(gen[547]),
			.S(gen[548]),
			.SE(gen[549]),

			.SELF(gen[453]),
			.cell_state(gen[453])
		); 

/******************* CELL 454 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell454 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[358]),
			.N(gen[359]),
			.NE(gen[360]),

			.O(gen[453]),
			.E(gen[455]),

			.SO(gen[548]),
			.S(gen[549]),
			.SE(gen[550]),

			.SELF(gen[454]),
			.cell_state(gen[454])
		); 

/******************* CELL 455 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell455 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[359]),
			.N(gen[360]),
			.NE(gen[361]),

			.O(gen[454]),
			.E(gen[456]),

			.SO(gen[549]),
			.S(gen[550]),
			.SE(gen[551]),

			.SELF(gen[455]),
			.cell_state(gen[455])
		); 

/******************* CELL 456 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell456 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[360]),
			.N(gen[361]),
			.NE(gen[362]),

			.O(gen[455]),
			.E(gen[457]),

			.SO(gen[550]),
			.S(gen[551]),
			.SE(gen[552]),

			.SELF(gen[456]),
			.cell_state(gen[456])
		); 

/******************* CELL 457 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell457 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[361]),
			.N(gen[362]),
			.NE(gen[363]),

			.O(gen[456]),
			.E(gen[458]),

			.SO(gen[551]),
			.S(gen[552]),
			.SE(gen[553]),

			.SELF(gen[457]),
			.cell_state(gen[457])
		); 

/******************* CELL 458 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell458 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[362]),
			.N(gen[363]),
			.NE(gen[364]),

			.O(gen[457]),
			.E(gen[459]),

			.SO(gen[552]),
			.S(gen[553]),
			.SE(gen[554]),

			.SELF(gen[458]),
			.cell_state(gen[458])
		); 

/******************* CELL 459 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell459 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[363]),
			.N(gen[364]),
			.NE(gen[365]),

			.O(gen[458]),
			.E(gen[460]),

			.SO(gen[553]),
			.S(gen[554]),
			.SE(gen[555]),

			.SELF(gen[459]),
			.cell_state(gen[459])
		); 

/******************* CELL 460 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell460 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[364]),
			.N(gen[365]),
			.NE(gen[366]),

			.O(gen[459]),
			.E(gen[461]),

			.SO(gen[554]),
			.S(gen[555]),
			.SE(gen[556]),

			.SELF(gen[460]),
			.cell_state(gen[460])
		); 

/******************* CELL 461 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell461 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[365]),
			.N(gen[366]),
			.NE(gen[367]),

			.O(gen[460]),
			.E(gen[462]),

			.SO(gen[555]),
			.S(gen[556]),
			.SE(gen[557]),

			.SELF(gen[461]),
			.cell_state(gen[461])
		); 

/******************* CELL 462 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell462 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[366]),
			.N(gen[367]),
			.NE(gen[368]),

			.O(gen[461]),
			.E(gen[463]),

			.SO(gen[556]),
			.S(gen[557]),
			.SE(gen[558]),

			.SELF(gen[462]),
			.cell_state(gen[462])
		); 

/******************* CELL 463 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell463 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[367]),
			.N(gen[368]),
			.NE(gen[369]),

			.O(gen[462]),
			.E(gen[464]),

			.SO(gen[557]),
			.S(gen[558]),
			.SE(gen[559]),

			.SELF(gen[463]),
			.cell_state(gen[463])
		); 

/******************* CELL 464 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell464 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[368]),
			.N(gen[369]),
			.NE(gen[370]),

			.O(gen[463]),
			.E(gen[465]),

			.SO(gen[558]),
			.S(gen[559]),
			.SE(gen[560]),

			.SELF(gen[464]),
			.cell_state(gen[464])
		); 

/******************* CELL 465 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell465 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[369]),
			.N(gen[370]),
			.NE(gen[371]),

			.O(gen[464]),
			.E(gen[466]),

			.SO(gen[559]),
			.S(gen[560]),
			.SE(gen[561]),

			.SELF(gen[465]),
			.cell_state(gen[465])
		); 

/******************* CELL 466 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell466 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[370]),
			.N(gen[371]),
			.NE(gen[372]),

			.O(gen[465]),
			.E(gen[467]),

			.SO(gen[560]),
			.S(gen[561]),
			.SE(gen[562]),

			.SELF(gen[466]),
			.cell_state(gen[466])
		); 

/******************* CELL 467 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell467 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[371]),
			.N(gen[372]),
			.NE(gen[373]),

			.O(gen[466]),
			.E(gen[468]),

			.SO(gen[561]),
			.S(gen[562]),
			.SE(gen[563]),

			.SELF(gen[467]),
			.cell_state(gen[467])
		); 

/******************* CELL 468 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell468 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[372]),
			.N(gen[373]),
			.NE(gen[374]),

			.O(gen[467]),
			.E(gen[469]),

			.SO(gen[562]),
			.S(gen[563]),
			.SE(gen[564]),

			.SELF(gen[468]),
			.cell_state(gen[468])
		); 

/******************* CELL 469 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell469 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[373]),
			.N(gen[374]),
			.NE(gen[375]),

			.O(gen[468]),
			.E(gen[470]),

			.SO(gen[563]),
			.S(gen[564]),
			.SE(gen[565]),

			.SELF(gen[469]),
			.cell_state(gen[469])
		); 

/******************* CELL 470 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell470 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[374]),
			.N(gen[375]),
			.NE(gen[376]),

			.O(gen[469]),
			.E(gen[471]),

			.SO(gen[564]),
			.S(gen[565]),
			.SE(gen[566]),

			.SELF(gen[470]),
			.cell_state(gen[470])
		); 

/******************* CELL 471 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell471 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[375]),
			.N(gen[376]),
			.NE(gen[377]),

			.O(gen[470]),
			.E(gen[472]),

			.SO(gen[565]),
			.S(gen[566]),
			.SE(gen[567]),

			.SELF(gen[471]),
			.cell_state(gen[471])
		); 

/******************* CELL 472 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell472 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[376]),
			.N(gen[377]),
			.NE(gen[378]),

			.O(gen[471]),
			.E(gen[473]),

			.SO(gen[566]),
			.S(gen[567]),
			.SE(gen[568]),

			.SELF(gen[472]),
			.cell_state(gen[472])
		); 

/******************* CELL 473 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell473 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[377]),
			.N(gen[378]),
			.NE(gen[379]),

			.O(gen[472]),
			.E(gen[474]),

			.SO(gen[567]),
			.S(gen[568]),
			.SE(gen[569]),

			.SELF(gen[473]),
			.cell_state(gen[473])
		); 

/******************* CELL 474 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell474 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[378]),
			.N(gen[379]),
			.NE(gen[378]),

			.O(gen[473]),
			.E(gen[473]),

			.SO(gen[568]),
			.S(gen[569]),
			.SE(gen[568]),

			.SELF(gen[474]),
			.cell_state(gen[474])
		); 

/******************* CELL 475 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell475 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[381]),
			.N(gen[380]),
			.NE(gen[381]),

			.O(gen[476]),
			.E(gen[476]),

			.SO(gen[571]),
			.S(gen[570]),
			.SE(gen[571]),

			.SELF(gen[475]),
			.cell_state(gen[475])
		); 

/******************* CELL 476 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell476 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[380]),
			.N(gen[381]),
			.NE(gen[382]),

			.O(gen[475]),
			.E(gen[477]),

			.SO(gen[570]),
			.S(gen[571]),
			.SE(gen[572]),

			.SELF(gen[476]),
			.cell_state(gen[476])
		); 

/******************* CELL 477 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell477 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[381]),
			.N(gen[382]),
			.NE(gen[383]),

			.O(gen[476]),
			.E(gen[478]),

			.SO(gen[571]),
			.S(gen[572]),
			.SE(gen[573]),

			.SELF(gen[477]),
			.cell_state(gen[477])
		); 

/******************* CELL 478 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell478 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[382]),
			.N(gen[383]),
			.NE(gen[384]),

			.O(gen[477]),
			.E(gen[479]),

			.SO(gen[572]),
			.S(gen[573]),
			.SE(gen[574]),

			.SELF(gen[478]),
			.cell_state(gen[478])
		); 

/******************* CELL 479 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell479 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[383]),
			.N(gen[384]),
			.NE(gen[385]),

			.O(gen[478]),
			.E(gen[480]),

			.SO(gen[573]),
			.S(gen[574]),
			.SE(gen[575]),

			.SELF(gen[479]),
			.cell_state(gen[479])
		); 

/******************* CELL 480 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell480 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[384]),
			.N(gen[385]),
			.NE(gen[386]),

			.O(gen[479]),
			.E(gen[481]),

			.SO(gen[574]),
			.S(gen[575]),
			.SE(gen[576]),

			.SELF(gen[480]),
			.cell_state(gen[480])
		); 

/******************* CELL 481 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell481 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[385]),
			.N(gen[386]),
			.NE(gen[387]),

			.O(gen[480]),
			.E(gen[482]),

			.SO(gen[575]),
			.S(gen[576]),
			.SE(gen[577]),

			.SELF(gen[481]),
			.cell_state(gen[481])
		); 

/******************* CELL 482 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell482 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[386]),
			.N(gen[387]),
			.NE(gen[388]),

			.O(gen[481]),
			.E(gen[483]),

			.SO(gen[576]),
			.S(gen[577]),
			.SE(gen[578]),

			.SELF(gen[482]),
			.cell_state(gen[482])
		); 

/******************* CELL 483 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell483 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[387]),
			.N(gen[388]),
			.NE(gen[389]),

			.O(gen[482]),
			.E(gen[484]),

			.SO(gen[577]),
			.S(gen[578]),
			.SE(gen[579]),

			.SELF(gen[483]),
			.cell_state(gen[483])
		); 

/******************* CELL 484 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell484 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[388]),
			.N(gen[389]),
			.NE(gen[390]),

			.O(gen[483]),
			.E(gen[485]),

			.SO(gen[578]),
			.S(gen[579]),
			.SE(gen[580]),

			.SELF(gen[484]),
			.cell_state(gen[484])
		); 

/******************* CELL 485 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell485 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[389]),
			.N(gen[390]),
			.NE(gen[391]),

			.O(gen[484]),
			.E(gen[486]),

			.SO(gen[579]),
			.S(gen[580]),
			.SE(gen[581]),

			.SELF(gen[485]),
			.cell_state(gen[485])
		); 

/******************* CELL 486 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell486 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[390]),
			.N(gen[391]),
			.NE(gen[392]),

			.O(gen[485]),
			.E(gen[487]),

			.SO(gen[580]),
			.S(gen[581]),
			.SE(gen[582]),

			.SELF(gen[486]),
			.cell_state(gen[486])
		); 

/******************* CELL 487 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell487 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[391]),
			.N(gen[392]),
			.NE(gen[393]),

			.O(gen[486]),
			.E(gen[488]),

			.SO(gen[581]),
			.S(gen[582]),
			.SE(gen[583]),

			.SELF(gen[487]),
			.cell_state(gen[487])
		); 

/******************* CELL 488 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell488 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[392]),
			.N(gen[393]),
			.NE(gen[394]),

			.O(gen[487]),
			.E(gen[489]),

			.SO(gen[582]),
			.S(gen[583]),
			.SE(gen[584]),

			.SELF(gen[488]),
			.cell_state(gen[488])
		); 

/******************* CELL 489 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell489 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[393]),
			.N(gen[394]),
			.NE(gen[395]),

			.O(gen[488]),
			.E(gen[490]),

			.SO(gen[583]),
			.S(gen[584]),
			.SE(gen[585]),

			.SELF(gen[489]),
			.cell_state(gen[489])
		); 

/******************* CELL 490 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell490 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[394]),
			.N(gen[395]),
			.NE(gen[396]),

			.O(gen[489]),
			.E(gen[491]),

			.SO(gen[584]),
			.S(gen[585]),
			.SE(gen[586]),

			.SELF(gen[490]),
			.cell_state(gen[490])
		); 

/******************* CELL 491 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell491 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[395]),
			.N(gen[396]),
			.NE(gen[397]),

			.O(gen[490]),
			.E(gen[492]),

			.SO(gen[585]),
			.S(gen[586]),
			.SE(gen[587]),

			.SELF(gen[491]),
			.cell_state(gen[491])
		); 

/******************* CELL 492 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell492 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[396]),
			.N(gen[397]),
			.NE(gen[398]),

			.O(gen[491]),
			.E(gen[493]),

			.SO(gen[586]),
			.S(gen[587]),
			.SE(gen[588]),

			.SELF(gen[492]),
			.cell_state(gen[492])
		); 

/******************* CELL 493 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell493 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[397]),
			.N(gen[398]),
			.NE(gen[399]),

			.O(gen[492]),
			.E(gen[494]),

			.SO(gen[587]),
			.S(gen[588]),
			.SE(gen[589]),

			.SELF(gen[493]),
			.cell_state(gen[493])
		); 

/******************* CELL 494 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell494 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[398]),
			.N(gen[399]),
			.NE(gen[400]),

			.O(gen[493]),
			.E(gen[495]),

			.SO(gen[588]),
			.S(gen[589]),
			.SE(gen[590]),

			.SELF(gen[494]),
			.cell_state(gen[494])
		); 

/******************* CELL 495 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell495 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[399]),
			.N(gen[400]),
			.NE(gen[401]),

			.O(gen[494]),
			.E(gen[496]),

			.SO(gen[589]),
			.S(gen[590]),
			.SE(gen[591]),

			.SELF(gen[495]),
			.cell_state(gen[495])
		); 

/******************* CELL 496 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell496 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[400]),
			.N(gen[401]),
			.NE(gen[402]),

			.O(gen[495]),
			.E(gen[497]),

			.SO(gen[590]),
			.S(gen[591]),
			.SE(gen[592]),

			.SELF(gen[496]),
			.cell_state(gen[496])
		); 

/******************* CELL 497 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell497 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[401]),
			.N(gen[402]),
			.NE(gen[403]),

			.O(gen[496]),
			.E(gen[498]),

			.SO(gen[591]),
			.S(gen[592]),
			.SE(gen[593]),

			.SELF(gen[497]),
			.cell_state(gen[497])
		); 

/******************* CELL 498 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell498 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[402]),
			.N(gen[403]),
			.NE(gen[404]),

			.O(gen[497]),
			.E(gen[499]),

			.SO(gen[592]),
			.S(gen[593]),
			.SE(gen[594]),

			.SELF(gen[498]),
			.cell_state(gen[498])
		); 

/******************* CELL 499 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell499 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[403]),
			.N(gen[404]),
			.NE(gen[405]),

			.O(gen[498]),
			.E(gen[500]),

			.SO(gen[593]),
			.S(gen[594]),
			.SE(gen[595]),

			.SELF(gen[499]),
			.cell_state(gen[499])
		); 

/******************* CELL 500 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell500 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[404]),
			.N(gen[405]),
			.NE(gen[406]),

			.O(gen[499]),
			.E(gen[501]),

			.SO(gen[594]),
			.S(gen[595]),
			.SE(gen[596]),

			.SELF(gen[500]),
			.cell_state(gen[500])
		); 

/******************* CELL 501 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell501 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[405]),
			.N(gen[406]),
			.NE(gen[407]),

			.O(gen[500]),
			.E(gen[502]),

			.SO(gen[595]),
			.S(gen[596]),
			.SE(gen[597]),

			.SELF(gen[501]),
			.cell_state(gen[501])
		); 

/******************* CELL 502 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell502 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[406]),
			.N(gen[407]),
			.NE(gen[408]),

			.O(gen[501]),
			.E(gen[503]),

			.SO(gen[596]),
			.S(gen[597]),
			.SE(gen[598]),

			.SELF(gen[502]),
			.cell_state(gen[502])
		); 

/******************* CELL 503 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell503 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[407]),
			.N(gen[408]),
			.NE(gen[409]),

			.O(gen[502]),
			.E(gen[504]),

			.SO(gen[597]),
			.S(gen[598]),
			.SE(gen[599]),

			.SELF(gen[503]),
			.cell_state(gen[503])
		); 

/******************* CELL 504 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell504 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[408]),
			.N(gen[409]),
			.NE(gen[410]),

			.O(gen[503]),
			.E(gen[505]),

			.SO(gen[598]),
			.S(gen[599]),
			.SE(gen[600]),

			.SELF(gen[504]),
			.cell_state(gen[504])
		); 

/******************* CELL 505 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell505 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[409]),
			.N(gen[410]),
			.NE(gen[411]),

			.O(gen[504]),
			.E(gen[506]),

			.SO(gen[599]),
			.S(gen[600]),
			.SE(gen[601]),

			.SELF(gen[505]),
			.cell_state(gen[505])
		); 

/******************* CELL 506 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell506 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[410]),
			.N(gen[411]),
			.NE(gen[412]),

			.O(gen[505]),
			.E(gen[507]),

			.SO(gen[600]),
			.S(gen[601]),
			.SE(gen[602]),

			.SELF(gen[506]),
			.cell_state(gen[506])
		); 

/******************* CELL 507 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell507 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[411]),
			.N(gen[412]),
			.NE(gen[413]),

			.O(gen[506]),
			.E(gen[508]),

			.SO(gen[601]),
			.S(gen[602]),
			.SE(gen[603]),

			.SELF(gen[507]),
			.cell_state(gen[507])
		); 

/******************* CELL 508 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell508 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[412]),
			.N(gen[413]),
			.NE(gen[414]),

			.O(gen[507]),
			.E(gen[509]),

			.SO(gen[602]),
			.S(gen[603]),
			.SE(gen[604]),

			.SELF(gen[508]),
			.cell_state(gen[508])
		); 

/******************* CELL 509 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell509 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[413]),
			.N(gen[414]),
			.NE(gen[415]),

			.O(gen[508]),
			.E(gen[510]),

			.SO(gen[603]),
			.S(gen[604]),
			.SE(gen[605]),

			.SELF(gen[509]),
			.cell_state(gen[509])
		); 

/******************* CELL 510 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell510 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[414]),
			.N(gen[415]),
			.NE(gen[416]),

			.O(gen[509]),
			.E(gen[511]),

			.SO(gen[604]),
			.S(gen[605]),
			.SE(gen[606]),

			.SELF(gen[510]),
			.cell_state(gen[510])
		); 

/******************* CELL 511 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell511 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[415]),
			.N(gen[416]),
			.NE(gen[417]),

			.O(gen[510]),
			.E(gen[512]),

			.SO(gen[605]),
			.S(gen[606]),
			.SE(gen[607]),

			.SELF(gen[511]),
			.cell_state(gen[511])
		); 

/******************* CELL 512 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell512 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[416]),
			.N(gen[417]),
			.NE(gen[418]),

			.O(gen[511]),
			.E(gen[513]),

			.SO(gen[606]),
			.S(gen[607]),
			.SE(gen[608]),

			.SELF(gen[512]),
			.cell_state(gen[512])
		); 

/******************* CELL 513 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell513 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[417]),
			.N(gen[418]),
			.NE(gen[419]),

			.O(gen[512]),
			.E(gen[514]),

			.SO(gen[607]),
			.S(gen[608]),
			.SE(gen[609]),

			.SELF(gen[513]),
			.cell_state(gen[513])
		); 

/******************* CELL 514 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell514 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[418]),
			.N(gen[419]),
			.NE(gen[420]),

			.O(gen[513]),
			.E(gen[515]),

			.SO(gen[608]),
			.S(gen[609]),
			.SE(gen[610]),

			.SELF(gen[514]),
			.cell_state(gen[514])
		); 

/******************* CELL 515 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell515 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[419]),
			.N(gen[420]),
			.NE(gen[421]),

			.O(gen[514]),
			.E(gen[516]),

			.SO(gen[609]),
			.S(gen[610]),
			.SE(gen[611]),

			.SELF(gen[515]),
			.cell_state(gen[515])
		); 

/******************* CELL 516 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell516 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[420]),
			.N(gen[421]),
			.NE(gen[422]),

			.O(gen[515]),
			.E(gen[517]),

			.SO(gen[610]),
			.S(gen[611]),
			.SE(gen[612]),

			.SELF(gen[516]),
			.cell_state(gen[516])
		); 

/******************* CELL 517 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell517 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[421]),
			.N(gen[422]),
			.NE(gen[423]),

			.O(gen[516]),
			.E(gen[518]),

			.SO(gen[611]),
			.S(gen[612]),
			.SE(gen[613]),

			.SELF(gen[517]),
			.cell_state(gen[517])
		); 

/******************* CELL 518 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell518 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[422]),
			.N(gen[423]),
			.NE(gen[424]),

			.O(gen[517]),
			.E(gen[519]),

			.SO(gen[612]),
			.S(gen[613]),
			.SE(gen[614]),

			.SELF(gen[518]),
			.cell_state(gen[518])
		); 

/******************* CELL 519 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell519 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[423]),
			.N(gen[424]),
			.NE(gen[425]),

			.O(gen[518]),
			.E(gen[520]),

			.SO(gen[613]),
			.S(gen[614]),
			.SE(gen[615]),

			.SELF(gen[519]),
			.cell_state(gen[519])
		); 

/******************* CELL 520 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell520 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[424]),
			.N(gen[425]),
			.NE(gen[426]),

			.O(gen[519]),
			.E(gen[521]),

			.SO(gen[614]),
			.S(gen[615]),
			.SE(gen[616]),

			.SELF(gen[520]),
			.cell_state(gen[520])
		); 

/******************* CELL 521 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell521 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[425]),
			.N(gen[426]),
			.NE(gen[427]),

			.O(gen[520]),
			.E(gen[522]),

			.SO(gen[615]),
			.S(gen[616]),
			.SE(gen[617]),

			.SELF(gen[521]),
			.cell_state(gen[521])
		); 

/******************* CELL 522 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell522 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[426]),
			.N(gen[427]),
			.NE(gen[428]),

			.O(gen[521]),
			.E(gen[523]),

			.SO(gen[616]),
			.S(gen[617]),
			.SE(gen[618]),

			.SELF(gen[522]),
			.cell_state(gen[522])
		); 

/******************* CELL 523 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell523 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[427]),
			.N(gen[428]),
			.NE(gen[429]),

			.O(gen[522]),
			.E(gen[524]),

			.SO(gen[617]),
			.S(gen[618]),
			.SE(gen[619]),

			.SELF(gen[523]),
			.cell_state(gen[523])
		); 

/******************* CELL 524 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell524 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[428]),
			.N(gen[429]),
			.NE(gen[430]),

			.O(gen[523]),
			.E(gen[525]),

			.SO(gen[618]),
			.S(gen[619]),
			.SE(gen[620]),

			.SELF(gen[524]),
			.cell_state(gen[524])
		); 

/******************* CELL 525 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell525 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[429]),
			.N(gen[430]),
			.NE(gen[431]),

			.O(gen[524]),
			.E(gen[526]),

			.SO(gen[619]),
			.S(gen[620]),
			.SE(gen[621]),

			.SELF(gen[525]),
			.cell_state(gen[525])
		); 

/******************* CELL 526 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell526 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[430]),
			.N(gen[431]),
			.NE(gen[432]),

			.O(gen[525]),
			.E(gen[527]),

			.SO(gen[620]),
			.S(gen[621]),
			.SE(gen[622]),

			.SELF(gen[526]),
			.cell_state(gen[526])
		); 

/******************* CELL 527 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell527 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[431]),
			.N(gen[432]),
			.NE(gen[433]),

			.O(gen[526]),
			.E(gen[528]),

			.SO(gen[621]),
			.S(gen[622]),
			.SE(gen[623]),

			.SELF(gen[527]),
			.cell_state(gen[527])
		); 

/******************* CELL 528 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell528 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[432]),
			.N(gen[433]),
			.NE(gen[434]),

			.O(gen[527]),
			.E(gen[529]),

			.SO(gen[622]),
			.S(gen[623]),
			.SE(gen[624]),

			.SELF(gen[528]),
			.cell_state(gen[528])
		); 

/******************* CELL 529 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell529 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[433]),
			.N(gen[434]),
			.NE(gen[435]),

			.O(gen[528]),
			.E(gen[530]),

			.SO(gen[623]),
			.S(gen[624]),
			.SE(gen[625]),

			.SELF(gen[529]),
			.cell_state(gen[529])
		); 

/******************* CELL 530 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell530 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[434]),
			.N(gen[435]),
			.NE(gen[436]),

			.O(gen[529]),
			.E(gen[531]),

			.SO(gen[624]),
			.S(gen[625]),
			.SE(gen[626]),

			.SELF(gen[530]),
			.cell_state(gen[530])
		); 

/******************* CELL 531 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell531 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[435]),
			.N(gen[436]),
			.NE(gen[437]),

			.O(gen[530]),
			.E(gen[532]),

			.SO(gen[625]),
			.S(gen[626]),
			.SE(gen[627]),

			.SELF(gen[531]),
			.cell_state(gen[531])
		); 

/******************* CELL 532 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell532 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[436]),
			.N(gen[437]),
			.NE(gen[438]),

			.O(gen[531]),
			.E(gen[533]),

			.SO(gen[626]),
			.S(gen[627]),
			.SE(gen[628]),

			.SELF(gen[532]),
			.cell_state(gen[532])
		); 

/******************* CELL 533 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell533 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[437]),
			.N(gen[438]),
			.NE(gen[439]),

			.O(gen[532]),
			.E(gen[534]),

			.SO(gen[627]),
			.S(gen[628]),
			.SE(gen[629]),

			.SELF(gen[533]),
			.cell_state(gen[533])
		); 

/******************* CELL 534 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell534 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[438]),
			.N(gen[439]),
			.NE(gen[440]),

			.O(gen[533]),
			.E(gen[535]),

			.SO(gen[628]),
			.S(gen[629]),
			.SE(gen[630]),

			.SELF(gen[534]),
			.cell_state(gen[534])
		); 

/******************* CELL 535 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell535 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[439]),
			.N(gen[440]),
			.NE(gen[441]),

			.O(gen[534]),
			.E(gen[536]),

			.SO(gen[629]),
			.S(gen[630]),
			.SE(gen[631]),

			.SELF(gen[535]),
			.cell_state(gen[535])
		); 

/******************* CELL 536 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell536 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[440]),
			.N(gen[441]),
			.NE(gen[442]),

			.O(gen[535]),
			.E(gen[537]),

			.SO(gen[630]),
			.S(gen[631]),
			.SE(gen[632]),

			.SELF(gen[536]),
			.cell_state(gen[536])
		); 

/******************* CELL 537 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell537 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[441]),
			.N(gen[442]),
			.NE(gen[443]),

			.O(gen[536]),
			.E(gen[538]),

			.SO(gen[631]),
			.S(gen[632]),
			.SE(gen[633]),

			.SELF(gen[537]),
			.cell_state(gen[537])
		); 

/******************* CELL 538 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell538 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[442]),
			.N(gen[443]),
			.NE(gen[444]),

			.O(gen[537]),
			.E(gen[539]),

			.SO(gen[632]),
			.S(gen[633]),
			.SE(gen[634]),

			.SELF(gen[538]),
			.cell_state(gen[538])
		); 

/******************* CELL 539 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell539 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[443]),
			.N(gen[444]),
			.NE(gen[445]),

			.O(gen[538]),
			.E(gen[540]),

			.SO(gen[633]),
			.S(gen[634]),
			.SE(gen[635]),

			.SELF(gen[539]),
			.cell_state(gen[539])
		); 

/******************* CELL 540 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell540 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[444]),
			.N(gen[445]),
			.NE(gen[446]),

			.O(gen[539]),
			.E(gen[541]),

			.SO(gen[634]),
			.S(gen[635]),
			.SE(gen[636]),

			.SELF(gen[540]),
			.cell_state(gen[540])
		); 

/******************* CELL 541 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell541 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[445]),
			.N(gen[446]),
			.NE(gen[447]),

			.O(gen[540]),
			.E(gen[542]),

			.SO(gen[635]),
			.S(gen[636]),
			.SE(gen[637]),

			.SELF(gen[541]),
			.cell_state(gen[541])
		); 

/******************* CELL 542 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell542 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[446]),
			.N(gen[447]),
			.NE(gen[448]),

			.O(gen[541]),
			.E(gen[543]),

			.SO(gen[636]),
			.S(gen[637]),
			.SE(gen[638]),

			.SELF(gen[542]),
			.cell_state(gen[542])
		); 

/******************* CELL 543 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell543 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[447]),
			.N(gen[448]),
			.NE(gen[449]),

			.O(gen[542]),
			.E(gen[544]),

			.SO(gen[637]),
			.S(gen[638]),
			.SE(gen[639]),

			.SELF(gen[543]),
			.cell_state(gen[543])
		); 

/******************* CELL 544 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell544 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[448]),
			.N(gen[449]),
			.NE(gen[450]),

			.O(gen[543]),
			.E(gen[545]),

			.SO(gen[638]),
			.S(gen[639]),
			.SE(gen[640]),

			.SELF(gen[544]),
			.cell_state(gen[544])
		); 

/******************* CELL 545 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell545 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[449]),
			.N(gen[450]),
			.NE(gen[451]),

			.O(gen[544]),
			.E(gen[546]),

			.SO(gen[639]),
			.S(gen[640]),
			.SE(gen[641]),

			.SELF(gen[545]),
			.cell_state(gen[545])
		); 

/******************* CELL 546 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell546 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[450]),
			.N(gen[451]),
			.NE(gen[452]),

			.O(gen[545]),
			.E(gen[547]),

			.SO(gen[640]),
			.S(gen[641]),
			.SE(gen[642]),

			.SELF(gen[546]),
			.cell_state(gen[546])
		); 

/******************* CELL 547 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell547 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[451]),
			.N(gen[452]),
			.NE(gen[453]),

			.O(gen[546]),
			.E(gen[548]),

			.SO(gen[641]),
			.S(gen[642]),
			.SE(gen[643]),

			.SELF(gen[547]),
			.cell_state(gen[547])
		); 

/******************* CELL 548 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell548 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[452]),
			.N(gen[453]),
			.NE(gen[454]),

			.O(gen[547]),
			.E(gen[549]),

			.SO(gen[642]),
			.S(gen[643]),
			.SE(gen[644]),

			.SELF(gen[548]),
			.cell_state(gen[548])
		); 

/******************* CELL 549 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell549 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[453]),
			.N(gen[454]),
			.NE(gen[455]),

			.O(gen[548]),
			.E(gen[550]),

			.SO(gen[643]),
			.S(gen[644]),
			.SE(gen[645]),

			.SELF(gen[549]),
			.cell_state(gen[549])
		); 

/******************* CELL 550 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell550 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[454]),
			.N(gen[455]),
			.NE(gen[456]),

			.O(gen[549]),
			.E(gen[551]),

			.SO(gen[644]),
			.S(gen[645]),
			.SE(gen[646]),

			.SELF(gen[550]),
			.cell_state(gen[550])
		); 

/******************* CELL 551 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell551 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[455]),
			.N(gen[456]),
			.NE(gen[457]),

			.O(gen[550]),
			.E(gen[552]),

			.SO(gen[645]),
			.S(gen[646]),
			.SE(gen[647]),

			.SELF(gen[551]),
			.cell_state(gen[551])
		); 

/******************* CELL 552 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell552 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[456]),
			.N(gen[457]),
			.NE(gen[458]),

			.O(gen[551]),
			.E(gen[553]),

			.SO(gen[646]),
			.S(gen[647]),
			.SE(gen[648]),

			.SELF(gen[552]),
			.cell_state(gen[552])
		); 

/******************* CELL 553 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell553 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[457]),
			.N(gen[458]),
			.NE(gen[459]),

			.O(gen[552]),
			.E(gen[554]),

			.SO(gen[647]),
			.S(gen[648]),
			.SE(gen[649]),

			.SELF(gen[553]),
			.cell_state(gen[553])
		); 

/******************* CELL 554 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell554 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[458]),
			.N(gen[459]),
			.NE(gen[460]),

			.O(gen[553]),
			.E(gen[555]),

			.SO(gen[648]),
			.S(gen[649]),
			.SE(gen[650]),

			.SELF(gen[554]),
			.cell_state(gen[554])
		); 

/******************* CELL 555 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell555 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[459]),
			.N(gen[460]),
			.NE(gen[461]),

			.O(gen[554]),
			.E(gen[556]),

			.SO(gen[649]),
			.S(gen[650]),
			.SE(gen[651]),

			.SELF(gen[555]),
			.cell_state(gen[555])
		); 

/******************* CELL 556 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell556 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[460]),
			.N(gen[461]),
			.NE(gen[462]),

			.O(gen[555]),
			.E(gen[557]),

			.SO(gen[650]),
			.S(gen[651]),
			.SE(gen[652]),

			.SELF(gen[556]),
			.cell_state(gen[556])
		); 

/******************* CELL 557 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell557 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[461]),
			.N(gen[462]),
			.NE(gen[463]),

			.O(gen[556]),
			.E(gen[558]),

			.SO(gen[651]),
			.S(gen[652]),
			.SE(gen[653]),

			.SELF(gen[557]),
			.cell_state(gen[557])
		); 

/******************* CELL 558 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell558 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[462]),
			.N(gen[463]),
			.NE(gen[464]),

			.O(gen[557]),
			.E(gen[559]),

			.SO(gen[652]),
			.S(gen[653]),
			.SE(gen[654]),

			.SELF(gen[558]),
			.cell_state(gen[558])
		); 

/******************* CELL 559 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell559 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[463]),
			.N(gen[464]),
			.NE(gen[465]),

			.O(gen[558]),
			.E(gen[560]),

			.SO(gen[653]),
			.S(gen[654]),
			.SE(gen[655]),

			.SELF(gen[559]),
			.cell_state(gen[559])
		); 

/******************* CELL 560 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell560 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[464]),
			.N(gen[465]),
			.NE(gen[466]),

			.O(gen[559]),
			.E(gen[561]),

			.SO(gen[654]),
			.S(gen[655]),
			.SE(gen[656]),

			.SELF(gen[560]),
			.cell_state(gen[560])
		); 

/******************* CELL 561 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell561 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[465]),
			.N(gen[466]),
			.NE(gen[467]),

			.O(gen[560]),
			.E(gen[562]),

			.SO(gen[655]),
			.S(gen[656]),
			.SE(gen[657]),

			.SELF(gen[561]),
			.cell_state(gen[561])
		); 

/******************* CELL 562 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell562 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[466]),
			.N(gen[467]),
			.NE(gen[468]),

			.O(gen[561]),
			.E(gen[563]),

			.SO(gen[656]),
			.S(gen[657]),
			.SE(gen[658]),

			.SELF(gen[562]),
			.cell_state(gen[562])
		); 

/******************* CELL 563 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell563 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[467]),
			.N(gen[468]),
			.NE(gen[469]),

			.O(gen[562]),
			.E(gen[564]),

			.SO(gen[657]),
			.S(gen[658]),
			.SE(gen[659]),

			.SELF(gen[563]),
			.cell_state(gen[563])
		); 

/******************* CELL 564 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell564 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[468]),
			.N(gen[469]),
			.NE(gen[470]),

			.O(gen[563]),
			.E(gen[565]),

			.SO(gen[658]),
			.S(gen[659]),
			.SE(gen[660]),

			.SELF(gen[564]),
			.cell_state(gen[564])
		); 

/******************* CELL 565 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell565 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[469]),
			.N(gen[470]),
			.NE(gen[471]),

			.O(gen[564]),
			.E(gen[566]),

			.SO(gen[659]),
			.S(gen[660]),
			.SE(gen[661]),

			.SELF(gen[565]),
			.cell_state(gen[565])
		); 

/******************* CELL 566 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell566 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[470]),
			.N(gen[471]),
			.NE(gen[472]),

			.O(gen[565]),
			.E(gen[567]),

			.SO(gen[660]),
			.S(gen[661]),
			.SE(gen[662]),

			.SELF(gen[566]),
			.cell_state(gen[566])
		); 

/******************* CELL 567 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell567 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[471]),
			.N(gen[472]),
			.NE(gen[473]),

			.O(gen[566]),
			.E(gen[568]),

			.SO(gen[661]),
			.S(gen[662]),
			.SE(gen[663]),

			.SELF(gen[567]),
			.cell_state(gen[567])
		); 

/******************* CELL 568 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell568 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[472]),
			.N(gen[473]),
			.NE(gen[474]),

			.O(gen[567]),
			.E(gen[569]),

			.SO(gen[662]),
			.S(gen[663]),
			.SE(gen[664]),

			.SELF(gen[568]),
			.cell_state(gen[568])
		); 

/******************* CELL 569 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell569 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[473]),
			.N(gen[474]),
			.NE(gen[473]),

			.O(gen[568]),
			.E(gen[568]),

			.SO(gen[663]),
			.S(gen[664]),
			.SE(gen[663]),

			.SELF(gen[569]),
			.cell_state(gen[569])
		); 

/******************* CELL 570 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell570 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[476]),
			.N(gen[475]),
			.NE(gen[476]),

			.O(gen[571]),
			.E(gen[571]),

			.SO(gen[666]),
			.S(gen[665]),
			.SE(gen[666]),

			.SELF(gen[570]),
			.cell_state(gen[570])
		); 

/******************* CELL 571 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell571 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[475]),
			.N(gen[476]),
			.NE(gen[477]),

			.O(gen[570]),
			.E(gen[572]),

			.SO(gen[665]),
			.S(gen[666]),
			.SE(gen[667]),

			.SELF(gen[571]),
			.cell_state(gen[571])
		); 

/******************* CELL 572 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell572 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[476]),
			.N(gen[477]),
			.NE(gen[478]),

			.O(gen[571]),
			.E(gen[573]),

			.SO(gen[666]),
			.S(gen[667]),
			.SE(gen[668]),

			.SELF(gen[572]),
			.cell_state(gen[572])
		); 

/******************* CELL 573 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell573 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[477]),
			.N(gen[478]),
			.NE(gen[479]),

			.O(gen[572]),
			.E(gen[574]),

			.SO(gen[667]),
			.S(gen[668]),
			.SE(gen[669]),

			.SELF(gen[573]),
			.cell_state(gen[573])
		); 

/******************* CELL 574 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell574 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[478]),
			.N(gen[479]),
			.NE(gen[480]),

			.O(gen[573]),
			.E(gen[575]),

			.SO(gen[668]),
			.S(gen[669]),
			.SE(gen[670]),

			.SELF(gen[574]),
			.cell_state(gen[574])
		); 

/******************* CELL 575 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell575 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[479]),
			.N(gen[480]),
			.NE(gen[481]),

			.O(gen[574]),
			.E(gen[576]),

			.SO(gen[669]),
			.S(gen[670]),
			.SE(gen[671]),

			.SELF(gen[575]),
			.cell_state(gen[575])
		); 

/******************* CELL 576 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell576 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[480]),
			.N(gen[481]),
			.NE(gen[482]),

			.O(gen[575]),
			.E(gen[577]),

			.SO(gen[670]),
			.S(gen[671]),
			.SE(gen[672]),

			.SELF(gen[576]),
			.cell_state(gen[576])
		); 

/******************* CELL 577 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell577 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[481]),
			.N(gen[482]),
			.NE(gen[483]),

			.O(gen[576]),
			.E(gen[578]),

			.SO(gen[671]),
			.S(gen[672]),
			.SE(gen[673]),

			.SELF(gen[577]),
			.cell_state(gen[577])
		); 

/******************* CELL 578 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell578 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[482]),
			.N(gen[483]),
			.NE(gen[484]),

			.O(gen[577]),
			.E(gen[579]),

			.SO(gen[672]),
			.S(gen[673]),
			.SE(gen[674]),

			.SELF(gen[578]),
			.cell_state(gen[578])
		); 

/******************* CELL 579 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell579 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[483]),
			.N(gen[484]),
			.NE(gen[485]),

			.O(gen[578]),
			.E(gen[580]),

			.SO(gen[673]),
			.S(gen[674]),
			.SE(gen[675]),

			.SELF(gen[579]),
			.cell_state(gen[579])
		); 

/******************* CELL 580 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell580 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[484]),
			.N(gen[485]),
			.NE(gen[486]),

			.O(gen[579]),
			.E(gen[581]),

			.SO(gen[674]),
			.S(gen[675]),
			.SE(gen[676]),

			.SELF(gen[580]),
			.cell_state(gen[580])
		); 

/******************* CELL 581 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell581 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[485]),
			.N(gen[486]),
			.NE(gen[487]),

			.O(gen[580]),
			.E(gen[582]),

			.SO(gen[675]),
			.S(gen[676]),
			.SE(gen[677]),

			.SELF(gen[581]),
			.cell_state(gen[581])
		); 

/******************* CELL 582 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell582 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[486]),
			.N(gen[487]),
			.NE(gen[488]),

			.O(gen[581]),
			.E(gen[583]),

			.SO(gen[676]),
			.S(gen[677]),
			.SE(gen[678]),

			.SELF(gen[582]),
			.cell_state(gen[582])
		); 

/******************* CELL 583 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell583 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[487]),
			.N(gen[488]),
			.NE(gen[489]),

			.O(gen[582]),
			.E(gen[584]),

			.SO(gen[677]),
			.S(gen[678]),
			.SE(gen[679]),

			.SELF(gen[583]),
			.cell_state(gen[583])
		); 

/******************* CELL 584 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell584 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[488]),
			.N(gen[489]),
			.NE(gen[490]),

			.O(gen[583]),
			.E(gen[585]),

			.SO(gen[678]),
			.S(gen[679]),
			.SE(gen[680]),

			.SELF(gen[584]),
			.cell_state(gen[584])
		); 

/******************* CELL 585 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell585 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[489]),
			.N(gen[490]),
			.NE(gen[491]),

			.O(gen[584]),
			.E(gen[586]),

			.SO(gen[679]),
			.S(gen[680]),
			.SE(gen[681]),

			.SELF(gen[585]),
			.cell_state(gen[585])
		); 

/******************* CELL 586 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell586 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[490]),
			.N(gen[491]),
			.NE(gen[492]),

			.O(gen[585]),
			.E(gen[587]),

			.SO(gen[680]),
			.S(gen[681]),
			.SE(gen[682]),

			.SELF(gen[586]),
			.cell_state(gen[586])
		); 

/******************* CELL 587 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell587 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[491]),
			.N(gen[492]),
			.NE(gen[493]),

			.O(gen[586]),
			.E(gen[588]),

			.SO(gen[681]),
			.S(gen[682]),
			.SE(gen[683]),

			.SELF(gen[587]),
			.cell_state(gen[587])
		); 

/******************* CELL 588 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell588 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[492]),
			.N(gen[493]),
			.NE(gen[494]),

			.O(gen[587]),
			.E(gen[589]),

			.SO(gen[682]),
			.S(gen[683]),
			.SE(gen[684]),

			.SELF(gen[588]),
			.cell_state(gen[588])
		); 

/******************* CELL 589 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell589 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[493]),
			.N(gen[494]),
			.NE(gen[495]),

			.O(gen[588]),
			.E(gen[590]),

			.SO(gen[683]),
			.S(gen[684]),
			.SE(gen[685]),

			.SELF(gen[589]),
			.cell_state(gen[589])
		); 

/******************* CELL 590 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell590 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[494]),
			.N(gen[495]),
			.NE(gen[496]),

			.O(gen[589]),
			.E(gen[591]),

			.SO(gen[684]),
			.S(gen[685]),
			.SE(gen[686]),

			.SELF(gen[590]),
			.cell_state(gen[590])
		); 

/******************* CELL 591 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell591 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[495]),
			.N(gen[496]),
			.NE(gen[497]),

			.O(gen[590]),
			.E(gen[592]),

			.SO(gen[685]),
			.S(gen[686]),
			.SE(gen[687]),

			.SELF(gen[591]),
			.cell_state(gen[591])
		); 

/******************* CELL 592 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell592 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[496]),
			.N(gen[497]),
			.NE(gen[498]),

			.O(gen[591]),
			.E(gen[593]),

			.SO(gen[686]),
			.S(gen[687]),
			.SE(gen[688]),

			.SELF(gen[592]),
			.cell_state(gen[592])
		); 

/******************* CELL 593 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell593 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[497]),
			.N(gen[498]),
			.NE(gen[499]),

			.O(gen[592]),
			.E(gen[594]),

			.SO(gen[687]),
			.S(gen[688]),
			.SE(gen[689]),

			.SELF(gen[593]),
			.cell_state(gen[593])
		); 

/******************* CELL 594 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell594 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[498]),
			.N(gen[499]),
			.NE(gen[500]),

			.O(gen[593]),
			.E(gen[595]),

			.SO(gen[688]),
			.S(gen[689]),
			.SE(gen[690]),

			.SELF(gen[594]),
			.cell_state(gen[594])
		); 

/******************* CELL 595 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell595 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[499]),
			.N(gen[500]),
			.NE(gen[501]),

			.O(gen[594]),
			.E(gen[596]),

			.SO(gen[689]),
			.S(gen[690]),
			.SE(gen[691]),

			.SELF(gen[595]),
			.cell_state(gen[595])
		); 

/******************* CELL 596 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell596 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[500]),
			.N(gen[501]),
			.NE(gen[502]),

			.O(gen[595]),
			.E(gen[597]),

			.SO(gen[690]),
			.S(gen[691]),
			.SE(gen[692]),

			.SELF(gen[596]),
			.cell_state(gen[596])
		); 

/******************* CELL 597 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell597 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[501]),
			.N(gen[502]),
			.NE(gen[503]),

			.O(gen[596]),
			.E(gen[598]),

			.SO(gen[691]),
			.S(gen[692]),
			.SE(gen[693]),

			.SELF(gen[597]),
			.cell_state(gen[597])
		); 

/******************* CELL 598 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell598 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[502]),
			.N(gen[503]),
			.NE(gen[504]),

			.O(gen[597]),
			.E(gen[599]),

			.SO(gen[692]),
			.S(gen[693]),
			.SE(gen[694]),

			.SELF(gen[598]),
			.cell_state(gen[598])
		); 

/******************* CELL 599 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell599 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[503]),
			.N(gen[504]),
			.NE(gen[505]),

			.O(gen[598]),
			.E(gen[600]),

			.SO(gen[693]),
			.S(gen[694]),
			.SE(gen[695]),

			.SELF(gen[599]),
			.cell_state(gen[599])
		); 

/******************* CELL 600 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell600 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[504]),
			.N(gen[505]),
			.NE(gen[506]),

			.O(gen[599]),
			.E(gen[601]),

			.SO(gen[694]),
			.S(gen[695]),
			.SE(gen[696]),

			.SELF(gen[600]),
			.cell_state(gen[600])
		); 

/******************* CELL 601 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell601 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[505]),
			.N(gen[506]),
			.NE(gen[507]),

			.O(gen[600]),
			.E(gen[602]),

			.SO(gen[695]),
			.S(gen[696]),
			.SE(gen[697]),

			.SELF(gen[601]),
			.cell_state(gen[601])
		); 

/******************* CELL 602 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell602 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[506]),
			.N(gen[507]),
			.NE(gen[508]),

			.O(gen[601]),
			.E(gen[603]),

			.SO(gen[696]),
			.S(gen[697]),
			.SE(gen[698]),

			.SELF(gen[602]),
			.cell_state(gen[602])
		); 

/******************* CELL 603 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell603 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[507]),
			.N(gen[508]),
			.NE(gen[509]),

			.O(gen[602]),
			.E(gen[604]),

			.SO(gen[697]),
			.S(gen[698]),
			.SE(gen[699]),

			.SELF(gen[603]),
			.cell_state(gen[603])
		); 

/******************* CELL 604 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell604 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[508]),
			.N(gen[509]),
			.NE(gen[510]),

			.O(gen[603]),
			.E(gen[605]),

			.SO(gen[698]),
			.S(gen[699]),
			.SE(gen[700]),

			.SELF(gen[604]),
			.cell_state(gen[604])
		); 

/******************* CELL 605 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell605 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[509]),
			.N(gen[510]),
			.NE(gen[511]),

			.O(gen[604]),
			.E(gen[606]),

			.SO(gen[699]),
			.S(gen[700]),
			.SE(gen[701]),

			.SELF(gen[605]),
			.cell_state(gen[605])
		); 

/******************* CELL 606 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell606 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[510]),
			.N(gen[511]),
			.NE(gen[512]),

			.O(gen[605]),
			.E(gen[607]),

			.SO(gen[700]),
			.S(gen[701]),
			.SE(gen[702]),

			.SELF(gen[606]),
			.cell_state(gen[606])
		); 

/******************* CELL 607 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell607 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[511]),
			.N(gen[512]),
			.NE(gen[513]),

			.O(gen[606]),
			.E(gen[608]),

			.SO(gen[701]),
			.S(gen[702]),
			.SE(gen[703]),

			.SELF(gen[607]),
			.cell_state(gen[607])
		); 

/******************* CELL 608 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell608 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[512]),
			.N(gen[513]),
			.NE(gen[514]),

			.O(gen[607]),
			.E(gen[609]),

			.SO(gen[702]),
			.S(gen[703]),
			.SE(gen[704]),

			.SELF(gen[608]),
			.cell_state(gen[608])
		); 

/******************* CELL 609 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell609 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[513]),
			.N(gen[514]),
			.NE(gen[515]),

			.O(gen[608]),
			.E(gen[610]),

			.SO(gen[703]),
			.S(gen[704]),
			.SE(gen[705]),

			.SELF(gen[609]),
			.cell_state(gen[609])
		); 

/******************* CELL 610 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell610 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[514]),
			.N(gen[515]),
			.NE(gen[516]),

			.O(gen[609]),
			.E(gen[611]),

			.SO(gen[704]),
			.S(gen[705]),
			.SE(gen[706]),

			.SELF(gen[610]),
			.cell_state(gen[610])
		); 

/******************* CELL 611 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell611 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[515]),
			.N(gen[516]),
			.NE(gen[517]),

			.O(gen[610]),
			.E(gen[612]),

			.SO(gen[705]),
			.S(gen[706]),
			.SE(gen[707]),

			.SELF(gen[611]),
			.cell_state(gen[611])
		); 

/******************* CELL 612 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell612 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[516]),
			.N(gen[517]),
			.NE(gen[518]),

			.O(gen[611]),
			.E(gen[613]),

			.SO(gen[706]),
			.S(gen[707]),
			.SE(gen[708]),

			.SELF(gen[612]),
			.cell_state(gen[612])
		); 

/******************* CELL 613 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell613 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[517]),
			.N(gen[518]),
			.NE(gen[519]),

			.O(gen[612]),
			.E(gen[614]),

			.SO(gen[707]),
			.S(gen[708]),
			.SE(gen[709]),

			.SELF(gen[613]),
			.cell_state(gen[613])
		); 

/******************* CELL 614 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell614 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[518]),
			.N(gen[519]),
			.NE(gen[520]),

			.O(gen[613]),
			.E(gen[615]),

			.SO(gen[708]),
			.S(gen[709]),
			.SE(gen[710]),

			.SELF(gen[614]),
			.cell_state(gen[614])
		); 

/******************* CELL 615 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell615 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[519]),
			.N(gen[520]),
			.NE(gen[521]),

			.O(gen[614]),
			.E(gen[616]),

			.SO(gen[709]),
			.S(gen[710]),
			.SE(gen[711]),

			.SELF(gen[615]),
			.cell_state(gen[615])
		); 

/******************* CELL 616 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell616 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[520]),
			.N(gen[521]),
			.NE(gen[522]),

			.O(gen[615]),
			.E(gen[617]),

			.SO(gen[710]),
			.S(gen[711]),
			.SE(gen[712]),

			.SELF(gen[616]),
			.cell_state(gen[616])
		); 

/******************* CELL 617 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell617 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[521]),
			.N(gen[522]),
			.NE(gen[523]),

			.O(gen[616]),
			.E(gen[618]),

			.SO(gen[711]),
			.S(gen[712]),
			.SE(gen[713]),

			.SELF(gen[617]),
			.cell_state(gen[617])
		); 

/******************* CELL 618 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell618 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[522]),
			.N(gen[523]),
			.NE(gen[524]),

			.O(gen[617]),
			.E(gen[619]),

			.SO(gen[712]),
			.S(gen[713]),
			.SE(gen[714]),

			.SELF(gen[618]),
			.cell_state(gen[618])
		); 

/******************* CELL 619 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell619 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[523]),
			.N(gen[524]),
			.NE(gen[525]),

			.O(gen[618]),
			.E(gen[620]),

			.SO(gen[713]),
			.S(gen[714]),
			.SE(gen[715]),

			.SELF(gen[619]),
			.cell_state(gen[619])
		); 

/******************* CELL 620 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell620 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[524]),
			.N(gen[525]),
			.NE(gen[526]),

			.O(gen[619]),
			.E(gen[621]),

			.SO(gen[714]),
			.S(gen[715]),
			.SE(gen[716]),

			.SELF(gen[620]),
			.cell_state(gen[620])
		); 

/******************* CELL 621 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell621 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[525]),
			.N(gen[526]),
			.NE(gen[527]),

			.O(gen[620]),
			.E(gen[622]),

			.SO(gen[715]),
			.S(gen[716]),
			.SE(gen[717]),

			.SELF(gen[621]),
			.cell_state(gen[621])
		); 

/******************* CELL 622 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell622 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[526]),
			.N(gen[527]),
			.NE(gen[528]),

			.O(gen[621]),
			.E(gen[623]),

			.SO(gen[716]),
			.S(gen[717]),
			.SE(gen[718]),

			.SELF(gen[622]),
			.cell_state(gen[622])
		); 

/******************* CELL 623 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell623 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[527]),
			.N(gen[528]),
			.NE(gen[529]),

			.O(gen[622]),
			.E(gen[624]),

			.SO(gen[717]),
			.S(gen[718]),
			.SE(gen[719]),

			.SELF(gen[623]),
			.cell_state(gen[623])
		); 

/******************* CELL 624 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell624 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[528]),
			.N(gen[529]),
			.NE(gen[530]),

			.O(gen[623]),
			.E(gen[625]),

			.SO(gen[718]),
			.S(gen[719]),
			.SE(gen[720]),

			.SELF(gen[624]),
			.cell_state(gen[624])
		); 

/******************* CELL 625 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell625 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[529]),
			.N(gen[530]),
			.NE(gen[531]),

			.O(gen[624]),
			.E(gen[626]),

			.SO(gen[719]),
			.S(gen[720]),
			.SE(gen[721]),

			.SELF(gen[625]),
			.cell_state(gen[625])
		); 

/******************* CELL 626 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell626 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[530]),
			.N(gen[531]),
			.NE(gen[532]),

			.O(gen[625]),
			.E(gen[627]),

			.SO(gen[720]),
			.S(gen[721]),
			.SE(gen[722]),

			.SELF(gen[626]),
			.cell_state(gen[626])
		); 

/******************* CELL 627 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell627 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[531]),
			.N(gen[532]),
			.NE(gen[533]),

			.O(gen[626]),
			.E(gen[628]),

			.SO(gen[721]),
			.S(gen[722]),
			.SE(gen[723]),

			.SELF(gen[627]),
			.cell_state(gen[627])
		); 

/******************* CELL 628 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell628 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[532]),
			.N(gen[533]),
			.NE(gen[534]),

			.O(gen[627]),
			.E(gen[629]),

			.SO(gen[722]),
			.S(gen[723]),
			.SE(gen[724]),

			.SELF(gen[628]),
			.cell_state(gen[628])
		); 

/******************* CELL 629 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell629 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[533]),
			.N(gen[534]),
			.NE(gen[535]),

			.O(gen[628]),
			.E(gen[630]),

			.SO(gen[723]),
			.S(gen[724]),
			.SE(gen[725]),

			.SELF(gen[629]),
			.cell_state(gen[629])
		); 

/******************* CELL 630 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell630 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[534]),
			.N(gen[535]),
			.NE(gen[536]),

			.O(gen[629]),
			.E(gen[631]),

			.SO(gen[724]),
			.S(gen[725]),
			.SE(gen[726]),

			.SELF(gen[630]),
			.cell_state(gen[630])
		); 

/******************* CELL 631 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell631 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[535]),
			.N(gen[536]),
			.NE(gen[537]),

			.O(gen[630]),
			.E(gen[632]),

			.SO(gen[725]),
			.S(gen[726]),
			.SE(gen[727]),

			.SELF(gen[631]),
			.cell_state(gen[631])
		); 

/******************* CELL 632 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell632 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[536]),
			.N(gen[537]),
			.NE(gen[538]),

			.O(gen[631]),
			.E(gen[633]),

			.SO(gen[726]),
			.S(gen[727]),
			.SE(gen[728]),

			.SELF(gen[632]),
			.cell_state(gen[632])
		); 

/******************* CELL 633 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell633 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[537]),
			.N(gen[538]),
			.NE(gen[539]),

			.O(gen[632]),
			.E(gen[634]),

			.SO(gen[727]),
			.S(gen[728]),
			.SE(gen[729]),

			.SELF(gen[633]),
			.cell_state(gen[633])
		); 

/******************* CELL 634 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell634 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[538]),
			.N(gen[539]),
			.NE(gen[540]),

			.O(gen[633]),
			.E(gen[635]),

			.SO(gen[728]),
			.S(gen[729]),
			.SE(gen[730]),

			.SELF(gen[634]),
			.cell_state(gen[634])
		); 

/******************* CELL 635 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell635 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[539]),
			.N(gen[540]),
			.NE(gen[541]),

			.O(gen[634]),
			.E(gen[636]),

			.SO(gen[729]),
			.S(gen[730]),
			.SE(gen[731]),

			.SELF(gen[635]),
			.cell_state(gen[635])
		); 

/******************* CELL 636 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell636 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[540]),
			.N(gen[541]),
			.NE(gen[542]),

			.O(gen[635]),
			.E(gen[637]),

			.SO(gen[730]),
			.S(gen[731]),
			.SE(gen[732]),

			.SELF(gen[636]),
			.cell_state(gen[636])
		); 

/******************* CELL 637 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell637 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[541]),
			.N(gen[542]),
			.NE(gen[543]),

			.O(gen[636]),
			.E(gen[638]),

			.SO(gen[731]),
			.S(gen[732]),
			.SE(gen[733]),

			.SELF(gen[637]),
			.cell_state(gen[637])
		); 

/******************* CELL 638 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell638 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[542]),
			.N(gen[543]),
			.NE(gen[544]),

			.O(gen[637]),
			.E(gen[639]),

			.SO(gen[732]),
			.S(gen[733]),
			.SE(gen[734]),

			.SELF(gen[638]),
			.cell_state(gen[638])
		); 

/******************* CELL 639 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell639 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[543]),
			.N(gen[544]),
			.NE(gen[545]),

			.O(gen[638]),
			.E(gen[640]),

			.SO(gen[733]),
			.S(gen[734]),
			.SE(gen[735]),

			.SELF(gen[639]),
			.cell_state(gen[639])
		); 

/******************* CELL 640 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell640 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[544]),
			.N(gen[545]),
			.NE(gen[546]),

			.O(gen[639]),
			.E(gen[641]),

			.SO(gen[734]),
			.S(gen[735]),
			.SE(gen[736]),

			.SELF(gen[640]),
			.cell_state(gen[640])
		); 

/******************* CELL 641 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell641 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[545]),
			.N(gen[546]),
			.NE(gen[547]),

			.O(gen[640]),
			.E(gen[642]),

			.SO(gen[735]),
			.S(gen[736]),
			.SE(gen[737]),

			.SELF(gen[641]),
			.cell_state(gen[641])
		); 

/******************* CELL 642 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell642 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[546]),
			.N(gen[547]),
			.NE(gen[548]),

			.O(gen[641]),
			.E(gen[643]),

			.SO(gen[736]),
			.S(gen[737]),
			.SE(gen[738]),

			.SELF(gen[642]),
			.cell_state(gen[642])
		); 

/******************* CELL 643 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell643 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[547]),
			.N(gen[548]),
			.NE(gen[549]),

			.O(gen[642]),
			.E(gen[644]),

			.SO(gen[737]),
			.S(gen[738]),
			.SE(gen[739]),

			.SELF(gen[643]),
			.cell_state(gen[643])
		); 

/******************* CELL 644 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell644 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[548]),
			.N(gen[549]),
			.NE(gen[550]),

			.O(gen[643]),
			.E(gen[645]),

			.SO(gen[738]),
			.S(gen[739]),
			.SE(gen[740]),

			.SELF(gen[644]),
			.cell_state(gen[644])
		); 

/******************* CELL 645 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell645 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[549]),
			.N(gen[550]),
			.NE(gen[551]),

			.O(gen[644]),
			.E(gen[646]),

			.SO(gen[739]),
			.S(gen[740]),
			.SE(gen[741]),

			.SELF(gen[645]),
			.cell_state(gen[645])
		); 

/******************* CELL 646 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell646 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[550]),
			.N(gen[551]),
			.NE(gen[552]),

			.O(gen[645]),
			.E(gen[647]),

			.SO(gen[740]),
			.S(gen[741]),
			.SE(gen[742]),

			.SELF(gen[646]),
			.cell_state(gen[646])
		); 

/******************* CELL 647 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell647 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[551]),
			.N(gen[552]),
			.NE(gen[553]),

			.O(gen[646]),
			.E(gen[648]),

			.SO(gen[741]),
			.S(gen[742]),
			.SE(gen[743]),

			.SELF(gen[647]),
			.cell_state(gen[647])
		); 

/******************* CELL 648 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell648 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[552]),
			.N(gen[553]),
			.NE(gen[554]),

			.O(gen[647]),
			.E(gen[649]),

			.SO(gen[742]),
			.S(gen[743]),
			.SE(gen[744]),

			.SELF(gen[648]),
			.cell_state(gen[648])
		); 

/******************* CELL 649 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell649 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[553]),
			.N(gen[554]),
			.NE(gen[555]),

			.O(gen[648]),
			.E(gen[650]),

			.SO(gen[743]),
			.S(gen[744]),
			.SE(gen[745]),

			.SELF(gen[649]),
			.cell_state(gen[649])
		); 

/******************* CELL 650 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell650 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[554]),
			.N(gen[555]),
			.NE(gen[556]),

			.O(gen[649]),
			.E(gen[651]),

			.SO(gen[744]),
			.S(gen[745]),
			.SE(gen[746]),

			.SELF(gen[650]),
			.cell_state(gen[650])
		); 

/******************* CELL 651 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell651 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[555]),
			.N(gen[556]),
			.NE(gen[557]),

			.O(gen[650]),
			.E(gen[652]),

			.SO(gen[745]),
			.S(gen[746]),
			.SE(gen[747]),

			.SELF(gen[651]),
			.cell_state(gen[651])
		); 

/******************* CELL 652 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell652 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[556]),
			.N(gen[557]),
			.NE(gen[558]),

			.O(gen[651]),
			.E(gen[653]),

			.SO(gen[746]),
			.S(gen[747]),
			.SE(gen[748]),

			.SELF(gen[652]),
			.cell_state(gen[652])
		); 

/******************* CELL 653 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell653 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[557]),
			.N(gen[558]),
			.NE(gen[559]),

			.O(gen[652]),
			.E(gen[654]),

			.SO(gen[747]),
			.S(gen[748]),
			.SE(gen[749]),

			.SELF(gen[653]),
			.cell_state(gen[653])
		); 

/******************* CELL 654 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell654 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[558]),
			.N(gen[559]),
			.NE(gen[560]),

			.O(gen[653]),
			.E(gen[655]),

			.SO(gen[748]),
			.S(gen[749]),
			.SE(gen[750]),

			.SELF(gen[654]),
			.cell_state(gen[654])
		); 

/******************* CELL 655 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell655 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[559]),
			.N(gen[560]),
			.NE(gen[561]),

			.O(gen[654]),
			.E(gen[656]),

			.SO(gen[749]),
			.S(gen[750]),
			.SE(gen[751]),

			.SELF(gen[655]),
			.cell_state(gen[655])
		); 

/******************* CELL 656 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell656 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[560]),
			.N(gen[561]),
			.NE(gen[562]),

			.O(gen[655]),
			.E(gen[657]),

			.SO(gen[750]),
			.S(gen[751]),
			.SE(gen[752]),

			.SELF(gen[656]),
			.cell_state(gen[656])
		); 

/******************* CELL 657 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell657 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[561]),
			.N(gen[562]),
			.NE(gen[563]),

			.O(gen[656]),
			.E(gen[658]),

			.SO(gen[751]),
			.S(gen[752]),
			.SE(gen[753]),

			.SELF(gen[657]),
			.cell_state(gen[657])
		); 

/******************* CELL 658 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell658 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[562]),
			.N(gen[563]),
			.NE(gen[564]),

			.O(gen[657]),
			.E(gen[659]),

			.SO(gen[752]),
			.S(gen[753]),
			.SE(gen[754]),

			.SELF(gen[658]),
			.cell_state(gen[658])
		); 

/******************* CELL 659 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell659 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[563]),
			.N(gen[564]),
			.NE(gen[565]),

			.O(gen[658]),
			.E(gen[660]),

			.SO(gen[753]),
			.S(gen[754]),
			.SE(gen[755]),

			.SELF(gen[659]),
			.cell_state(gen[659])
		); 

/******************* CELL 660 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell660 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[564]),
			.N(gen[565]),
			.NE(gen[566]),

			.O(gen[659]),
			.E(gen[661]),

			.SO(gen[754]),
			.S(gen[755]),
			.SE(gen[756]),

			.SELF(gen[660]),
			.cell_state(gen[660])
		); 

/******************* CELL 661 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell661 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[565]),
			.N(gen[566]),
			.NE(gen[567]),

			.O(gen[660]),
			.E(gen[662]),

			.SO(gen[755]),
			.S(gen[756]),
			.SE(gen[757]),

			.SELF(gen[661]),
			.cell_state(gen[661])
		); 

/******************* CELL 662 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell662 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[566]),
			.N(gen[567]),
			.NE(gen[568]),

			.O(gen[661]),
			.E(gen[663]),

			.SO(gen[756]),
			.S(gen[757]),
			.SE(gen[758]),

			.SELF(gen[662]),
			.cell_state(gen[662])
		); 

/******************* CELL 663 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell663 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[567]),
			.N(gen[568]),
			.NE(gen[569]),

			.O(gen[662]),
			.E(gen[664]),

			.SO(gen[757]),
			.S(gen[758]),
			.SE(gen[759]),

			.SELF(gen[663]),
			.cell_state(gen[663])
		); 

/******************* CELL 664 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell664 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[568]),
			.N(gen[569]),
			.NE(gen[568]),

			.O(gen[663]),
			.E(gen[663]),

			.SO(gen[758]),
			.S(gen[759]),
			.SE(gen[758]),

			.SELF(gen[664]),
			.cell_state(gen[664])
		); 

/******************* CELL 665 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell665 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[571]),
			.N(gen[570]),
			.NE(gen[571]),

			.O(gen[666]),
			.E(gen[666]),

			.SO(gen[761]),
			.S(gen[760]),
			.SE(gen[761]),

			.SELF(gen[665]),
			.cell_state(gen[665])
		); 

/******************* CELL 666 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell666 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[570]),
			.N(gen[571]),
			.NE(gen[572]),

			.O(gen[665]),
			.E(gen[667]),

			.SO(gen[760]),
			.S(gen[761]),
			.SE(gen[762]),

			.SELF(gen[666]),
			.cell_state(gen[666])
		); 

/******************* CELL 667 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell667 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[571]),
			.N(gen[572]),
			.NE(gen[573]),

			.O(gen[666]),
			.E(gen[668]),

			.SO(gen[761]),
			.S(gen[762]),
			.SE(gen[763]),

			.SELF(gen[667]),
			.cell_state(gen[667])
		); 

/******************* CELL 668 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell668 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[572]),
			.N(gen[573]),
			.NE(gen[574]),

			.O(gen[667]),
			.E(gen[669]),

			.SO(gen[762]),
			.S(gen[763]),
			.SE(gen[764]),

			.SELF(gen[668]),
			.cell_state(gen[668])
		); 

/******************* CELL 669 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell669 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[573]),
			.N(gen[574]),
			.NE(gen[575]),

			.O(gen[668]),
			.E(gen[670]),

			.SO(gen[763]),
			.S(gen[764]),
			.SE(gen[765]),

			.SELF(gen[669]),
			.cell_state(gen[669])
		); 

/******************* CELL 670 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell670 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[574]),
			.N(gen[575]),
			.NE(gen[576]),

			.O(gen[669]),
			.E(gen[671]),

			.SO(gen[764]),
			.S(gen[765]),
			.SE(gen[766]),

			.SELF(gen[670]),
			.cell_state(gen[670])
		); 

/******************* CELL 671 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell671 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[575]),
			.N(gen[576]),
			.NE(gen[577]),

			.O(gen[670]),
			.E(gen[672]),

			.SO(gen[765]),
			.S(gen[766]),
			.SE(gen[767]),

			.SELF(gen[671]),
			.cell_state(gen[671])
		); 

/******************* CELL 672 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell672 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[576]),
			.N(gen[577]),
			.NE(gen[578]),

			.O(gen[671]),
			.E(gen[673]),

			.SO(gen[766]),
			.S(gen[767]),
			.SE(gen[768]),

			.SELF(gen[672]),
			.cell_state(gen[672])
		); 

/******************* CELL 673 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell673 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[577]),
			.N(gen[578]),
			.NE(gen[579]),

			.O(gen[672]),
			.E(gen[674]),

			.SO(gen[767]),
			.S(gen[768]),
			.SE(gen[769]),

			.SELF(gen[673]),
			.cell_state(gen[673])
		); 

/******************* CELL 674 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell674 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[578]),
			.N(gen[579]),
			.NE(gen[580]),

			.O(gen[673]),
			.E(gen[675]),

			.SO(gen[768]),
			.S(gen[769]),
			.SE(gen[770]),

			.SELF(gen[674]),
			.cell_state(gen[674])
		); 

/******************* CELL 675 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell675 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[579]),
			.N(gen[580]),
			.NE(gen[581]),

			.O(gen[674]),
			.E(gen[676]),

			.SO(gen[769]),
			.S(gen[770]),
			.SE(gen[771]),

			.SELF(gen[675]),
			.cell_state(gen[675])
		); 

/******************* CELL 676 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell676 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[580]),
			.N(gen[581]),
			.NE(gen[582]),

			.O(gen[675]),
			.E(gen[677]),

			.SO(gen[770]),
			.S(gen[771]),
			.SE(gen[772]),

			.SELF(gen[676]),
			.cell_state(gen[676])
		); 

/******************* CELL 677 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell677 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[581]),
			.N(gen[582]),
			.NE(gen[583]),

			.O(gen[676]),
			.E(gen[678]),

			.SO(gen[771]),
			.S(gen[772]),
			.SE(gen[773]),

			.SELF(gen[677]),
			.cell_state(gen[677])
		); 

/******************* CELL 678 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell678 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[582]),
			.N(gen[583]),
			.NE(gen[584]),

			.O(gen[677]),
			.E(gen[679]),

			.SO(gen[772]),
			.S(gen[773]),
			.SE(gen[774]),

			.SELF(gen[678]),
			.cell_state(gen[678])
		); 

/******************* CELL 679 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell679 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[583]),
			.N(gen[584]),
			.NE(gen[585]),

			.O(gen[678]),
			.E(gen[680]),

			.SO(gen[773]),
			.S(gen[774]),
			.SE(gen[775]),

			.SELF(gen[679]),
			.cell_state(gen[679])
		); 

/******************* CELL 680 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell680 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[584]),
			.N(gen[585]),
			.NE(gen[586]),

			.O(gen[679]),
			.E(gen[681]),

			.SO(gen[774]),
			.S(gen[775]),
			.SE(gen[776]),

			.SELF(gen[680]),
			.cell_state(gen[680])
		); 

/******************* CELL 681 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell681 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[585]),
			.N(gen[586]),
			.NE(gen[587]),

			.O(gen[680]),
			.E(gen[682]),

			.SO(gen[775]),
			.S(gen[776]),
			.SE(gen[777]),

			.SELF(gen[681]),
			.cell_state(gen[681])
		); 

/******************* CELL 682 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell682 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[586]),
			.N(gen[587]),
			.NE(gen[588]),

			.O(gen[681]),
			.E(gen[683]),

			.SO(gen[776]),
			.S(gen[777]),
			.SE(gen[778]),

			.SELF(gen[682]),
			.cell_state(gen[682])
		); 

/******************* CELL 683 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell683 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[587]),
			.N(gen[588]),
			.NE(gen[589]),

			.O(gen[682]),
			.E(gen[684]),

			.SO(gen[777]),
			.S(gen[778]),
			.SE(gen[779]),

			.SELF(gen[683]),
			.cell_state(gen[683])
		); 

/******************* CELL 684 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell684 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[588]),
			.N(gen[589]),
			.NE(gen[590]),

			.O(gen[683]),
			.E(gen[685]),

			.SO(gen[778]),
			.S(gen[779]),
			.SE(gen[780]),

			.SELF(gen[684]),
			.cell_state(gen[684])
		); 

/******************* CELL 685 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell685 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[589]),
			.N(gen[590]),
			.NE(gen[591]),

			.O(gen[684]),
			.E(gen[686]),

			.SO(gen[779]),
			.S(gen[780]),
			.SE(gen[781]),

			.SELF(gen[685]),
			.cell_state(gen[685])
		); 

/******************* CELL 686 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell686 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[590]),
			.N(gen[591]),
			.NE(gen[592]),

			.O(gen[685]),
			.E(gen[687]),

			.SO(gen[780]),
			.S(gen[781]),
			.SE(gen[782]),

			.SELF(gen[686]),
			.cell_state(gen[686])
		); 

/******************* CELL 687 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell687 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[591]),
			.N(gen[592]),
			.NE(gen[593]),

			.O(gen[686]),
			.E(gen[688]),

			.SO(gen[781]),
			.S(gen[782]),
			.SE(gen[783]),

			.SELF(gen[687]),
			.cell_state(gen[687])
		); 

/******************* CELL 688 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell688 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[592]),
			.N(gen[593]),
			.NE(gen[594]),

			.O(gen[687]),
			.E(gen[689]),

			.SO(gen[782]),
			.S(gen[783]),
			.SE(gen[784]),

			.SELF(gen[688]),
			.cell_state(gen[688])
		); 

/******************* CELL 689 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell689 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[593]),
			.N(gen[594]),
			.NE(gen[595]),

			.O(gen[688]),
			.E(gen[690]),

			.SO(gen[783]),
			.S(gen[784]),
			.SE(gen[785]),

			.SELF(gen[689]),
			.cell_state(gen[689])
		); 

/******************* CELL 690 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell690 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[594]),
			.N(gen[595]),
			.NE(gen[596]),

			.O(gen[689]),
			.E(gen[691]),

			.SO(gen[784]),
			.S(gen[785]),
			.SE(gen[786]),

			.SELF(gen[690]),
			.cell_state(gen[690])
		); 

/******************* CELL 691 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell691 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[595]),
			.N(gen[596]),
			.NE(gen[597]),

			.O(gen[690]),
			.E(gen[692]),

			.SO(gen[785]),
			.S(gen[786]),
			.SE(gen[787]),

			.SELF(gen[691]),
			.cell_state(gen[691])
		); 

/******************* CELL 692 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell692 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[596]),
			.N(gen[597]),
			.NE(gen[598]),

			.O(gen[691]),
			.E(gen[693]),

			.SO(gen[786]),
			.S(gen[787]),
			.SE(gen[788]),

			.SELF(gen[692]),
			.cell_state(gen[692])
		); 

/******************* CELL 693 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell693 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[597]),
			.N(gen[598]),
			.NE(gen[599]),

			.O(gen[692]),
			.E(gen[694]),

			.SO(gen[787]),
			.S(gen[788]),
			.SE(gen[789]),

			.SELF(gen[693]),
			.cell_state(gen[693])
		); 

/******************* CELL 694 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell694 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[598]),
			.N(gen[599]),
			.NE(gen[600]),

			.O(gen[693]),
			.E(gen[695]),

			.SO(gen[788]),
			.S(gen[789]),
			.SE(gen[790]),

			.SELF(gen[694]),
			.cell_state(gen[694])
		); 

/******************* CELL 695 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell695 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[599]),
			.N(gen[600]),
			.NE(gen[601]),

			.O(gen[694]),
			.E(gen[696]),

			.SO(gen[789]),
			.S(gen[790]),
			.SE(gen[791]),

			.SELF(gen[695]),
			.cell_state(gen[695])
		); 

/******************* CELL 696 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell696 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[600]),
			.N(gen[601]),
			.NE(gen[602]),

			.O(gen[695]),
			.E(gen[697]),

			.SO(gen[790]),
			.S(gen[791]),
			.SE(gen[792]),

			.SELF(gen[696]),
			.cell_state(gen[696])
		); 

/******************* CELL 697 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell697 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[601]),
			.N(gen[602]),
			.NE(gen[603]),

			.O(gen[696]),
			.E(gen[698]),

			.SO(gen[791]),
			.S(gen[792]),
			.SE(gen[793]),

			.SELF(gen[697]),
			.cell_state(gen[697])
		); 

/******************* CELL 698 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell698 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[602]),
			.N(gen[603]),
			.NE(gen[604]),

			.O(gen[697]),
			.E(gen[699]),

			.SO(gen[792]),
			.S(gen[793]),
			.SE(gen[794]),

			.SELF(gen[698]),
			.cell_state(gen[698])
		); 

/******************* CELL 699 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell699 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[603]),
			.N(gen[604]),
			.NE(gen[605]),

			.O(gen[698]),
			.E(gen[700]),

			.SO(gen[793]),
			.S(gen[794]),
			.SE(gen[795]),

			.SELF(gen[699]),
			.cell_state(gen[699])
		); 

/******************* CELL 700 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell700 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[604]),
			.N(gen[605]),
			.NE(gen[606]),

			.O(gen[699]),
			.E(gen[701]),

			.SO(gen[794]),
			.S(gen[795]),
			.SE(gen[796]),

			.SELF(gen[700]),
			.cell_state(gen[700])
		); 

/******************* CELL 701 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell701 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[605]),
			.N(gen[606]),
			.NE(gen[607]),

			.O(gen[700]),
			.E(gen[702]),

			.SO(gen[795]),
			.S(gen[796]),
			.SE(gen[797]),

			.SELF(gen[701]),
			.cell_state(gen[701])
		); 

/******************* CELL 702 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell702 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[606]),
			.N(gen[607]),
			.NE(gen[608]),

			.O(gen[701]),
			.E(gen[703]),

			.SO(gen[796]),
			.S(gen[797]),
			.SE(gen[798]),

			.SELF(gen[702]),
			.cell_state(gen[702])
		); 

/******************* CELL 703 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell703 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[607]),
			.N(gen[608]),
			.NE(gen[609]),

			.O(gen[702]),
			.E(gen[704]),

			.SO(gen[797]),
			.S(gen[798]),
			.SE(gen[799]),

			.SELF(gen[703]),
			.cell_state(gen[703])
		); 

/******************* CELL 704 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell704 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[608]),
			.N(gen[609]),
			.NE(gen[610]),

			.O(gen[703]),
			.E(gen[705]),

			.SO(gen[798]),
			.S(gen[799]),
			.SE(gen[800]),

			.SELF(gen[704]),
			.cell_state(gen[704])
		); 

/******************* CELL 705 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell705 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[609]),
			.N(gen[610]),
			.NE(gen[611]),

			.O(gen[704]),
			.E(gen[706]),

			.SO(gen[799]),
			.S(gen[800]),
			.SE(gen[801]),

			.SELF(gen[705]),
			.cell_state(gen[705])
		); 

/******************* CELL 706 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell706 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[610]),
			.N(gen[611]),
			.NE(gen[612]),

			.O(gen[705]),
			.E(gen[707]),

			.SO(gen[800]),
			.S(gen[801]),
			.SE(gen[802]),

			.SELF(gen[706]),
			.cell_state(gen[706])
		); 

/******************* CELL 707 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell707 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[611]),
			.N(gen[612]),
			.NE(gen[613]),

			.O(gen[706]),
			.E(gen[708]),

			.SO(gen[801]),
			.S(gen[802]),
			.SE(gen[803]),

			.SELF(gen[707]),
			.cell_state(gen[707])
		); 

/******************* CELL 708 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell708 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[612]),
			.N(gen[613]),
			.NE(gen[614]),

			.O(gen[707]),
			.E(gen[709]),

			.SO(gen[802]),
			.S(gen[803]),
			.SE(gen[804]),

			.SELF(gen[708]),
			.cell_state(gen[708])
		); 

/******************* CELL 709 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell709 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[613]),
			.N(gen[614]),
			.NE(gen[615]),

			.O(gen[708]),
			.E(gen[710]),

			.SO(gen[803]),
			.S(gen[804]),
			.SE(gen[805]),

			.SELF(gen[709]),
			.cell_state(gen[709])
		); 

/******************* CELL 710 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell710 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[614]),
			.N(gen[615]),
			.NE(gen[616]),

			.O(gen[709]),
			.E(gen[711]),

			.SO(gen[804]),
			.S(gen[805]),
			.SE(gen[806]),

			.SELF(gen[710]),
			.cell_state(gen[710])
		); 

/******************* CELL 711 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell711 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[615]),
			.N(gen[616]),
			.NE(gen[617]),

			.O(gen[710]),
			.E(gen[712]),

			.SO(gen[805]),
			.S(gen[806]),
			.SE(gen[807]),

			.SELF(gen[711]),
			.cell_state(gen[711])
		); 

/******************* CELL 712 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell712 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[616]),
			.N(gen[617]),
			.NE(gen[618]),

			.O(gen[711]),
			.E(gen[713]),

			.SO(gen[806]),
			.S(gen[807]),
			.SE(gen[808]),

			.SELF(gen[712]),
			.cell_state(gen[712])
		); 

/******************* CELL 713 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell713 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[617]),
			.N(gen[618]),
			.NE(gen[619]),

			.O(gen[712]),
			.E(gen[714]),

			.SO(gen[807]),
			.S(gen[808]),
			.SE(gen[809]),

			.SELF(gen[713]),
			.cell_state(gen[713])
		); 

/******************* CELL 714 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell714 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[618]),
			.N(gen[619]),
			.NE(gen[620]),

			.O(gen[713]),
			.E(gen[715]),

			.SO(gen[808]),
			.S(gen[809]),
			.SE(gen[810]),

			.SELF(gen[714]),
			.cell_state(gen[714])
		); 

/******************* CELL 715 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell715 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[619]),
			.N(gen[620]),
			.NE(gen[621]),

			.O(gen[714]),
			.E(gen[716]),

			.SO(gen[809]),
			.S(gen[810]),
			.SE(gen[811]),

			.SELF(gen[715]),
			.cell_state(gen[715])
		); 

/******************* CELL 716 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell716 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[620]),
			.N(gen[621]),
			.NE(gen[622]),

			.O(gen[715]),
			.E(gen[717]),

			.SO(gen[810]),
			.S(gen[811]),
			.SE(gen[812]),

			.SELF(gen[716]),
			.cell_state(gen[716])
		); 

/******************* CELL 717 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell717 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[621]),
			.N(gen[622]),
			.NE(gen[623]),

			.O(gen[716]),
			.E(gen[718]),

			.SO(gen[811]),
			.S(gen[812]),
			.SE(gen[813]),

			.SELF(gen[717]),
			.cell_state(gen[717])
		); 

/******************* CELL 718 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell718 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[622]),
			.N(gen[623]),
			.NE(gen[624]),

			.O(gen[717]),
			.E(gen[719]),

			.SO(gen[812]),
			.S(gen[813]),
			.SE(gen[814]),

			.SELF(gen[718]),
			.cell_state(gen[718])
		); 

/******************* CELL 719 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell719 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[623]),
			.N(gen[624]),
			.NE(gen[625]),

			.O(gen[718]),
			.E(gen[720]),

			.SO(gen[813]),
			.S(gen[814]),
			.SE(gen[815]),

			.SELF(gen[719]),
			.cell_state(gen[719])
		); 

/******************* CELL 720 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell720 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[624]),
			.N(gen[625]),
			.NE(gen[626]),

			.O(gen[719]),
			.E(gen[721]),

			.SO(gen[814]),
			.S(gen[815]),
			.SE(gen[816]),

			.SELF(gen[720]),
			.cell_state(gen[720])
		); 

/******************* CELL 721 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell721 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[625]),
			.N(gen[626]),
			.NE(gen[627]),

			.O(gen[720]),
			.E(gen[722]),

			.SO(gen[815]),
			.S(gen[816]),
			.SE(gen[817]),

			.SELF(gen[721]),
			.cell_state(gen[721])
		); 

/******************* CELL 722 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell722 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[626]),
			.N(gen[627]),
			.NE(gen[628]),

			.O(gen[721]),
			.E(gen[723]),

			.SO(gen[816]),
			.S(gen[817]),
			.SE(gen[818]),

			.SELF(gen[722]),
			.cell_state(gen[722])
		); 

/******************* CELL 723 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell723 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[627]),
			.N(gen[628]),
			.NE(gen[629]),

			.O(gen[722]),
			.E(gen[724]),

			.SO(gen[817]),
			.S(gen[818]),
			.SE(gen[819]),

			.SELF(gen[723]),
			.cell_state(gen[723])
		); 

/******************* CELL 724 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell724 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[628]),
			.N(gen[629]),
			.NE(gen[630]),

			.O(gen[723]),
			.E(gen[725]),

			.SO(gen[818]),
			.S(gen[819]),
			.SE(gen[820]),

			.SELF(gen[724]),
			.cell_state(gen[724])
		); 

/******************* CELL 725 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell725 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[629]),
			.N(gen[630]),
			.NE(gen[631]),

			.O(gen[724]),
			.E(gen[726]),

			.SO(gen[819]),
			.S(gen[820]),
			.SE(gen[821]),

			.SELF(gen[725]),
			.cell_state(gen[725])
		); 

/******************* CELL 726 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell726 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[630]),
			.N(gen[631]),
			.NE(gen[632]),

			.O(gen[725]),
			.E(gen[727]),

			.SO(gen[820]),
			.S(gen[821]),
			.SE(gen[822]),

			.SELF(gen[726]),
			.cell_state(gen[726])
		); 

/******************* CELL 727 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell727 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[631]),
			.N(gen[632]),
			.NE(gen[633]),

			.O(gen[726]),
			.E(gen[728]),

			.SO(gen[821]),
			.S(gen[822]),
			.SE(gen[823]),

			.SELF(gen[727]),
			.cell_state(gen[727])
		); 

/******************* CELL 728 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell728 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[632]),
			.N(gen[633]),
			.NE(gen[634]),

			.O(gen[727]),
			.E(gen[729]),

			.SO(gen[822]),
			.S(gen[823]),
			.SE(gen[824]),

			.SELF(gen[728]),
			.cell_state(gen[728])
		); 

/******************* CELL 729 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell729 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[633]),
			.N(gen[634]),
			.NE(gen[635]),

			.O(gen[728]),
			.E(gen[730]),

			.SO(gen[823]),
			.S(gen[824]),
			.SE(gen[825]),

			.SELF(gen[729]),
			.cell_state(gen[729])
		); 

/******************* CELL 730 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell730 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[634]),
			.N(gen[635]),
			.NE(gen[636]),

			.O(gen[729]),
			.E(gen[731]),

			.SO(gen[824]),
			.S(gen[825]),
			.SE(gen[826]),

			.SELF(gen[730]),
			.cell_state(gen[730])
		); 

/******************* CELL 731 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell731 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[635]),
			.N(gen[636]),
			.NE(gen[637]),

			.O(gen[730]),
			.E(gen[732]),

			.SO(gen[825]),
			.S(gen[826]),
			.SE(gen[827]),

			.SELF(gen[731]),
			.cell_state(gen[731])
		); 

/******************* CELL 732 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell732 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[636]),
			.N(gen[637]),
			.NE(gen[638]),

			.O(gen[731]),
			.E(gen[733]),

			.SO(gen[826]),
			.S(gen[827]),
			.SE(gen[828]),

			.SELF(gen[732]),
			.cell_state(gen[732])
		); 

/******************* CELL 733 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell733 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[637]),
			.N(gen[638]),
			.NE(gen[639]),

			.O(gen[732]),
			.E(gen[734]),

			.SO(gen[827]),
			.S(gen[828]),
			.SE(gen[829]),

			.SELF(gen[733]),
			.cell_state(gen[733])
		); 

/******************* CELL 734 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell734 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[638]),
			.N(gen[639]),
			.NE(gen[640]),

			.O(gen[733]),
			.E(gen[735]),

			.SO(gen[828]),
			.S(gen[829]),
			.SE(gen[830]),

			.SELF(gen[734]),
			.cell_state(gen[734])
		); 

/******************* CELL 735 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell735 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[639]),
			.N(gen[640]),
			.NE(gen[641]),

			.O(gen[734]),
			.E(gen[736]),

			.SO(gen[829]),
			.S(gen[830]),
			.SE(gen[831]),

			.SELF(gen[735]),
			.cell_state(gen[735])
		); 

/******************* CELL 736 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell736 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[640]),
			.N(gen[641]),
			.NE(gen[642]),

			.O(gen[735]),
			.E(gen[737]),

			.SO(gen[830]),
			.S(gen[831]),
			.SE(gen[832]),

			.SELF(gen[736]),
			.cell_state(gen[736])
		); 

/******************* CELL 737 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell737 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[641]),
			.N(gen[642]),
			.NE(gen[643]),

			.O(gen[736]),
			.E(gen[738]),

			.SO(gen[831]),
			.S(gen[832]),
			.SE(gen[833]),

			.SELF(gen[737]),
			.cell_state(gen[737])
		); 

/******************* CELL 738 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell738 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[642]),
			.N(gen[643]),
			.NE(gen[644]),

			.O(gen[737]),
			.E(gen[739]),

			.SO(gen[832]),
			.S(gen[833]),
			.SE(gen[834]),

			.SELF(gen[738]),
			.cell_state(gen[738])
		); 

/******************* CELL 739 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell739 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[643]),
			.N(gen[644]),
			.NE(gen[645]),

			.O(gen[738]),
			.E(gen[740]),

			.SO(gen[833]),
			.S(gen[834]),
			.SE(gen[835]),

			.SELF(gen[739]),
			.cell_state(gen[739])
		); 

/******************* CELL 740 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell740 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[644]),
			.N(gen[645]),
			.NE(gen[646]),

			.O(gen[739]),
			.E(gen[741]),

			.SO(gen[834]),
			.S(gen[835]),
			.SE(gen[836]),

			.SELF(gen[740]),
			.cell_state(gen[740])
		); 

/******************* CELL 741 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell741 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[645]),
			.N(gen[646]),
			.NE(gen[647]),

			.O(gen[740]),
			.E(gen[742]),

			.SO(gen[835]),
			.S(gen[836]),
			.SE(gen[837]),

			.SELF(gen[741]),
			.cell_state(gen[741])
		); 

/******************* CELL 742 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell742 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[646]),
			.N(gen[647]),
			.NE(gen[648]),

			.O(gen[741]),
			.E(gen[743]),

			.SO(gen[836]),
			.S(gen[837]),
			.SE(gen[838]),

			.SELF(gen[742]),
			.cell_state(gen[742])
		); 

/******************* CELL 743 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell743 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[647]),
			.N(gen[648]),
			.NE(gen[649]),

			.O(gen[742]),
			.E(gen[744]),

			.SO(gen[837]),
			.S(gen[838]),
			.SE(gen[839]),

			.SELF(gen[743]),
			.cell_state(gen[743])
		); 

/******************* CELL 744 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell744 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[648]),
			.N(gen[649]),
			.NE(gen[650]),

			.O(gen[743]),
			.E(gen[745]),

			.SO(gen[838]),
			.S(gen[839]),
			.SE(gen[840]),

			.SELF(gen[744]),
			.cell_state(gen[744])
		); 

/******************* CELL 745 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell745 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[649]),
			.N(gen[650]),
			.NE(gen[651]),

			.O(gen[744]),
			.E(gen[746]),

			.SO(gen[839]),
			.S(gen[840]),
			.SE(gen[841]),

			.SELF(gen[745]),
			.cell_state(gen[745])
		); 

/******************* CELL 746 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell746 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[650]),
			.N(gen[651]),
			.NE(gen[652]),

			.O(gen[745]),
			.E(gen[747]),

			.SO(gen[840]),
			.S(gen[841]),
			.SE(gen[842]),

			.SELF(gen[746]),
			.cell_state(gen[746])
		); 

/******************* CELL 747 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell747 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[651]),
			.N(gen[652]),
			.NE(gen[653]),

			.O(gen[746]),
			.E(gen[748]),

			.SO(gen[841]),
			.S(gen[842]),
			.SE(gen[843]),

			.SELF(gen[747]),
			.cell_state(gen[747])
		); 

/******************* CELL 748 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell748 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[652]),
			.N(gen[653]),
			.NE(gen[654]),

			.O(gen[747]),
			.E(gen[749]),

			.SO(gen[842]),
			.S(gen[843]),
			.SE(gen[844]),

			.SELF(gen[748]),
			.cell_state(gen[748])
		); 

/******************* CELL 749 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell749 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[653]),
			.N(gen[654]),
			.NE(gen[655]),

			.O(gen[748]),
			.E(gen[750]),

			.SO(gen[843]),
			.S(gen[844]),
			.SE(gen[845]),

			.SELF(gen[749]),
			.cell_state(gen[749])
		); 

/******************* CELL 750 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell750 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[654]),
			.N(gen[655]),
			.NE(gen[656]),

			.O(gen[749]),
			.E(gen[751]),

			.SO(gen[844]),
			.S(gen[845]),
			.SE(gen[846]),

			.SELF(gen[750]),
			.cell_state(gen[750])
		); 

/******************* CELL 751 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell751 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[655]),
			.N(gen[656]),
			.NE(gen[657]),

			.O(gen[750]),
			.E(gen[752]),

			.SO(gen[845]),
			.S(gen[846]),
			.SE(gen[847]),

			.SELF(gen[751]),
			.cell_state(gen[751])
		); 

/******************* CELL 752 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell752 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[656]),
			.N(gen[657]),
			.NE(gen[658]),

			.O(gen[751]),
			.E(gen[753]),

			.SO(gen[846]),
			.S(gen[847]),
			.SE(gen[848]),

			.SELF(gen[752]),
			.cell_state(gen[752])
		); 

/******************* CELL 753 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell753 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[657]),
			.N(gen[658]),
			.NE(gen[659]),

			.O(gen[752]),
			.E(gen[754]),

			.SO(gen[847]),
			.S(gen[848]),
			.SE(gen[849]),

			.SELF(gen[753]),
			.cell_state(gen[753])
		); 

/******************* CELL 754 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell754 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[658]),
			.N(gen[659]),
			.NE(gen[660]),

			.O(gen[753]),
			.E(gen[755]),

			.SO(gen[848]),
			.S(gen[849]),
			.SE(gen[850]),

			.SELF(gen[754]),
			.cell_state(gen[754])
		); 

/******************* CELL 755 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell755 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[659]),
			.N(gen[660]),
			.NE(gen[661]),

			.O(gen[754]),
			.E(gen[756]),

			.SO(gen[849]),
			.S(gen[850]),
			.SE(gen[851]),

			.SELF(gen[755]),
			.cell_state(gen[755])
		); 

/******************* CELL 756 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell756 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[660]),
			.N(gen[661]),
			.NE(gen[662]),

			.O(gen[755]),
			.E(gen[757]),

			.SO(gen[850]),
			.S(gen[851]),
			.SE(gen[852]),

			.SELF(gen[756]),
			.cell_state(gen[756])
		); 

/******************* CELL 757 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell757 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[661]),
			.N(gen[662]),
			.NE(gen[663]),

			.O(gen[756]),
			.E(gen[758]),

			.SO(gen[851]),
			.S(gen[852]),
			.SE(gen[853]),

			.SELF(gen[757]),
			.cell_state(gen[757])
		); 

/******************* CELL 758 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell758 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[662]),
			.N(gen[663]),
			.NE(gen[664]),

			.O(gen[757]),
			.E(gen[759]),

			.SO(gen[852]),
			.S(gen[853]),
			.SE(gen[854]),

			.SELF(gen[758]),
			.cell_state(gen[758])
		); 

/******************* CELL 759 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell759 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[663]),
			.N(gen[664]),
			.NE(gen[663]),

			.O(gen[758]),
			.E(gen[758]),

			.SO(gen[853]),
			.S(gen[854]),
			.SE(gen[853]),

			.SELF(gen[759]),
			.cell_state(gen[759])
		); 

/******************* CELL 760 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell760 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[666]),
			.N(gen[665]),
			.NE(gen[666]),

			.O(gen[761]),
			.E(gen[761]),

			.SO(gen[856]),
			.S(gen[855]),
			.SE(gen[856]),

			.SELF(gen[760]),
			.cell_state(gen[760])
		); 

/******************* CELL 761 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell761 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[665]),
			.N(gen[666]),
			.NE(gen[667]),

			.O(gen[760]),
			.E(gen[762]),

			.SO(gen[855]),
			.S(gen[856]),
			.SE(gen[857]),

			.SELF(gen[761]),
			.cell_state(gen[761])
		); 

/******************* CELL 762 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell762 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[666]),
			.N(gen[667]),
			.NE(gen[668]),

			.O(gen[761]),
			.E(gen[763]),

			.SO(gen[856]),
			.S(gen[857]),
			.SE(gen[858]),

			.SELF(gen[762]),
			.cell_state(gen[762])
		); 

/******************* CELL 763 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell763 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[667]),
			.N(gen[668]),
			.NE(gen[669]),

			.O(gen[762]),
			.E(gen[764]),

			.SO(gen[857]),
			.S(gen[858]),
			.SE(gen[859]),

			.SELF(gen[763]),
			.cell_state(gen[763])
		); 

/******************* CELL 764 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell764 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[668]),
			.N(gen[669]),
			.NE(gen[670]),

			.O(gen[763]),
			.E(gen[765]),

			.SO(gen[858]),
			.S(gen[859]),
			.SE(gen[860]),

			.SELF(gen[764]),
			.cell_state(gen[764])
		); 

/******************* CELL 765 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell765 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[669]),
			.N(gen[670]),
			.NE(gen[671]),

			.O(gen[764]),
			.E(gen[766]),

			.SO(gen[859]),
			.S(gen[860]),
			.SE(gen[861]),

			.SELF(gen[765]),
			.cell_state(gen[765])
		); 

/******************* CELL 766 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell766 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[670]),
			.N(gen[671]),
			.NE(gen[672]),

			.O(gen[765]),
			.E(gen[767]),

			.SO(gen[860]),
			.S(gen[861]),
			.SE(gen[862]),

			.SELF(gen[766]),
			.cell_state(gen[766])
		); 

/******************* CELL 767 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell767 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[671]),
			.N(gen[672]),
			.NE(gen[673]),

			.O(gen[766]),
			.E(gen[768]),

			.SO(gen[861]),
			.S(gen[862]),
			.SE(gen[863]),

			.SELF(gen[767]),
			.cell_state(gen[767])
		); 

/******************* CELL 768 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell768 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[672]),
			.N(gen[673]),
			.NE(gen[674]),

			.O(gen[767]),
			.E(gen[769]),

			.SO(gen[862]),
			.S(gen[863]),
			.SE(gen[864]),

			.SELF(gen[768]),
			.cell_state(gen[768])
		); 

/******************* CELL 769 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell769 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[673]),
			.N(gen[674]),
			.NE(gen[675]),

			.O(gen[768]),
			.E(gen[770]),

			.SO(gen[863]),
			.S(gen[864]),
			.SE(gen[865]),

			.SELF(gen[769]),
			.cell_state(gen[769])
		); 

/******************* CELL 770 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell770 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[674]),
			.N(gen[675]),
			.NE(gen[676]),

			.O(gen[769]),
			.E(gen[771]),

			.SO(gen[864]),
			.S(gen[865]),
			.SE(gen[866]),

			.SELF(gen[770]),
			.cell_state(gen[770])
		); 

/******************* CELL 771 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell771 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[675]),
			.N(gen[676]),
			.NE(gen[677]),

			.O(gen[770]),
			.E(gen[772]),

			.SO(gen[865]),
			.S(gen[866]),
			.SE(gen[867]),

			.SELF(gen[771]),
			.cell_state(gen[771])
		); 

/******************* CELL 772 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell772 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[676]),
			.N(gen[677]),
			.NE(gen[678]),

			.O(gen[771]),
			.E(gen[773]),

			.SO(gen[866]),
			.S(gen[867]),
			.SE(gen[868]),

			.SELF(gen[772]),
			.cell_state(gen[772])
		); 

/******************* CELL 773 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell773 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[677]),
			.N(gen[678]),
			.NE(gen[679]),

			.O(gen[772]),
			.E(gen[774]),

			.SO(gen[867]),
			.S(gen[868]),
			.SE(gen[869]),

			.SELF(gen[773]),
			.cell_state(gen[773])
		); 

/******************* CELL 774 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell774 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[678]),
			.N(gen[679]),
			.NE(gen[680]),

			.O(gen[773]),
			.E(gen[775]),

			.SO(gen[868]),
			.S(gen[869]),
			.SE(gen[870]),

			.SELF(gen[774]),
			.cell_state(gen[774])
		); 

/******************* CELL 775 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell775 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[679]),
			.N(gen[680]),
			.NE(gen[681]),

			.O(gen[774]),
			.E(gen[776]),

			.SO(gen[869]),
			.S(gen[870]),
			.SE(gen[871]),

			.SELF(gen[775]),
			.cell_state(gen[775])
		); 

/******************* CELL 776 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell776 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[680]),
			.N(gen[681]),
			.NE(gen[682]),

			.O(gen[775]),
			.E(gen[777]),

			.SO(gen[870]),
			.S(gen[871]),
			.SE(gen[872]),

			.SELF(gen[776]),
			.cell_state(gen[776])
		); 

/******************* CELL 777 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell777 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[681]),
			.N(gen[682]),
			.NE(gen[683]),

			.O(gen[776]),
			.E(gen[778]),

			.SO(gen[871]),
			.S(gen[872]),
			.SE(gen[873]),

			.SELF(gen[777]),
			.cell_state(gen[777])
		); 

/******************* CELL 778 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell778 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[682]),
			.N(gen[683]),
			.NE(gen[684]),

			.O(gen[777]),
			.E(gen[779]),

			.SO(gen[872]),
			.S(gen[873]),
			.SE(gen[874]),

			.SELF(gen[778]),
			.cell_state(gen[778])
		); 

/******************* CELL 779 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell779 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[683]),
			.N(gen[684]),
			.NE(gen[685]),

			.O(gen[778]),
			.E(gen[780]),

			.SO(gen[873]),
			.S(gen[874]),
			.SE(gen[875]),

			.SELF(gen[779]),
			.cell_state(gen[779])
		); 

/******************* CELL 780 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell780 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[684]),
			.N(gen[685]),
			.NE(gen[686]),

			.O(gen[779]),
			.E(gen[781]),

			.SO(gen[874]),
			.S(gen[875]),
			.SE(gen[876]),

			.SELF(gen[780]),
			.cell_state(gen[780])
		); 

/******************* CELL 781 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell781 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[685]),
			.N(gen[686]),
			.NE(gen[687]),

			.O(gen[780]),
			.E(gen[782]),

			.SO(gen[875]),
			.S(gen[876]),
			.SE(gen[877]),

			.SELF(gen[781]),
			.cell_state(gen[781])
		); 

/******************* CELL 782 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell782 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[686]),
			.N(gen[687]),
			.NE(gen[688]),

			.O(gen[781]),
			.E(gen[783]),

			.SO(gen[876]),
			.S(gen[877]),
			.SE(gen[878]),

			.SELF(gen[782]),
			.cell_state(gen[782])
		); 

/******************* CELL 783 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell783 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[687]),
			.N(gen[688]),
			.NE(gen[689]),

			.O(gen[782]),
			.E(gen[784]),

			.SO(gen[877]),
			.S(gen[878]),
			.SE(gen[879]),

			.SELF(gen[783]),
			.cell_state(gen[783])
		); 

/******************* CELL 784 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell784 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[688]),
			.N(gen[689]),
			.NE(gen[690]),

			.O(gen[783]),
			.E(gen[785]),

			.SO(gen[878]),
			.S(gen[879]),
			.SE(gen[880]),

			.SELF(gen[784]),
			.cell_state(gen[784])
		); 

/******************* CELL 785 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell785 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[689]),
			.N(gen[690]),
			.NE(gen[691]),

			.O(gen[784]),
			.E(gen[786]),

			.SO(gen[879]),
			.S(gen[880]),
			.SE(gen[881]),

			.SELF(gen[785]),
			.cell_state(gen[785])
		); 

/******************* CELL 786 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell786 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[690]),
			.N(gen[691]),
			.NE(gen[692]),

			.O(gen[785]),
			.E(gen[787]),

			.SO(gen[880]),
			.S(gen[881]),
			.SE(gen[882]),

			.SELF(gen[786]),
			.cell_state(gen[786])
		); 

/******************* CELL 787 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell787 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[691]),
			.N(gen[692]),
			.NE(gen[693]),

			.O(gen[786]),
			.E(gen[788]),

			.SO(gen[881]),
			.S(gen[882]),
			.SE(gen[883]),

			.SELF(gen[787]),
			.cell_state(gen[787])
		); 

/******************* CELL 788 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell788 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[692]),
			.N(gen[693]),
			.NE(gen[694]),

			.O(gen[787]),
			.E(gen[789]),

			.SO(gen[882]),
			.S(gen[883]),
			.SE(gen[884]),

			.SELF(gen[788]),
			.cell_state(gen[788])
		); 

/******************* CELL 789 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell789 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[693]),
			.N(gen[694]),
			.NE(gen[695]),

			.O(gen[788]),
			.E(gen[790]),

			.SO(gen[883]),
			.S(gen[884]),
			.SE(gen[885]),

			.SELF(gen[789]),
			.cell_state(gen[789])
		); 

/******************* CELL 790 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell790 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[694]),
			.N(gen[695]),
			.NE(gen[696]),

			.O(gen[789]),
			.E(gen[791]),

			.SO(gen[884]),
			.S(gen[885]),
			.SE(gen[886]),

			.SELF(gen[790]),
			.cell_state(gen[790])
		); 

/******************* CELL 791 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell791 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[695]),
			.N(gen[696]),
			.NE(gen[697]),

			.O(gen[790]),
			.E(gen[792]),

			.SO(gen[885]),
			.S(gen[886]),
			.SE(gen[887]),

			.SELF(gen[791]),
			.cell_state(gen[791])
		); 

/******************* CELL 792 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell792 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[696]),
			.N(gen[697]),
			.NE(gen[698]),

			.O(gen[791]),
			.E(gen[793]),

			.SO(gen[886]),
			.S(gen[887]),
			.SE(gen[888]),

			.SELF(gen[792]),
			.cell_state(gen[792])
		); 

/******************* CELL 793 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell793 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[697]),
			.N(gen[698]),
			.NE(gen[699]),

			.O(gen[792]),
			.E(gen[794]),

			.SO(gen[887]),
			.S(gen[888]),
			.SE(gen[889]),

			.SELF(gen[793]),
			.cell_state(gen[793])
		); 

/******************* CELL 794 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell794 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[698]),
			.N(gen[699]),
			.NE(gen[700]),

			.O(gen[793]),
			.E(gen[795]),

			.SO(gen[888]),
			.S(gen[889]),
			.SE(gen[890]),

			.SELF(gen[794]),
			.cell_state(gen[794])
		); 

/******************* CELL 795 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell795 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[699]),
			.N(gen[700]),
			.NE(gen[701]),

			.O(gen[794]),
			.E(gen[796]),

			.SO(gen[889]),
			.S(gen[890]),
			.SE(gen[891]),

			.SELF(gen[795]),
			.cell_state(gen[795])
		); 

/******************* CELL 796 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell796 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[700]),
			.N(gen[701]),
			.NE(gen[702]),

			.O(gen[795]),
			.E(gen[797]),

			.SO(gen[890]),
			.S(gen[891]),
			.SE(gen[892]),

			.SELF(gen[796]),
			.cell_state(gen[796])
		); 

/******************* CELL 797 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell797 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[701]),
			.N(gen[702]),
			.NE(gen[703]),

			.O(gen[796]),
			.E(gen[798]),

			.SO(gen[891]),
			.S(gen[892]),
			.SE(gen[893]),

			.SELF(gen[797]),
			.cell_state(gen[797])
		); 

/******************* CELL 798 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell798 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[702]),
			.N(gen[703]),
			.NE(gen[704]),

			.O(gen[797]),
			.E(gen[799]),

			.SO(gen[892]),
			.S(gen[893]),
			.SE(gen[894]),

			.SELF(gen[798]),
			.cell_state(gen[798])
		); 

/******************* CELL 799 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell799 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[703]),
			.N(gen[704]),
			.NE(gen[705]),

			.O(gen[798]),
			.E(gen[800]),

			.SO(gen[893]),
			.S(gen[894]),
			.SE(gen[895]),

			.SELF(gen[799]),
			.cell_state(gen[799])
		); 

/******************* CELL 800 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell800 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[704]),
			.N(gen[705]),
			.NE(gen[706]),

			.O(gen[799]),
			.E(gen[801]),

			.SO(gen[894]),
			.S(gen[895]),
			.SE(gen[896]),

			.SELF(gen[800]),
			.cell_state(gen[800])
		); 

/******************* CELL 801 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell801 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[705]),
			.N(gen[706]),
			.NE(gen[707]),

			.O(gen[800]),
			.E(gen[802]),

			.SO(gen[895]),
			.S(gen[896]),
			.SE(gen[897]),

			.SELF(gen[801]),
			.cell_state(gen[801])
		); 

/******************* CELL 802 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell802 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[706]),
			.N(gen[707]),
			.NE(gen[708]),

			.O(gen[801]),
			.E(gen[803]),

			.SO(gen[896]),
			.S(gen[897]),
			.SE(gen[898]),

			.SELF(gen[802]),
			.cell_state(gen[802])
		); 

/******************* CELL 803 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell803 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[707]),
			.N(gen[708]),
			.NE(gen[709]),

			.O(gen[802]),
			.E(gen[804]),

			.SO(gen[897]),
			.S(gen[898]),
			.SE(gen[899]),

			.SELF(gen[803]),
			.cell_state(gen[803])
		); 

/******************* CELL 804 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell804 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[708]),
			.N(gen[709]),
			.NE(gen[710]),

			.O(gen[803]),
			.E(gen[805]),

			.SO(gen[898]),
			.S(gen[899]),
			.SE(gen[900]),

			.SELF(gen[804]),
			.cell_state(gen[804])
		); 

/******************* CELL 805 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell805 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[709]),
			.N(gen[710]),
			.NE(gen[711]),

			.O(gen[804]),
			.E(gen[806]),

			.SO(gen[899]),
			.S(gen[900]),
			.SE(gen[901]),

			.SELF(gen[805]),
			.cell_state(gen[805])
		); 

/******************* CELL 806 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell806 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[710]),
			.N(gen[711]),
			.NE(gen[712]),

			.O(gen[805]),
			.E(gen[807]),

			.SO(gen[900]),
			.S(gen[901]),
			.SE(gen[902]),

			.SELF(gen[806]),
			.cell_state(gen[806])
		); 

/******************* CELL 807 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell807 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[711]),
			.N(gen[712]),
			.NE(gen[713]),

			.O(gen[806]),
			.E(gen[808]),

			.SO(gen[901]),
			.S(gen[902]),
			.SE(gen[903]),

			.SELF(gen[807]),
			.cell_state(gen[807])
		); 

/******************* CELL 808 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell808 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[712]),
			.N(gen[713]),
			.NE(gen[714]),

			.O(gen[807]),
			.E(gen[809]),

			.SO(gen[902]),
			.S(gen[903]),
			.SE(gen[904]),

			.SELF(gen[808]),
			.cell_state(gen[808])
		); 

/******************* CELL 809 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell809 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[713]),
			.N(gen[714]),
			.NE(gen[715]),

			.O(gen[808]),
			.E(gen[810]),

			.SO(gen[903]),
			.S(gen[904]),
			.SE(gen[905]),

			.SELF(gen[809]),
			.cell_state(gen[809])
		); 

/******************* CELL 810 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell810 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[714]),
			.N(gen[715]),
			.NE(gen[716]),

			.O(gen[809]),
			.E(gen[811]),

			.SO(gen[904]),
			.S(gen[905]),
			.SE(gen[906]),

			.SELF(gen[810]),
			.cell_state(gen[810])
		); 

/******************* CELL 811 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell811 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[715]),
			.N(gen[716]),
			.NE(gen[717]),

			.O(gen[810]),
			.E(gen[812]),

			.SO(gen[905]),
			.S(gen[906]),
			.SE(gen[907]),

			.SELF(gen[811]),
			.cell_state(gen[811])
		); 

/******************* CELL 812 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell812 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[716]),
			.N(gen[717]),
			.NE(gen[718]),

			.O(gen[811]),
			.E(gen[813]),

			.SO(gen[906]),
			.S(gen[907]),
			.SE(gen[908]),

			.SELF(gen[812]),
			.cell_state(gen[812])
		); 

/******************* CELL 813 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell813 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[717]),
			.N(gen[718]),
			.NE(gen[719]),

			.O(gen[812]),
			.E(gen[814]),

			.SO(gen[907]),
			.S(gen[908]),
			.SE(gen[909]),

			.SELF(gen[813]),
			.cell_state(gen[813])
		); 

/******************* CELL 814 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell814 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[718]),
			.N(gen[719]),
			.NE(gen[720]),

			.O(gen[813]),
			.E(gen[815]),

			.SO(gen[908]),
			.S(gen[909]),
			.SE(gen[910]),

			.SELF(gen[814]),
			.cell_state(gen[814])
		); 

/******************* CELL 815 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell815 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[719]),
			.N(gen[720]),
			.NE(gen[721]),

			.O(gen[814]),
			.E(gen[816]),

			.SO(gen[909]),
			.S(gen[910]),
			.SE(gen[911]),

			.SELF(gen[815]),
			.cell_state(gen[815])
		); 

/******************* CELL 816 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell816 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[720]),
			.N(gen[721]),
			.NE(gen[722]),

			.O(gen[815]),
			.E(gen[817]),

			.SO(gen[910]),
			.S(gen[911]),
			.SE(gen[912]),

			.SELF(gen[816]),
			.cell_state(gen[816])
		); 

/******************* CELL 817 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell817 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[721]),
			.N(gen[722]),
			.NE(gen[723]),

			.O(gen[816]),
			.E(gen[818]),

			.SO(gen[911]),
			.S(gen[912]),
			.SE(gen[913]),

			.SELF(gen[817]),
			.cell_state(gen[817])
		); 

/******************* CELL 818 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell818 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[722]),
			.N(gen[723]),
			.NE(gen[724]),

			.O(gen[817]),
			.E(gen[819]),

			.SO(gen[912]),
			.S(gen[913]),
			.SE(gen[914]),

			.SELF(gen[818]),
			.cell_state(gen[818])
		); 

/******************* CELL 819 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell819 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[723]),
			.N(gen[724]),
			.NE(gen[725]),

			.O(gen[818]),
			.E(gen[820]),

			.SO(gen[913]),
			.S(gen[914]),
			.SE(gen[915]),

			.SELF(gen[819]),
			.cell_state(gen[819])
		); 

/******************* CELL 820 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell820 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[724]),
			.N(gen[725]),
			.NE(gen[726]),

			.O(gen[819]),
			.E(gen[821]),

			.SO(gen[914]),
			.S(gen[915]),
			.SE(gen[916]),

			.SELF(gen[820]),
			.cell_state(gen[820])
		); 

/******************* CELL 821 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell821 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[725]),
			.N(gen[726]),
			.NE(gen[727]),

			.O(gen[820]),
			.E(gen[822]),

			.SO(gen[915]),
			.S(gen[916]),
			.SE(gen[917]),

			.SELF(gen[821]),
			.cell_state(gen[821])
		); 

/******************* CELL 822 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell822 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[726]),
			.N(gen[727]),
			.NE(gen[728]),

			.O(gen[821]),
			.E(gen[823]),

			.SO(gen[916]),
			.S(gen[917]),
			.SE(gen[918]),

			.SELF(gen[822]),
			.cell_state(gen[822])
		); 

/******************* CELL 823 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell823 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[727]),
			.N(gen[728]),
			.NE(gen[729]),

			.O(gen[822]),
			.E(gen[824]),

			.SO(gen[917]),
			.S(gen[918]),
			.SE(gen[919]),

			.SELF(gen[823]),
			.cell_state(gen[823])
		); 

/******************* CELL 824 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell824 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[728]),
			.N(gen[729]),
			.NE(gen[730]),

			.O(gen[823]),
			.E(gen[825]),

			.SO(gen[918]),
			.S(gen[919]),
			.SE(gen[920]),

			.SELF(gen[824]),
			.cell_state(gen[824])
		); 

/******************* CELL 825 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell825 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[729]),
			.N(gen[730]),
			.NE(gen[731]),

			.O(gen[824]),
			.E(gen[826]),

			.SO(gen[919]),
			.S(gen[920]),
			.SE(gen[921]),

			.SELF(gen[825]),
			.cell_state(gen[825])
		); 

/******************* CELL 826 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell826 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[730]),
			.N(gen[731]),
			.NE(gen[732]),

			.O(gen[825]),
			.E(gen[827]),

			.SO(gen[920]),
			.S(gen[921]),
			.SE(gen[922]),

			.SELF(gen[826]),
			.cell_state(gen[826])
		); 

/******************* CELL 827 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell827 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[731]),
			.N(gen[732]),
			.NE(gen[733]),

			.O(gen[826]),
			.E(gen[828]),

			.SO(gen[921]),
			.S(gen[922]),
			.SE(gen[923]),

			.SELF(gen[827]),
			.cell_state(gen[827])
		); 

/******************* CELL 828 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell828 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[732]),
			.N(gen[733]),
			.NE(gen[734]),

			.O(gen[827]),
			.E(gen[829]),

			.SO(gen[922]),
			.S(gen[923]),
			.SE(gen[924]),

			.SELF(gen[828]),
			.cell_state(gen[828])
		); 

/******************* CELL 829 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell829 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[733]),
			.N(gen[734]),
			.NE(gen[735]),

			.O(gen[828]),
			.E(gen[830]),

			.SO(gen[923]),
			.S(gen[924]),
			.SE(gen[925]),

			.SELF(gen[829]),
			.cell_state(gen[829])
		); 

/******************* CELL 830 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell830 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[734]),
			.N(gen[735]),
			.NE(gen[736]),

			.O(gen[829]),
			.E(gen[831]),

			.SO(gen[924]),
			.S(gen[925]),
			.SE(gen[926]),

			.SELF(gen[830]),
			.cell_state(gen[830])
		); 

/******************* CELL 831 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell831 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[735]),
			.N(gen[736]),
			.NE(gen[737]),

			.O(gen[830]),
			.E(gen[832]),

			.SO(gen[925]),
			.S(gen[926]),
			.SE(gen[927]),

			.SELF(gen[831]),
			.cell_state(gen[831])
		); 

/******************* CELL 832 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell832 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[736]),
			.N(gen[737]),
			.NE(gen[738]),

			.O(gen[831]),
			.E(gen[833]),

			.SO(gen[926]),
			.S(gen[927]),
			.SE(gen[928]),

			.SELF(gen[832]),
			.cell_state(gen[832])
		); 

/******************* CELL 833 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell833 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[737]),
			.N(gen[738]),
			.NE(gen[739]),

			.O(gen[832]),
			.E(gen[834]),

			.SO(gen[927]),
			.S(gen[928]),
			.SE(gen[929]),

			.SELF(gen[833]),
			.cell_state(gen[833])
		); 

/******************* CELL 834 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell834 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[738]),
			.N(gen[739]),
			.NE(gen[740]),

			.O(gen[833]),
			.E(gen[835]),

			.SO(gen[928]),
			.S(gen[929]),
			.SE(gen[930]),

			.SELF(gen[834]),
			.cell_state(gen[834])
		); 

/******************* CELL 835 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell835 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[739]),
			.N(gen[740]),
			.NE(gen[741]),

			.O(gen[834]),
			.E(gen[836]),

			.SO(gen[929]),
			.S(gen[930]),
			.SE(gen[931]),

			.SELF(gen[835]),
			.cell_state(gen[835])
		); 

/******************* CELL 836 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell836 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[740]),
			.N(gen[741]),
			.NE(gen[742]),

			.O(gen[835]),
			.E(gen[837]),

			.SO(gen[930]),
			.S(gen[931]),
			.SE(gen[932]),

			.SELF(gen[836]),
			.cell_state(gen[836])
		); 

/******************* CELL 837 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell837 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[741]),
			.N(gen[742]),
			.NE(gen[743]),

			.O(gen[836]),
			.E(gen[838]),

			.SO(gen[931]),
			.S(gen[932]),
			.SE(gen[933]),

			.SELF(gen[837]),
			.cell_state(gen[837])
		); 

/******************* CELL 838 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell838 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[742]),
			.N(gen[743]),
			.NE(gen[744]),

			.O(gen[837]),
			.E(gen[839]),

			.SO(gen[932]),
			.S(gen[933]),
			.SE(gen[934]),

			.SELF(gen[838]),
			.cell_state(gen[838])
		); 

/******************* CELL 839 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell839 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[743]),
			.N(gen[744]),
			.NE(gen[745]),

			.O(gen[838]),
			.E(gen[840]),

			.SO(gen[933]),
			.S(gen[934]),
			.SE(gen[935]),

			.SELF(gen[839]),
			.cell_state(gen[839])
		); 

/******************* CELL 840 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell840 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[744]),
			.N(gen[745]),
			.NE(gen[746]),

			.O(gen[839]),
			.E(gen[841]),

			.SO(gen[934]),
			.S(gen[935]),
			.SE(gen[936]),

			.SELF(gen[840]),
			.cell_state(gen[840])
		); 

/******************* CELL 841 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell841 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[745]),
			.N(gen[746]),
			.NE(gen[747]),

			.O(gen[840]),
			.E(gen[842]),

			.SO(gen[935]),
			.S(gen[936]),
			.SE(gen[937]),

			.SELF(gen[841]),
			.cell_state(gen[841])
		); 

/******************* CELL 842 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell842 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[746]),
			.N(gen[747]),
			.NE(gen[748]),

			.O(gen[841]),
			.E(gen[843]),

			.SO(gen[936]),
			.S(gen[937]),
			.SE(gen[938]),

			.SELF(gen[842]),
			.cell_state(gen[842])
		); 

/******************* CELL 843 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell843 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[747]),
			.N(gen[748]),
			.NE(gen[749]),

			.O(gen[842]),
			.E(gen[844]),

			.SO(gen[937]),
			.S(gen[938]),
			.SE(gen[939]),

			.SELF(gen[843]),
			.cell_state(gen[843])
		); 

/******************* CELL 844 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell844 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[748]),
			.N(gen[749]),
			.NE(gen[750]),

			.O(gen[843]),
			.E(gen[845]),

			.SO(gen[938]),
			.S(gen[939]),
			.SE(gen[940]),

			.SELF(gen[844]),
			.cell_state(gen[844])
		); 

/******************* CELL 845 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell845 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[749]),
			.N(gen[750]),
			.NE(gen[751]),

			.O(gen[844]),
			.E(gen[846]),

			.SO(gen[939]),
			.S(gen[940]),
			.SE(gen[941]),

			.SELF(gen[845]),
			.cell_state(gen[845])
		); 

/******************* CELL 846 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell846 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[750]),
			.N(gen[751]),
			.NE(gen[752]),

			.O(gen[845]),
			.E(gen[847]),

			.SO(gen[940]),
			.S(gen[941]),
			.SE(gen[942]),

			.SELF(gen[846]),
			.cell_state(gen[846])
		); 

/******************* CELL 847 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell847 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[751]),
			.N(gen[752]),
			.NE(gen[753]),

			.O(gen[846]),
			.E(gen[848]),

			.SO(gen[941]),
			.S(gen[942]),
			.SE(gen[943]),

			.SELF(gen[847]),
			.cell_state(gen[847])
		); 

/******************* CELL 848 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell848 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[752]),
			.N(gen[753]),
			.NE(gen[754]),

			.O(gen[847]),
			.E(gen[849]),

			.SO(gen[942]),
			.S(gen[943]),
			.SE(gen[944]),

			.SELF(gen[848]),
			.cell_state(gen[848])
		); 

/******************* CELL 849 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell849 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[753]),
			.N(gen[754]),
			.NE(gen[755]),

			.O(gen[848]),
			.E(gen[850]),

			.SO(gen[943]),
			.S(gen[944]),
			.SE(gen[945]),

			.SELF(gen[849]),
			.cell_state(gen[849])
		); 

/******************* CELL 850 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell850 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[754]),
			.N(gen[755]),
			.NE(gen[756]),

			.O(gen[849]),
			.E(gen[851]),

			.SO(gen[944]),
			.S(gen[945]),
			.SE(gen[946]),

			.SELF(gen[850]),
			.cell_state(gen[850])
		); 

/******************* CELL 851 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell851 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[755]),
			.N(gen[756]),
			.NE(gen[757]),

			.O(gen[850]),
			.E(gen[852]),

			.SO(gen[945]),
			.S(gen[946]),
			.SE(gen[947]),

			.SELF(gen[851]),
			.cell_state(gen[851])
		); 

/******************* CELL 852 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell852 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[756]),
			.N(gen[757]),
			.NE(gen[758]),

			.O(gen[851]),
			.E(gen[853]),

			.SO(gen[946]),
			.S(gen[947]),
			.SE(gen[948]),

			.SELF(gen[852]),
			.cell_state(gen[852])
		); 

/******************* CELL 853 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell853 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[757]),
			.N(gen[758]),
			.NE(gen[759]),

			.O(gen[852]),
			.E(gen[854]),

			.SO(gen[947]),
			.S(gen[948]),
			.SE(gen[949]),

			.SELF(gen[853]),
			.cell_state(gen[853])
		); 

/******************* CELL 854 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell854 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[758]),
			.N(gen[759]),
			.NE(gen[758]),

			.O(gen[853]),
			.E(gen[853]),

			.SO(gen[948]),
			.S(gen[949]),
			.SE(gen[948]),

			.SELF(gen[854]),
			.cell_state(gen[854])
		); 

/******************* CELL 855 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell855 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[761]),
			.N(gen[760]),
			.NE(gen[761]),

			.O(gen[856]),
			.E(gen[856]),

			.SO(gen[951]),
			.S(gen[950]),
			.SE(gen[951]),

			.SELF(gen[855]),
			.cell_state(gen[855])
		); 

/******************* CELL 856 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell856 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[760]),
			.N(gen[761]),
			.NE(gen[762]),

			.O(gen[855]),
			.E(gen[857]),

			.SO(gen[950]),
			.S(gen[951]),
			.SE(gen[952]),

			.SELF(gen[856]),
			.cell_state(gen[856])
		); 

/******************* CELL 857 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell857 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[761]),
			.N(gen[762]),
			.NE(gen[763]),

			.O(gen[856]),
			.E(gen[858]),

			.SO(gen[951]),
			.S(gen[952]),
			.SE(gen[953]),

			.SELF(gen[857]),
			.cell_state(gen[857])
		); 

/******************* CELL 858 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell858 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[762]),
			.N(gen[763]),
			.NE(gen[764]),

			.O(gen[857]),
			.E(gen[859]),

			.SO(gen[952]),
			.S(gen[953]),
			.SE(gen[954]),

			.SELF(gen[858]),
			.cell_state(gen[858])
		); 

/******************* CELL 859 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell859 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[763]),
			.N(gen[764]),
			.NE(gen[765]),

			.O(gen[858]),
			.E(gen[860]),

			.SO(gen[953]),
			.S(gen[954]),
			.SE(gen[955]),

			.SELF(gen[859]),
			.cell_state(gen[859])
		); 

/******************* CELL 860 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell860 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[764]),
			.N(gen[765]),
			.NE(gen[766]),

			.O(gen[859]),
			.E(gen[861]),

			.SO(gen[954]),
			.S(gen[955]),
			.SE(gen[956]),

			.SELF(gen[860]),
			.cell_state(gen[860])
		); 

/******************* CELL 861 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell861 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[765]),
			.N(gen[766]),
			.NE(gen[767]),

			.O(gen[860]),
			.E(gen[862]),

			.SO(gen[955]),
			.S(gen[956]),
			.SE(gen[957]),

			.SELF(gen[861]),
			.cell_state(gen[861])
		); 

/******************* CELL 862 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell862 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[766]),
			.N(gen[767]),
			.NE(gen[768]),

			.O(gen[861]),
			.E(gen[863]),

			.SO(gen[956]),
			.S(gen[957]),
			.SE(gen[958]),

			.SELF(gen[862]),
			.cell_state(gen[862])
		); 

/******************* CELL 863 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell863 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[767]),
			.N(gen[768]),
			.NE(gen[769]),

			.O(gen[862]),
			.E(gen[864]),

			.SO(gen[957]),
			.S(gen[958]),
			.SE(gen[959]),

			.SELF(gen[863]),
			.cell_state(gen[863])
		); 

/******************* CELL 864 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell864 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[768]),
			.N(gen[769]),
			.NE(gen[770]),

			.O(gen[863]),
			.E(gen[865]),

			.SO(gen[958]),
			.S(gen[959]),
			.SE(gen[960]),

			.SELF(gen[864]),
			.cell_state(gen[864])
		); 

/******************* CELL 865 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell865 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[769]),
			.N(gen[770]),
			.NE(gen[771]),

			.O(gen[864]),
			.E(gen[866]),

			.SO(gen[959]),
			.S(gen[960]),
			.SE(gen[961]),

			.SELF(gen[865]),
			.cell_state(gen[865])
		); 

/******************* CELL 866 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell866 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[770]),
			.N(gen[771]),
			.NE(gen[772]),

			.O(gen[865]),
			.E(gen[867]),

			.SO(gen[960]),
			.S(gen[961]),
			.SE(gen[962]),

			.SELF(gen[866]),
			.cell_state(gen[866])
		); 

/******************* CELL 867 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell867 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[771]),
			.N(gen[772]),
			.NE(gen[773]),

			.O(gen[866]),
			.E(gen[868]),

			.SO(gen[961]),
			.S(gen[962]),
			.SE(gen[963]),

			.SELF(gen[867]),
			.cell_state(gen[867])
		); 

/******************* CELL 868 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell868 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[772]),
			.N(gen[773]),
			.NE(gen[774]),

			.O(gen[867]),
			.E(gen[869]),

			.SO(gen[962]),
			.S(gen[963]),
			.SE(gen[964]),

			.SELF(gen[868]),
			.cell_state(gen[868])
		); 

/******************* CELL 869 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell869 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[773]),
			.N(gen[774]),
			.NE(gen[775]),

			.O(gen[868]),
			.E(gen[870]),

			.SO(gen[963]),
			.S(gen[964]),
			.SE(gen[965]),

			.SELF(gen[869]),
			.cell_state(gen[869])
		); 

/******************* CELL 870 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell870 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[774]),
			.N(gen[775]),
			.NE(gen[776]),

			.O(gen[869]),
			.E(gen[871]),

			.SO(gen[964]),
			.S(gen[965]),
			.SE(gen[966]),

			.SELF(gen[870]),
			.cell_state(gen[870])
		); 

/******************* CELL 871 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell871 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[775]),
			.N(gen[776]),
			.NE(gen[777]),

			.O(gen[870]),
			.E(gen[872]),

			.SO(gen[965]),
			.S(gen[966]),
			.SE(gen[967]),

			.SELF(gen[871]),
			.cell_state(gen[871])
		); 

/******************* CELL 872 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell872 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[776]),
			.N(gen[777]),
			.NE(gen[778]),

			.O(gen[871]),
			.E(gen[873]),

			.SO(gen[966]),
			.S(gen[967]),
			.SE(gen[968]),

			.SELF(gen[872]),
			.cell_state(gen[872])
		); 

/******************* CELL 873 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell873 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[777]),
			.N(gen[778]),
			.NE(gen[779]),

			.O(gen[872]),
			.E(gen[874]),

			.SO(gen[967]),
			.S(gen[968]),
			.SE(gen[969]),

			.SELF(gen[873]),
			.cell_state(gen[873])
		); 

/******************* CELL 874 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell874 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[778]),
			.N(gen[779]),
			.NE(gen[780]),

			.O(gen[873]),
			.E(gen[875]),

			.SO(gen[968]),
			.S(gen[969]),
			.SE(gen[970]),

			.SELF(gen[874]),
			.cell_state(gen[874])
		); 

/******************* CELL 875 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell875 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[779]),
			.N(gen[780]),
			.NE(gen[781]),

			.O(gen[874]),
			.E(gen[876]),

			.SO(gen[969]),
			.S(gen[970]),
			.SE(gen[971]),

			.SELF(gen[875]),
			.cell_state(gen[875])
		); 

/******************* CELL 876 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell876 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[780]),
			.N(gen[781]),
			.NE(gen[782]),

			.O(gen[875]),
			.E(gen[877]),

			.SO(gen[970]),
			.S(gen[971]),
			.SE(gen[972]),

			.SELF(gen[876]),
			.cell_state(gen[876])
		); 

/******************* CELL 877 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell877 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[781]),
			.N(gen[782]),
			.NE(gen[783]),

			.O(gen[876]),
			.E(gen[878]),

			.SO(gen[971]),
			.S(gen[972]),
			.SE(gen[973]),

			.SELF(gen[877]),
			.cell_state(gen[877])
		); 

/******************* CELL 878 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell878 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[782]),
			.N(gen[783]),
			.NE(gen[784]),

			.O(gen[877]),
			.E(gen[879]),

			.SO(gen[972]),
			.S(gen[973]),
			.SE(gen[974]),

			.SELF(gen[878]),
			.cell_state(gen[878])
		); 

/******************* CELL 879 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell879 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[783]),
			.N(gen[784]),
			.NE(gen[785]),

			.O(gen[878]),
			.E(gen[880]),

			.SO(gen[973]),
			.S(gen[974]),
			.SE(gen[975]),

			.SELF(gen[879]),
			.cell_state(gen[879])
		); 

/******************* CELL 880 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell880 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[784]),
			.N(gen[785]),
			.NE(gen[786]),

			.O(gen[879]),
			.E(gen[881]),

			.SO(gen[974]),
			.S(gen[975]),
			.SE(gen[976]),

			.SELF(gen[880]),
			.cell_state(gen[880])
		); 

/******************* CELL 881 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell881 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[785]),
			.N(gen[786]),
			.NE(gen[787]),

			.O(gen[880]),
			.E(gen[882]),

			.SO(gen[975]),
			.S(gen[976]),
			.SE(gen[977]),

			.SELF(gen[881]),
			.cell_state(gen[881])
		); 

/******************* CELL 882 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell882 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[786]),
			.N(gen[787]),
			.NE(gen[788]),

			.O(gen[881]),
			.E(gen[883]),

			.SO(gen[976]),
			.S(gen[977]),
			.SE(gen[978]),

			.SELF(gen[882]),
			.cell_state(gen[882])
		); 

/******************* CELL 883 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell883 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[787]),
			.N(gen[788]),
			.NE(gen[789]),

			.O(gen[882]),
			.E(gen[884]),

			.SO(gen[977]),
			.S(gen[978]),
			.SE(gen[979]),

			.SELF(gen[883]),
			.cell_state(gen[883])
		); 

/******************* CELL 884 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell884 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[788]),
			.N(gen[789]),
			.NE(gen[790]),

			.O(gen[883]),
			.E(gen[885]),

			.SO(gen[978]),
			.S(gen[979]),
			.SE(gen[980]),

			.SELF(gen[884]),
			.cell_state(gen[884])
		); 

/******************* CELL 885 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell885 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[789]),
			.N(gen[790]),
			.NE(gen[791]),

			.O(gen[884]),
			.E(gen[886]),

			.SO(gen[979]),
			.S(gen[980]),
			.SE(gen[981]),

			.SELF(gen[885]),
			.cell_state(gen[885])
		); 

/******************* CELL 886 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell886 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[790]),
			.N(gen[791]),
			.NE(gen[792]),

			.O(gen[885]),
			.E(gen[887]),

			.SO(gen[980]),
			.S(gen[981]),
			.SE(gen[982]),

			.SELF(gen[886]),
			.cell_state(gen[886])
		); 

/******************* CELL 887 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell887 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[791]),
			.N(gen[792]),
			.NE(gen[793]),

			.O(gen[886]),
			.E(gen[888]),

			.SO(gen[981]),
			.S(gen[982]),
			.SE(gen[983]),

			.SELF(gen[887]),
			.cell_state(gen[887])
		); 

/******************* CELL 888 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell888 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[792]),
			.N(gen[793]),
			.NE(gen[794]),

			.O(gen[887]),
			.E(gen[889]),

			.SO(gen[982]),
			.S(gen[983]),
			.SE(gen[984]),

			.SELF(gen[888]),
			.cell_state(gen[888])
		); 

/******************* CELL 889 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell889 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[793]),
			.N(gen[794]),
			.NE(gen[795]),

			.O(gen[888]),
			.E(gen[890]),

			.SO(gen[983]),
			.S(gen[984]),
			.SE(gen[985]),

			.SELF(gen[889]),
			.cell_state(gen[889])
		); 

/******************* CELL 890 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell890 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[794]),
			.N(gen[795]),
			.NE(gen[796]),

			.O(gen[889]),
			.E(gen[891]),

			.SO(gen[984]),
			.S(gen[985]),
			.SE(gen[986]),

			.SELF(gen[890]),
			.cell_state(gen[890])
		); 

/******************* CELL 891 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell891 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[795]),
			.N(gen[796]),
			.NE(gen[797]),

			.O(gen[890]),
			.E(gen[892]),

			.SO(gen[985]),
			.S(gen[986]),
			.SE(gen[987]),

			.SELF(gen[891]),
			.cell_state(gen[891])
		); 

/******************* CELL 892 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell892 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[796]),
			.N(gen[797]),
			.NE(gen[798]),

			.O(gen[891]),
			.E(gen[893]),

			.SO(gen[986]),
			.S(gen[987]),
			.SE(gen[988]),

			.SELF(gen[892]),
			.cell_state(gen[892])
		); 

/******************* CELL 893 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell893 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[797]),
			.N(gen[798]),
			.NE(gen[799]),

			.O(gen[892]),
			.E(gen[894]),

			.SO(gen[987]),
			.S(gen[988]),
			.SE(gen[989]),

			.SELF(gen[893]),
			.cell_state(gen[893])
		); 

/******************* CELL 894 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell894 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[798]),
			.N(gen[799]),
			.NE(gen[800]),

			.O(gen[893]),
			.E(gen[895]),

			.SO(gen[988]),
			.S(gen[989]),
			.SE(gen[990]),

			.SELF(gen[894]),
			.cell_state(gen[894])
		); 

/******************* CELL 895 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell895 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[799]),
			.N(gen[800]),
			.NE(gen[801]),

			.O(gen[894]),
			.E(gen[896]),

			.SO(gen[989]),
			.S(gen[990]),
			.SE(gen[991]),

			.SELF(gen[895]),
			.cell_state(gen[895])
		); 

/******************* CELL 896 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell896 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[800]),
			.N(gen[801]),
			.NE(gen[802]),

			.O(gen[895]),
			.E(gen[897]),

			.SO(gen[990]),
			.S(gen[991]),
			.SE(gen[992]),

			.SELF(gen[896]),
			.cell_state(gen[896])
		); 

/******************* CELL 897 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell897 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[801]),
			.N(gen[802]),
			.NE(gen[803]),

			.O(gen[896]),
			.E(gen[898]),

			.SO(gen[991]),
			.S(gen[992]),
			.SE(gen[993]),

			.SELF(gen[897]),
			.cell_state(gen[897])
		); 

/******************* CELL 898 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell898 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[802]),
			.N(gen[803]),
			.NE(gen[804]),

			.O(gen[897]),
			.E(gen[899]),

			.SO(gen[992]),
			.S(gen[993]),
			.SE(gen[994]),

			.SELF(gen[898]),
			.cell_state(gen[898])
		); 

/******************* CELL 899 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell899 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[803]),
			.N(gen[804]),
			.NE(gen[805]),

			.O(gen[898]),
			.E(gen[900]),

			.SO(gen[993]),
			.S(gen[994]),
			.SE(gen[995]),

			.SELF(gen[899]),
			.cell_state(gen[899])
		); 

/******************* CELL 900 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell900 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[804]),
			.N(gen[805]),
			.NE(gen[806]),

			.O(gen[899]),
			.E(gen[901]),

			.SO(gen[994]),
			.S(gen[995]),
			.SE(gen[996]),

			.SELF(gen[900]),
			.cell_state(gen[900])
		); 

/******************* CELL 901 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell901 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[805]),
			.N(gen[806]),
			.NE(gen[807]),

			.O(gen[900]),
			.E(gen[902]),

			.SO(gen[995]),
			.S(gen[996]),
			.SE(gen[997]),

			.SELF(gen[901]),
			.cell_state(gen[901])
		); 

/******************* CELL 902 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell902 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[806]),
			.N(gen[807]),
			.NE(gen[808]),

			.O(gen[901]),
			.E(gen[903]),

			.SO(gen[996]),
			.S(gen[997]),
			.SE(gen[998]),

			.SELF(gen[902]),
			.cell_state(gen[902])
		); 

/******************* CELL 903 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell903 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[807]),
			.N(gen[808]),
			.NE(gen[809]),

			.O(gen[902]),
			.E(gen[904]),

			.SO(gen[997]),
			.S(gen[998]),
			.SE(gen[999]),

			.SELF(gen[903]),
			.cell_state(gen[903])
		); 

/******************* CELL 904 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell904 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[808]),
			.N(gen[809]),
			.NE(gen[810]),

			.O(gen[903]),
			.E(gen[905]),

			.SO(gen[998]),
			.S(gen[999]),
			.SE(gen[1000]),

			.SELF(gen[904]),
			.cell_state(gen[904])
		); 

/******************* CELL 905 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell905 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[809]),
			.N(gen[810]),
			.NE(gen[811]),

			.O(gen[904]),
			.E(gen[906]),

			.SO(gen[999]),
			.S(gen[1000]),
			.SE(gen[1001]),

			.SELF(gen[905]),
			.cell_state(gen[905])
		); 

/******************* CELL 906 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell906 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[810]),
			.N(gen[811]),
			.NE(gen[812]),

			.O(gen[905]),
			.E(gen[907]),

			.SO(gen[1000]),
			.S(gen[1001]),
			.SE(gen[1002]),

			.SELF(gen[906]),
			.cell_state(gen[906])
		); 

/******************* CELL 907 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell907 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[811]),
			.N(gen[812]),
			.NE(gen[813]),

			.O(gen[906]),
			.E(gen[908]),

			.SO(gen[1001]),
			.S(gen[1002]),
			.SE(gen[1003]),

			.SELF(gen[907]),
			.cell_state(gen[907])
		); 

/******************* CELL 908 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell908 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[812]),
			.N(gen[813]),
			.NE(gen[814]),

			.O(gen[907]),
			.E(gen[909]),

			.SO(gen[1002]),
			.S(gen[1003]),
			.SE(gen[1004]),

			.SELF(gen[908]),
			.cell_state(gen[908])
		); 

/******************* CELL 909 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell909 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[813]),
			.N(gen[814]),
			.NE(gen[815]),

			.O(gen[908]),
			.E(gen[910]),

			.SO(gen[1003]),
			.S(gen[1004]),
			.SE(gen[1005]),

			.SELF(gen[909]),
			.cell_state(gen[909])
		); 

/******************* CELL 910 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell910 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[814]),
			.N(gen[815]),
			.NE(gen[816]),

			.O(gen[909]),
			.E(gen[911]),

			.SO(gen[1004]),
			.S(gen[1005]),
			.SE(gen[1006]),

			.SELF(gen[910]),
			.cell_state(gen[910])
		); 

/******************* CELL 911 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell911 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[815]),
			.N(gen[816]),
			.NE(gen[817]),

			.O(gen[910]),
			.E(gen[912]),

			.SO(gen[1005]),
			.S(gen[1006]),
			.SE(gen[1007]),

			.SELF(gen[911]),
			.cell_state(gen[911])
		); 

/******************* CELL 912 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell912 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[816]),
			.N(gen[817]),
			.NE(gen[818]),

			.O(gen[911]),
			.E(gen[913]),

			.SO(gen[1006]),
			.S(gen[1007]),
			.SE(gen[1008]),

			.SELF(gen[912]),
			.cell_state(gen[912])
		); 

/******************* CELL 913 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell913 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[817]),
			.N(gen[818]),
			.NE(gen[819]),

			.O(gen[912]),
			.E(gen[914]),

			.SO(gen[1007]),
			.S(gen[1008]),
			.SE(gen[1009]),

			.SELF(gen[913]),
			.cell_state(gen[913])
		); 

/******************* CELL 914 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell914 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[818]),
			.N(gen[819]),
			.NE(gen[820]),

			.O(gen[913]),
			.E(gen[915]),

			.SO(gen[1008]),
			.S(gen[1009]),
			.SE(gen[1010]),

			.SELF(gen[914]),
			.cell_state(gen[914])
		); 

/******************* CELL 915 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell915 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[819]),
			.N(gen[820]),
			.NE(gen[821]),

			.O(gen[914]),
			.E(gen[916]),

			.SO(gen[1009]),
			.S(gen[1010]),
			.SE(gen[1011]),

			.SELF(gen[915]),
			.cell_state(gen[915])
		); 

/******************* CELL 916 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell916 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[820]),
			.N(gen[821]),
			.NE(gen[822]),

			.O(gen[915]),
			.E(gen[917]),

			.SO(gen[1010]),
			.S(gen[1011]),
			.SE(gen[1012]),

			.SELF(gen[916]),
			.cell_state(gen[916])
		); 

/******************* CELL 917 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell917 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[821]),
			.N(gen[822]),
			.NE(gen[823]),

			.O(gen[916]),
			.E(gen[918]),

			.SO(gen[1011]),
			.S(gen[1012]),
			.SE(gen[1013]),

			.SELF(gen[917]),
			.cell_state(gen[917])
		); 

/******************* CELL 918 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell918 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[822]),
			.N(gen[823]),
			.NE(gen[824]),

			.O(gen[917]),
			.E(gen[919]),

			.SO(gen[1012]),
			.S(gen[1013]),
			.SE(gen[1014]),

			.SELF(gen[918]),
			.cell_state(gen[918])
		); 

/******************* CELL 919 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell919 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[823]),
			.N(gen[824]),
			.NE(gen[825]),

			.O(gen[918]),
			.E(gen[920]),

			.SO(gen[1013]),
			.S(gen[1014]),
			.SE(gen[1015]),

			.SELF(gen[919]),
			.cell_state(gen[919])
		); 

/******************* CELL 920 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell920 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[824]),
			.N(gen[825]),
			.NE(gen[826]),

			.O(gen[919]),
			.E(gen[921]),

			.SO(gen[1014]),
			.S(gen[1015]),
			.SE(gen[1016]),

			.SELF(gen[920]),
			.cell_state(gen[920])
		); 

/******************* CELL 921 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell921 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[825]),
			.N(gen[826]),
			.NE(gen[827]),

			.O(gen[920]),
			.E(gen[922]),

			.SO(gen[1015]),
			.S(gen[1016]),
			.SE(gen[1017]),

			.SELF(gen[921]),
			.cell_state(gen[921])
		); 

/******************* CELL 922 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell922 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[826]),
			.N(gen[827]),
			.NE(gen[828]),

			.O(gen[921]),
			.E(gen[923]),

			.SO(gen[1016]),
			.S(gen[1017]),
			.SE(gen[1018]),

			.SELF(gen[922]),
			.cell_state(gen[922])
		); 

/******************* CELL 923 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell923 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[827]),
			.N(gen[828]),
			.NE(gen[829]),

			.O(gen[922]),
			.E(gen[924]),

			.SO(gen[1017]),
			.S(gen[1018]),
			.SE(gen[1019]),

			.SELF(gen[923]),
			.cell_state(gen[923])
		); 

/******************* CELL 924 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell924 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[828]),
			.N(gen[829]),
			.NE(gen[830]),

			.O(gen[923]),
			.E(gen[925]),

			.SO(gen[1018]),
			.S(gen[1019]),
			.SE(gen[1020]),

			.SELF(gen[924]),
			.cell_state(gen[924])
		); 

/******************* CELL 925 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell925 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[829]),
			.N(gen[830]),
			.NE(gen[831]),

			.O(gen[924]),
			.E(gen[926]),

			.SO(gen[1019]),
			.S(gen[1020]),
			.SE(gen[1021]),

			.SELF(gen[925]),
			.cell_state(gen[925])
		); 

/******************* CELL 926 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell926 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[830]),
			.N(gen[831]),
			.NE(gen[832]),

			.O(gen[925]),
			.E(gen[927]),

			.SO(gen[1020]),
			.S(gen[1021]),
			.SE(gen[1022]),

			.SELF(gen[926]),
			.cell_state(gen[926])
		); 

/******************* CELL 927 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell927 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[831]),
			.N(gen[832]),
			.NE(gen[833]),

			.O(gen[926]),
			.E(gen[928]),

			.SO(gen[1021]),
			.S(gen[1022]),
			.SE(gen[1023]),

			.SELF(gen[927]),
			.cell_state(gen[927])
		); 

/******************* CELL 928 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell928 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[832]),
			.N(gen[833]),
			.NE(gen[834]),

			.O(gen[927]),
			.E(gen[929]),

			.SO(gen[1022]),
			.S(gen[1023]),
			.SE(gen[1024]),

			.SELF(gen[928]),
			.cell_state(gen[928])
		); 

/******************* CELL 929 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell929 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[833]),
			.N(gen[834]),
			.NE(gen[835]),

			.O(gen[928]),
			.E(gen[930]),

			.SO(gen[1023]),
			.S(gen[1024]),
			.SE(gen[1025]),

			.SELF(gen[929]),
			.cell_state(gen[929])
		); 

/******************* CELL 930 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell930 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[834]),
			.N(gen[835]),
			.NE(gen[836]),

			.O(gen[929]),
			.E(gen[931]),

			.SO(gen[1024]),
			.S(gen[1025]),
			.SE(gen[1026]),

			.SELF(gen[930]),
			.cell_state(gen[930])
		); 

/******************* CELL 931 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell931 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[835]),
			.N(gen[836]),
			.NE(gen[837]),

			.O(gen[930]),
			.E(gen[932]),

			.SO(gen[1025]),
			.S(gen[1026]),
			.SE(gen[1027]),

			.SELF(gen[931]),
			.cell_state(gen[931])
		); 

/******************* CELL 932 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell932 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[836]),
			.N(gen[837]),
			.NE(gen[838]),

			.O(gen[931]),
			.E(gen[933]),

			.SO(gen[1026]),
			.S(gen[1027]),
			.SE(gen[1028]),

			.SELF(gen[932]),
			.cell_state(gen[932])
		); 

/******************* CELL 933 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell933 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[837]),
			.N(gen[838]),
			.NE(gen[839]),

			.O(gen[932]),
			.E(gen[934]),

			.SO(gen[1027]),
			.S(gen[1028]),
			.SE(gen[1029]),

			.SELF(gen[933]),
			.cell_state(gen[933])
		); 

/******************* CELL 934 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell934 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[838]),
			.N(gen[839]),
			.NE(gen[840]),

			.O(gen[933]),
			.E(gen[935]),

			.SO(gen[1028]),
			.S(gen[1029]),
			.SE(gen[1030]),

			.SELF(gen[934]),
			.cell_state(gen[934])
		); 

/******************* CELL 935 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell935 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[839]),
			.N(gen[840]),
			.NE(gen[841]),

			.O(gen[934]),
			.E(gen[936]),

			.SO(gen[1029]),
			.S(gen[1030]),
			.SE(gen[1031]),

			.SELF(gen[935]),
			.cell_state(gen[935])
		); 

/******************* CELL 936 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell936 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[840]),
			.N(gen[841]),
			.NE(gen[842]),

			.O(gen[935]),
			.E(gen[937]),

			.SO(gen[1030]),
			.S(gen[1031]),
			.SE(gen[1032]),

			.SELF(gen[936]),
			.cell_state(gen[936])
		); 

/******************* CELL 937 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell937 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[841]),
			.N(gen[842]),
			.NE(gen[843]),

			.O(gen[936]),
			.E(gen[938]),

			.SO(gen[1031]),
			.S(gen[1032]),
			.SE(gen[1033]),

			.SELF(gen[937]),
			.cell_state(gen[937])
		); 

/******************* CELL 938 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell938 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[842]),
			.N(gen[843]),
			.NE(gen[844]),

			.O(gen[937]),
			.E(gen[939]),

			.SO(gen[1032]),
			.S(gen[1033]),
			.SE(gen[1034]),

			.SELF(gen[938]),
			.cell_state(gen[938])
		); 

/******************* CELL 939 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell939 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[843]),
			.N(gen[844]),
			.NE(gen[845]),

			.O(gen[938]),
			.E(gen[940]),

			.SO(gen[1033]),
			.S(gen[1034]),
			.SE(gen[1035]),

			.SELF(gen[939]),
			.cell_state(gen[939])
		); 

/******************* CELL 940 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell940 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[844]),
			.N(gen[845]),
			.NE(gen[846]),

			.O(gen[939]),
			.E(gen[941]),

			.SO(gen[1034]),
			.S(gen[1035]),
			.SE(gen[1036]),

			.SELF(gen[940]),
			.cell_state(gen[940])
		); 

/******************* CELL 941 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell941 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[845]),
			.N(gen[846]),
			.NE(gen[847]),

			.O(gen[940]),
			.E(gen[942]),

			.SO(gen[1035]),
			.S(gen[1036]),
			.SE(gen[1037]),

			.SELF(gen[941]),
			.cell_state(gen[941])
		); 

/******************* CELL 942 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell942 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[846]),
			.N(gen[847]),
			.NE(gen[848]),

			.O(gen[941]),
			.E(gen[943]),

			.SO(gen[1036]),
			.S(gen[1037]),
			.SE(gen[1038]),

			.SELF(gen[942]),
			.cell_state(gen[942])
		); 

/******************* CELL 943 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell943 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[847]),
			.N(gen[848]),
			.NE(gen[849]),

			.O(gen[942]),
			.E(gen[944]),

			.SO(gen[1037]),
			.S(gen[1038]),
			.SE(gen[1039]),

			.SELF(gen[943]),
			.cell_state(gen[943])
		); 

/******************* CELL 944 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell944 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[848]),
			.N(gen[849]),
			.NE(gen[850]),

			.O(gen[943]),
			.E(gen[945]),

			.SO(gen[1038]),
			.S(gen[1039]),
			.SE(gen[1040]),

			.SELF(gen[944]),
			.cell_state(gen[944])
		); 

/******************* CELL 945 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell945 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[849]),
			.N(gen[850]),
			.NE(gen[851]),

			.O(gen[944]),
			.E(gen[946]),

			.SO(gen[1039]),
			.S(gen[1040]),
			.SE(gen[1041]),

			.SELF(gen[945]),
			.cell_state(gen[945])
		); 

/******************* CELL 946 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell946 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[850]),
			.N(gen[851]),
			.NE(gen[852]),

			.O(gen[945]),
			.E(gen[947]),

			.SO(gen[1040]),
			.S(gen[1041]),
			.SE(gen[1042]),

			.SELF(gen[946]),
			.cell_state(gen[946])
		); 

/******************* CELL 947 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell947 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[851]),
			.N(gen[852]),
			.NE(gen[853]),

			.O(gen[946]),
			.E(gen[948]),

			.SO(gen[1041]),
			.S(gen[1042]),
			.SE(gen[1043]),

			.SELF(gen[947]),
			.cell_state(gen[947])
		); 

/******************* CELL 948 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell948 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[852]),
			.N(gen[853]),
			.NE(gen[854]),

			.O(gen[947]),
			.E(gen[949]),

			.SO(gen[1042]),
			.S(gen[1043]),
			.SE(gen[1044]),

			.SELF(gen[948]),
			.cell_state(gen[948])
		); 

/******************* CELL 949 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell949 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[853]),
			.N(gen[854]),
			.NE(gen[853]),

			.O(gen[948]),
			.E(gen[948]),

			.SO(gen[1043]),
			.S(gen[1044]),
			.SE(gen[1043]),

			.SELF(gen[949]),
			.cell_state(gen[949])
		); 

/******************* CELL 950 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell950 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[856]),
			.N(gen[855]),
			.NE(gen[856]),

			.O(gen[951]),
			.E(gen[951]),

			.SO(gen[1046]),
			.S(gen[1045]),
			.SE(gen[1046]),

			.SELF(gen[950]),
			.cell_state(gen[950])
		); 

/******************* CELL 951 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell951 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[855]),
			.N(gen[856]),
			.NE(gen[857]),

			.O(gen[950]),
			.E(gen[952]),

			.SO(gen[1045]),
			.S(gen[1046]),
			.SE(gen[1047]),

			.SELF(gen[951]),
			.cell_state(gen[951])
		); 

/******************* CELL 952 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell952 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[856]),
			.N(gen[857]),
			.NE(gen[858]),

			.O(gen[951]),
			.E(gen[953]),

			.SO(gen[1046]),
			.S(gen[1047]),
			.SE(gen[1048]),

			.SELF(gen[952]),
			.cell_state(gen[952])
		); 

/******************* CELL 953 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell953 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[857]),
			.N(gen[858]),
			.NE(gen[859]),

			.O(gen[952]),
			.E(gen[954]),

			.SO(gen[1047]),
			.S(gen[1048]),
			.SE(gen[1049]),

			.SELF(gen[953]),
			.cell_state(gen[953])
		); 

/******************* CELL 954 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell954 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[858]),
			.N(gen[859]),
			.NE(gen[860]),

			.O(gen[953]),
			.E(gen[955]),

			.SO(gen[1048]),
			.S(gen[1049]),
			.SE(gen[1050]),

			.SELF(gen[954]),
			.cell_state(gen[954])
		); 

/******************* CELL 955 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell955 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[859]),
			.N(gen[860]),
			.NE(gen[861]),

			.O(gen[954]),
			.E(gen[956]),

			.SO(gen[1049]),
			.S(gen[1050]),
			.SE(gen[1051]),

			.SELF(gen[955]),
			.cell_state(gen[955])
		); 

/******************* CELL 956 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell956 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[860]),
			.N(gen[861]),
			.NE(gen[862]),

			.O(gen[955]),
			.E(gen[957]),

			.SO(gen[1050]),
			.S(gen[1051]),
			.SE(gen[1052]),

			.SELF(gen[956]),
			.cell_state(gen[956])
		); 

/******************* CELL 957 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell957 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[861]),
			.N(gen[862]),
			.NE(gen[863]),

			.O(gen[956]),
			.E(gen[958]),

			.SO(gen[1051]),
			.S(gen[1052]),
			.SE(gen[1053]),

			.SELF(gen[957]),
			.cell_state(gen[957])
		); 

/******************* CELL 958 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell958 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[862]),
			.N(gen[863]),
			.NE(gen[864]),

			.O(gen[957]),
			.E(gen[959]),

			.SO(gen[1052]),
			.S(gen[1053]),
			.SE(gen[1054]),

			.SELF(gen[958]),
			.cell_state(gen[958])
		); 

/******************* CELL 959 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell959 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[863]),
			.N(gen[864]),
			.NE(gen[865]),

			.O(gen[958]),
			.E(gen[960]),

			.SO(gen[1053]),
			.S(gen[1054]),
			.SE(gen[1055]),

			.SELF(gen[959]),
			.cell_state(gen[959])
		); 

/******************* CELL 960 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell960 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[864]),
			.N(gen[865]),
			.NE(gen[866]),

			.O(gen[959]),
			.E(gen[961]),

			.SO(gen[1054]),
			.S(gen[1055]),
			.SE(gen[1056]),

			.SELF(gen[960]),
			.cell_state(gen[960])
		); 

/******************* CELL 961 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell961 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[865]),
			.N(gen[866]),
			.NE(gen[867]),

			.O(gen[960]),
			.E(gen[962]),

			.SO(gen[1055]),
			.S(gen[1056]),
			.SE(gen[1057]),

			.SELF(gen[961]),
			.cell_state(gen[961])
		); 

/******************* CELL 962 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell962 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[866]),
			.N(gen[867]),
			.NE(gen[868]),

			.O(gen[961]),
			.E(gen[963]),

			.SO(gen[1056]),
			.S(gen[1057]),
			.SE(gen[1058]),

			.SELF(gen[962]),
			.cell_state(gen[962])
		); 

/******************* CELL 963 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell963 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[867]),
			.N(gen[868]),
			.NE(gen[869]),

			.O(gen[962]),
			.E(gen[964]),

			.SO(gen[1057]),
			.S(gen[1058]),
			.SE(gen[1059]),

			.SELF(gen[963]),
			.cell_state(gen[963])
		); 

/******************* CELL 964 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell964 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[868]),
			.N(gen[869]),
			.NE(gen[870]),

			.O(gen[963]),
			.E(gen[965]),

			.SO(gen[1058]),
			.S(gen[1059]),
			.SE(gen[1060]),

			.SELF(gen[964]),
			.cell_state(gen[964])
		); 

/******************* CELL 965 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell965 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[869]),
			.N(gen[870]),
			.NE(gen[871]),

			.O(gen[964]),
			.E(gen[966]),

			.SO(gen[1059]),
			.S(gen[1060]),
			.SE(gen[1061]),

			.SELF(gen[965]),
			.cell_state(gen[965])
		); 

/******************* CELL 966 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell966 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[870]),
			.N(gen[871]),
			.NE(gen[872]),

			.O(gen[965]),
			.E(gen[967]),

			.SO(gen[1060]),
			.S(gen[1061]),
			.SE(gen[1062]),

			.SELF(gen[966]),
			.cell_state(gen[966])
		); 

/******************* CELL 967 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell967 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[871]),
			.N(gen[872]),
			.NE(gen[873]),

			.O(gen[966]),
			.E(gen[968]),

			.SO(gen[1061]),
			.S(gen[1062]),
			.SE(gen[1063]),

			.SELF(gen[967]),
			.cell_state(gen[967])
		); 

/******************* CELL 968 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell968 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[872]),
			.N(gen[873]),
			.NE(gen[874]),

			.O(gen[967]),
			.E(gen[969]),

			.SO(gen[1062]),
			.S(gen[1063]),
			.SE(gen[1064]),

			.SELF(gen[968]),
			.cell_state(gen[968])
		); 

/******************* CELL 969 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell969 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[873]),
			.N(gen[874]),
			.NE(gen[875]),

			.O(gen[968]),
			.E(gen[970]),

			.SO(gen[1063]),
			.S(gen[1064]),
			.SE(gen[1065]),

			.SELF(gen[969]),
			.cell_state(gen[969])
		); 

/******************* CELL 970 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell970 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[874]),
			.N(gen[875]),
			.NE(gen[876]),

			.O(gen[969]),
			.E(gen[971]),

			.SO(gen[1064]),
			.S(gen[1065]),
			.SE(gen[1066]),

			.SELF(gen[970]),
			.cell_state(gen[970])
		); 

/******************* CELL 971 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell971 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[875]),
			.N(gen[876]),
			.NE(gen[877]),

			.O(gen[970]),
			.E(gen[972]),

			.SO(gen[1065]),
			.S(gen[1066]),
			.SE(gen[1067]),

			.SELF(gen[971]),
			.cell_state(gen[971])
		); 

/******************* CELL 972 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell972 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[876]),
			.N(gen[877]),
			.NE(gen[878]),

			.O(gen[971]),
			.E(gen[973]),

			.SO(gen[1066]),
			.S(gen[1067]),
			.SE(gen[1068]),

			.SELF(gen[972]),
			.cell_state(gen[972])
		); 

/******************* CELL 973 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell973 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[877]),
			.N(gen[878]),
			.NE(gen[879]),

			.O(gen[972]),
			.E(gen[974]),

			.SO(gen[1067]),
			.S(gen[1068]),
			.SE(gen[1069]),

			.SELF(gen[973]),
			.cell_state(gen[973])
		); 

/******************* CELL 974 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell974 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[878]),
			.N(gen[879]),
			.NE(gen[880]),

			.O(gen[973]),
			.E(gen[975]),

			.SO(gen[1068]),
			.S(gen[1069]),
			.SE(gen[1070]),

			.SELF(gen[974]),
			.cell_state(gen[974])
		); 

/******************* CELL 975 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell975 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[879]),
			.N(gen[880]),
			.NE(gen[881]),

			.O(gen[974]),
			.E(gen[976]),

			.SO(gen[1069]),
			.S(gen[1070]),
			.SE(gen[1071]),

			.SELF(gen[975]),
			.cell_state(gen[975])
		); 

/******************* CELL 976 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell976 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[880]),
			.N(gen[881]),
			.NE(gen[882]),

			.O(gen[975]),
			.E(gen[977]),

			.SO(gen[1070]),
			.S(gen[1071]),
			.SE(gen[1072]),

			.SELF(gen[976]),
			.cell_state(gen[976])
		); 

/******************* CELL 977 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell977 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[881]),
			.N(gen[882]),
			.NE(gen[883]),

			.O(gen[976]),
			.E(gen[978]),

			.SO(gen[1071]),
			.S(gen[1072]),
			.SE(gen[1073]),

			.SELF(gen[977]),
			.cell_state(gen[977])
		); 

/******************* CELL 978 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell978 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[882]),
			.N(gen[883]),
			.NE(gen[884]),

			.O(gen[977]),
			.E(gen[979]),

			.SO(gen[1072]),
			.S(gen[1073]),
			.SE(gen[1074]),

			.SELF(gen[978]),
			.cell_state(gen[978])
		); 

/******************* CELL 979 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell979 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[883]),
			.N(gen[884]),
			.NE(gen[885]),

			.O(gen[978]),
			.E(gen[980]),

			.SO(gen[1073]),
			.S(gen[1074]),
			.SE(gen[1075]),

			.SELF(gen[979]),
			.cell_state(gen[979])
		); 

/******************* CELL 980 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell980 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[884]),
			.N(gen[885]),
			.NE(gen[886]),

			.O(gen[979]),
			.E(gen[981]),

			.SO(gen[1074]),
			.S(gen[1075]),
			.SE(gen[1076]),

			.SELF(gen[980]),
			.cell_state(gen[980])
		); 

/******************* CELL 981 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell981 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[885]),
			.N(gen[886]),
			.NE(gen[887]),

			.O(gen[980]),
			.E(gen[982]),

			.SO(gen[1075]),
			.S(gen[1076]),
			.SE(gen[1077]),

			.SELF(gen[981]),
			.cell_state(gen[981])
		); 

/******************* CELL 982 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell982 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[886]),
			.N(gen[887]),
			.NE(gen[888]),

			.O(gen[981]),
			.E(gen[983]),

			.SO(gen[1076]),
			.S(gen[1077]),
			.SE(gen[1078]),

			.SELF(gen[982]),
			.cell_state(gen[982])
		); 

/******************* CELL 983 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell983 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[887]),
			.N(gen[888]),
			.NE(gen[889]),

			.O(gen[982]),
			.E(gen[984]),

			.SO(gen[1077]),
			.S(gen[1078]),
			.SE(gen[1079]),

			.SELF(gen[983]),
			.cell_state(gen[983])
		); 

/******************* CELL 984 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell984 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[888]),
			.N(gen[889]),
			.NE(gen[890]),

			.O(gen[983]),
			.E(gen[985]),

			.SO(gen[1078]),
			.S(gen[1079]),
			.SE(gen[1080]),

			.SELF(gen[984]),
			.cell_state(gen[984])
		); 

/******************* CELL 985 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell985 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[889]),
			.N(gen[890]),
			.NE(gen[891]),

			.O(gen[984]),
			.E(gen[986]),

			.SO(gen[1079]),
			.S(gen[1080]),
			.SE(gen[1081]),

			.SELF(gen[985]),
			.cell_state(gen[985])
		); 

/******************* CELL 986 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell986 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[890]),
			.N(gen[891]),
			.NE(gen[892]),

			.O(gen[985]),
			.E(gen[987]),

			.SO(gen[1080]),
			.S(gen[1081]),
			.SE(gen[1082]),

			.SELF(gen[986]),
			.cell_state(gen[986])
		); 

/******************* CELL 987 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell987 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[891]),
			.N(gen[892]),
			.NE(gen[893]),

			.O(gen[986]),
			.E(gen[988]),

			.SO(gen[1081]),
			.S(gen[1082]),
			.SE(gen[1083]),

			.SELF(gen[987]),
			.cell_state(gen[987])
		); 

/******************* CELL 988 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell988 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[892]),
			.N(gen[893]),
			.NE(gen[894]),

			.O(gen[987]),
			.E(gen[989]),

			.SO(gen[1082]),
			.S(gen[1083]),
			.SE(gen[1084]),

			.SELF(gen[988]),
			.cell_state(gen[988])
		); 

/******************* CELL 989 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell989 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[893]),
			.N(gen[894]),
			.NE(gen[895]),

			.O(gen[988]),
			.E(gen[990]),

			.SO(gen[1083]),
			.S(gen[1084]),
			.SE(gen[1085]),

			.SELF(gen[989]),
			.cell_state(gen[989])
		); 

/******************* CELL 990 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell990 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[894]),
			.N(gen[895]),
			.NE(gen[896]),

			.O(gen[989]),
			.E(gen[991]),

			.SO(gen[1084]),
			.S(gen[1085]),
			.SE(gen[1086]),

			.SELF(gen[990]),
			.cell_state(gen[990])
		); 

/******************* CELL 991 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell991 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[895]),
			.N(gen[896]),
			.NE(gen[897]),

			.O(gen[990]),
			.E(gen[992]),

			.SO(gen[1085]),
			.S(gen[1086]),
			.SE(gen[1087]),

			.SELF(gen[991]),
			.cell_state(gen[991])
		); 

/******************* CELL 992 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell992 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[896]),
			.N(gen[897]),
			.NE(gen[898]),

			.O(gen[991]),
			.E(gen[993]),

			.SO(gen[1086]),
			.S(gen[1087]),
			.SE(gen[1088]),

			.SELF(gen[992]),
			.cell_state(gen[992])
		); 

/******************* CELL 993 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell993 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[897]),
			.N(gen[898]),
			.NE(gen[899]),

			.O(gen[992]),
			.E(gen[994]),

			.SO(gen[1087]),
			.S(gen[1088]),
			.SE(gen[1089]),

			.SELF(gen[993]),
			.cell_state(gen[993])
		); 

/******************* CELL 994 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell994 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[898]),
			.N(gen[899]),
			.NE(gen[900]),

			.O(gen[993]),
			.E(gen[995]),

			.SO(gen[1088]),
			.S(gen[1089]),
			.SE(gen[1090]),

			.SELF(gen[994]),
			.cell_state(gen[994])
		); 

/******************* CELL 995 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell995 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[899]),
			.N(gen[900]),
			.NE(gen[901]),

			.O(gen[994]),
			.E(gen[996]),

			.SO(gen[1089]),
			.S(gen[1090]),
			.SE(gen[1091]),

			.SELF(gen[995]),
			.cell_state(gen[995])
		); 

/******************* CELL 996 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell996 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[900]),
			.N(gen[901]),
			.NE(gen[902]),

			.O(gen[995]),
			.E(gen[997]),

			.SO(gen[1090]),
			.S(gen[1091]),
			.SE(gen[1092]),

			.SELF(gen[996]),
			.cell_state(gen[996])
		); 

/******************* CELL 997 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell997 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[901]),
			.N(gen[902]),
			.NE(gen[903]),

			.O(gen[996]),
			.E(gen[998]),

			.SO(gen[1091]),
			.S(gen[1092]),
			.SE(gen[1093]),

			.SELF(gen[997]),
			.cell_state(gen[997])
		); 

/******************* CELL 998 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell998 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[902]),
			.N(gen[903]),
			.NE(gen[904]),

			.O(gen[997]),
			.E(gen[999]),

			.SO(gen[1092]),
			.S(gen[1093]),
			.SE(gen[1094]),

			.SELF(gen[998]),
			.cell_state(gen[998])
		); 

/******************* CELL 999 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell999 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[903]),
			.N(gen[904]),
			.NE(gen[905]),

			.O(gen[998]),
			.E(gen[1000]),

			.SO(gen[1093]),
			.S(gen[1094]),
			.SE(gen[1095]),

			.SELF(gen[999]),
			.cell_state(gen[999])
		); 

/******************* CELL 1000 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1000 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[904]),
			.N(gen[905]),
			.NE(gen[906]),

			.O(gen[999]),
			.E(gen[1001]),

			.SO(gen[1094]),
			.S(gen[1095]),
			.SE(gen[1096]),

			.SELF(gen[1000]),
			.cell_state(gen[1000])
		); 

/******************* CELL 1001 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1001 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[905]),
			.N(gen[906]),
			.NE(gen[907]),

			.O(gen[1000]),
			.E(gen[1002]),

			.SO(gen[1095]),
			.S(gen[1096]),
			.SE(gen[1097]),

			.SELF(gen[1001]),
			.cell_state(gen[1001])
		); 

/******************* CELL 1002 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1002 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[906]),
			.N(gen[907]),
			.NE(gen[908]),

			.O(gen[1001]),
			.E(gen[1003]),

			.SO(gen[1096]),
			.S(gen[1097]),
			.SE(gen[1098]),

			.SELF(gen[1002]),
			.cell_state(gen[1002])
		); 

/******************* CELL 1003 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1003 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[907]),
			.N(gen[908]),
			.NE(gen[909]),

			.O(gen[1002]),
			.E(gen[1004]),

			.SO(gen[1097]),
			.S(gen[1098]),
			.SE(gen[1099]),

			.SELF(gen[1003]),
			.cell_state(gen[1003])
		); 

/******************* CELL 1004 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1004 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[908]),
			.N(gen[909]),
			.NE(gen[910]),

			.O(gen[1003]),
			.E(gen[1005]),

			.SO(gen[1098]),
			.S(gen[1099]),
			.SE(gen[1100]),

			.SELF(gen[1004]),
			.cell_state(gen[1004])
		); 

/******************* CELL 1005 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1005 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[909]),
			.N(gen[910]),
			.NE(gen[911]),

			.O(gen[1004]),
			.E(gen[1006]),

			.SO(gen[1099]),
			.S(gen[1100]),
			.SE(gen[1101]),

			.SELF(gen[1005]),
			.cell_state(gen[1005])
		); 

/******************* CELL 1006 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1006 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[910]),
			.N(gen[911]),
			.NE(gen[912]),

			.O(gen[1005]),
			.E(gen[1007]),

			.SO(gen[1100]),
			.S(gen[1101]),
			.SE(gen[1102]),

			.SELF(gen[1006]),
			.cell_state(gen[1006])
		); 

/******************* CELL 1007 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1007 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[911]),
			.N(gen[912]),
			.NE(gen[913]),

			.O(gen[1006]),
			.E(gen[1008]),

			.SO(gen[1101]),
			.S(gen[1102]),
			.SE(gen[1103]),

			.SELF(gen[1007]),
			.cell_state(gen[1007])
		); 

/******************* CELL 1008 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1008 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[912]),
			.N(gen[913]),
			.NE(gen[914]),

			.O(gen[1007]),
			.E(gen[1009]),

			.SO(gen[1102]),
			.S(gen[1103]),
			.SE(gen[1104]),

			.SELF(gen[1008]),
			.cell_state(gen[1008])
		); 

/******************* CELL 1009 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1009 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[913]),
			.N(gen[914]),
			.NE(gen[915]),

			.O(gen[1008]),
			.E(gen[1010]),

			.SO(gen[1103]),
			.S(gen[1104]),
			.SE(gen[1105]),

			.SELF(gen[1009]),
			.cell_state(gen[1009])
		); 

/******************* CELL 1010 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1010 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[914]),
			.N(gen[915]),
			.NE(gen[916]),

			.O(gen[1009]),
			.E(gen[1011]),

			.SO(gen[1104]),
			.S(gen[1105]),
			.SE(gen[1106]),

			.SELF(gen[1010]),
			.cell_state(gen[1010])
		); 

/******************* CELL 1011 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1011 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[915]),
			.N(gen[916]),
			.NE(gen[917]),

			.O(gen[1010]),
			.E(gen[1012]),

			.SO(gen[1105]),
			.S(gen[1106]),
			.SE(gen[1107]),

			.SELF(gen[1011]),
			.cell_state(gen[1011])
		); 

/******************* CELL 1012 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1012 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[916]),
			.N(gen[917]),
			.NE(gen[918]),

			.O(gen[1011]),
			.E(gen[1013]),

			.SO(gen[1106]),
			.S(gen[1107]),
			.SE(gen[1108]),

			.SELF(gen[1012]),
			.cell_state(gen[1012])
		); 

/******************* CELL 1013 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1013 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[917]),
			.N(gen[918]),
			.NE(gen[919]),

			.O(gen[1012]),
			.E(gen[1014]),

			.SO(gen[1107]),
			.S(gen[1108]),
			.SE(gen[1109]),

			.SELF(gen[1013]),
			.cell_state(gen[1013])
		); 

/******************* CELL 1014 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1014 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[918]),
			.N(gen[919]),
			.NE(gen[920]),

			.O(gen[1013]),
			.E(gen[1015]),

			.SO(gen[1108]),
			.S(gen[1109]),
			.SE(gen[1110]),

			.SELF(gen[1014]),
			.cell_state(gen[1014])
		); 

/******************* CELL 1015 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1015 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[919]),
			.N(gen[920]),
			.NE(gen[921]),

			.O(gen[1014]),
			.E(gen[1016]),

			.SO(gen[1109]),
			.S(gen[1110]),
			.SE(gen[1111]),

			.SELF(gen[1015]),
			.cell_state(gen[1015])
		); 

/******************* CELL 1016 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1016 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[920]),
			.N(gen[921]),
			.NE(gen[922]),

			.O(gen[1015]),
			.E(gen[1017]),

			.SO(gen[1110]),
			.S(gen[1111]),
			.SE(gen[1112]),

			.SELF(gen[1016]),
			.cell_state(gen[1016])
		); 

/******************* CELL 1017 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1017 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[921]),
			.N(gen[922]),
			.NE(gen[923]),

			.O(gen[1016]),
			.E(gen[1018]),

			.SO(gen[1111]),
			.S(gen[1112]),
			.SE(gen[1113]),

			.SELF(gen[1017]),
			.cell_state(gen[1017])
		); 

/******************* CELL 1018 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1018 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[922]),
			.N(gen[923]),
			.NE(gen[924]),

			.O(gen[1017]),
			.E(gen[1019]),

			.SO(gen[1112]),
			.S(gen[1113]),
			.SE(gen[1114]),

			.SELF(gen[1018]),
			.cell_state(gen[1018])
		); 

/******************* CELL 1019 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1019 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[923]),
			.N(gen[924]),
			.NE(gen[925]),

			.O(gen[1018]),
			.E(gen[1020]),

			.SO(gen[1113]),
			.S(gen[1114]),
			.SE(gen[1115]),

			.SELF(gen[1019]),
			.cell_state(gen[1019])
		); 

/******************* CELL 1020 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1020 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[924]),
			.N(gen[925]),
			.NE(gen[926]),

			.O(gen[1019]),
			.E(gen[1021]),

			.SO(gen[1114]),
			.S(gen[1115]),
			.SE(gen[1116]),

			.SELF(gen[1020]),
			.cell_state(gen[1020])
		); 

/******************* CELL 1021 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1021 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[925]),
			.N(gen[926]),
			.NE(gen[927]),

			.O(gen[1020]),
			.E(gen[1022]),

			.SO(gen[1115]),
			.S(gen[1116]),
			.SE(gen[1117]),

			.SELF(gen[1021]),
			.cell_state(gen[1021])
		); 

/******************* CELL 1022 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1022 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[926]),
			.N(gen[927]),
			.NE(gen[928]),

			.O(gen[1021]),
			.E(gen[1023]),

			.SO(gen[1116]),
			.S(gen[1117]),
			.SE(gen[1118]),

			.SELF(gen[1022]),
			.cell_state(gen[1022])
		); 

/******************* CELL 1023 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1023 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[927]),
			.N(gen[928]),
			.NE(gen[929]),

			.O(gen[1022]),
			.E(gen[1024]),

			.SO(gen[1117]),
			.S(gen[1118]),
			.SE(gen[1119]),

			.SELF(gen[1023]),
			.cell_state(gen[1023])
		); 

/******************* CELL 1024 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1024 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[928]),
			.N(gen[929]),
			.NE(gen[930]),

			.O(gen[1023]),
			.E(gen[1025]),

			.SO(gen[1118]),
			.S(gen[1119]),
			.SE(gen[1120]),

			.SELF(gen[1024]),
			.cell_state(gen[1024])
		); 

/******************* CELL 1025 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1025 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[929]),
			.N(gen[930]),
			.NE(gen[931]),

			.O(gen[1024]),
			.E(gen[1026]),

			.SO(gen[1119]),
			.S(gen[1120]),
			.SE(gen[1121]),

			.SELF(gen[1025]),
			.cell_state(gen[1025])
		); 

/******************* CELL 1026 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1026 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[930]),
			.N(gen[931]),
			.NE(gen[932]),

			.O(gen[1025]),
			.E(gen[1027]),

			.SO(gen[1120]),
			.S(gen[1121]),
			.SE(gen[1122]),

			.SELF(gen[1026]),
			.cell_state(gen[1026])
		); 

/******************* CELL 1027 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1027 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[931]),
			.N(gen[932]),
			.NE(gen[933]),

			.O(gen[1026]),
			.E(gen[1028]),

			.SO(gen[1121]),
			.S(gen[1122]),
			.SE(gen[1123]),

			.SELF(gen[1027]),
			.cell_state(gen[1027])
		); 

/******************* CELL 1028 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1028 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[932]),
			.N(gen[933]),
			.NE(gen[934]),

			.O(gen[1027]),
			.E(gen[1029]),

			.SO(gen[1122]),
			.S(gen[1123]),
			.SE(gen[1124]),

			.SELF(gen[1028]),
			.cell_state(gen[1028])
		); 

/******************* CELL 1029 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1029 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[933]),
			.N(gen[934]),
			.NE(gen[935]),

			.O(gen[1028]),
			.E(gen[1030]),

			.SO(gen[1123]),
			.S(gen[1124]),
			.SE(gen[1125]),

			.SELF(gen[1029]),
			.cell_state(gen[1029])
		); 

/******************* CELL 1030 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1030 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[934]),
			.N(gen[935]),
			.NE(gen[936]),

			.O(gen[1029]),
			.E(gen[1031]),

			.SO(gen[1124]),
			.S(gen[1125]),
			.SE(gen[1126]),

			.SELF(gen[1030]),
			.cell_state(gen[1030])
		); 

/******************* CELL 1031 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1031 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[935]),
			.N(gen[936]),
			.NE(gen[937]),

			.O(gen[1030]),
			.E(gen[1032]),

			.SO(gen[1125]),
			.S(gen[1126]),
			.SE(gen[1127]),

			.SELF(gen[1031]),
			.cell_state(gen[1031])
		); 

/******************* CELL 1032 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1032 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[936]),
			.N(gen[937]),
			.NE(gen[938]),

			.O(gen[1031]),
			.E(gen[1033]),

			.SO(gen[1126]),
			.S(gen[1127]),
			.SE(gen[1128]),

			.SELF(gen[1032]),
			.cell_state(gen[1032])
		); 

/******************* CELL 1033 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1033 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[937]),
			.N(gen[938]),
			.NE(gen[939]),

			.O(gen[1032]),
			.E(gen[1034]),

			.SO(gen[1127]),
			.S(gen[1128]),
			.SE(gen[1129]),

			.SELF(gen[1033]),
			.cell_state(gen[1033])
		); 

/******************* CELL 1034 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1034 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[938]),
			.N(gen[939]),
			.NE(gen[940]),

			.O(gen[1033]),
			.E(gen[1035]),

			.SO(gen[1128]),
			.S(gen[1129]),
			.SE(gen[1130]),

			.SELF(gen[1034]),
			.cell_state(gen[1034])
		); 

/******************* CELL 1035 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1035 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[939]),
			.N(gen[940]),
			.NE(gen[941]),

			.O(gen[1034]),
			.E(gen[1036]),

			.SO(gen[1129]),
			.S(gen[1130]),
			.SE(gen[1131]),

			.SELF(gen[1035]),
			.cell_state(gen[1035])
		); 

/******************* CELL 1036 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1036 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[940]),
			.N(gen[941]),
			.NE(gen[942]),

			.O(gen[1035]),
			.E(gen[1037]),

			.SO(gen[1130]),
			.S(gen[1131]),
			.SE(gen[1132]),

			.SELF(gen[1036]),
			.cell_state(gen[1036])
		); 

/******************* CELL 1037 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1037 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[941]),
			.N(gen[942]),
			.NE(gen[943]),

			.O(gen[1036]),
			.E(gen[1038]),

			.SO(gen[1131]),
			.S(gen[1132]),
			.SE(gen[1133]),

			.SELF(gen[1037]),
			.cell_state(gen[1037])
		); 

/******************* CELL 1038 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1038 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[942]),
			.N(gen[943]),
			.NE(gen[944]),

			.O(gen[1037]),
			.E(gen[1039]),

			.SO(gen[1132]),
			.S(gen[1133]),
			.SE(gen[1134]),

			.SELF(gen[1038]),
			.cell_state(gen[1038])
		); 

/******************* CELL 1039 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1039 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[943]),
			.N(gen[944]),
			.NE(gen[945]),

			.O(gen[1038]),
			.E(gen[1040]),

			.SO(gen[1133]),
			.S(gen[1134]),
			.SE(gen[1135]),

			.SELF(gen[1039]),
			.cell_state(gen[1039])
		); 

/******************* CELL 1040 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1040 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[944]),
			.N(gen[945]),
			.NE(gen[946]),

			.O(gen[1039]),
			.E(gen[1041]),

			.SO(gen[1134]),
			.S(gen[1135]),
			.SE(gen[1136]),

			.SELF(gen[1040]),
			.cell_state(gen[1040])
		); 

/******************* CELL 1041 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1041 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[945]),
			.N(gen[946]),
			.NE(gen[947]),

			.O(gen[1040]),
			.E(gen[1042]),

			.SO(gen[1135]),
			.S(gen[1136]),
			.SE(gen[1137]),

			.SELF(gen[1041]),
			.cell_state(gen[1041])
		); 

/******************* CELL 1042 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1042 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[946]),
			.N(gen[947]),
			.NE(gen[948]),

			.O(gen[1041]),
			.E(gen[1043]),

			.SO(gen[1136]),
			.S(gen[1137]),
			.SE(gen[1138]),

			.SELF(gen[1042]),
			.cell_state(gen[1042])
		); 

/******************* CELL 1043 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1043 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[947]),
			.N(gen[948]),
			.NE(gen[949]),

			.O(gen[1042]),
			.E(gen[1044]),

			.SO(gen[1137]),
			.S(gen[1138]),
			.SE(gen[1139]),

			.SELF(gen[1043]),
			.cell_state(gen[1043])
		); 

/******************* CELL 1044 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1044 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[948]),
			.N(gen[949]),
			.NE(gen[948]),

			.O(gen[1043]),
			.E(gen[1043]),

			.SO(gen[1138]),
			.S(gen[1139]),
			.SE(gen[1138]),

			.SELF(gen[1044]),
			.cell_state(gen[1044])
		); 

/******************* CELL 1045 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1045 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[951]),
			.N(gen[950]),
			.NE(gen[951]),

			.O(gen[1046]),
			.E(gen[1046]),

			.SO(gen[1141]),
			.S(gen[1140]),
			.SE(gen[1141]),

			.SELF(gen[1045]),
			.cell_state(gen[1045])
		); 

/******************* CELL 1046 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1046 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[950]),
			.N(gen[951]),
			.NE(gen[952]),

			.O(gen[1045]),
			.E(gen[1047]),

			.SO(gen[1140]),
			.S(gen[1141]),
			.SE(gen[1142]),

			.SELF(gen[1046]),
			.cell_state(gen[1046])
		); 

/******************* CELL 1047 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1047 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[951]),
			.N(gen[952]),
			.NE(gen[953]),

			.O(gen[1046]),
			.E(gen[1048]),

			.SO(gen[1141]),
			.S(gen[1142]),
			.SE(gen[1143]),

			.SELF(gen[1047]),
			.cell_state(gen[1047])
		); 

/******************* CELL 1048 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1048 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[952]),
			.N(gen[953]),
			.NE(gen[954]),

			.O(gen[1047]),
			.E(gen[1049]),

			.SO(gen[1142]),
			.S(gen[1143]),
			.SE(gen[1144]),

			.SELF(gen[1048]),
			.cell_state(gen[1048])
		); 

/******************* CELL 1049 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1049 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[953]),
			.N(gen[954]),
			.NE(gen[955]),

			.O(gen[1048]),
			.E(gen[1050]),

			.SO(gen[1143]),
			.S(gen[1144]),
			.SE(gen[1145]),

			.SELF(gen[1049]),
			.cell_state(gen[1049])
		); 

/******************* CELL 1050 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1050 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[954]),
			.N(gen[955]),
			.NE(gen[956]),

			.O(gen[1049]),
			.E(gen[1051]),

			.SO(gen[1144]),
			.S(gen[1145]),
			.SE(gen[1146]),

			.SELF(gen[1050]),
			.cell_state(gen[1050])
		); 

/******************* CELL 1051 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1051 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[955]),
			.N(gen[956]),
			.NE(gen[957]),

			.O(gen[1050]),
			.E(gen[1052]),

			.SO(gen[1145]),
			.S(gen[1146]),
			.SE(gen[1147]),

			.SELF(gen[1051]),
			.cell_state(gen[1051])
		); 

/******************* CELL 1052 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1052 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[956]),
			.N(gen[957]),
			.NE(gen[958]),

			.O(gen[1051]),
			.E(gen[1053]),

			.SO(gen[1146]),
			.S(gen[1147]),
			.SE(gen[1148]),

			.SELF(gen[1052]),
			.cell_state(gen[1052])
		); 

/******************* CELL 1053 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1053 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[957]),
			.N(gen[958]),
			.NE(gen[959]),

			.O(gen[1052]),
			.E(gen[1054]),

			.SO(gen[1147]),
			.S(gen[1148]),
			.SE(gen[1149]),

			.SELF(gen[1053]),
			.cell_state(gen[1053])
		); 

/******************* CELL 1054 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1054 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[958]),
			.N(gen[959]),
			.NE(gen[960]),

			.O(gen[1053]),
			.E(gen[1055]),

			.SO(gen[1148]),
			.S(gen[1149]),
			.SE(gen[1150]),

			.SELF(gen[1054]),
			.cell_state(gen[1054])
		); 

/******************* CELL 1055 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1055 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[959]),
			.N(gen[960]),
			.NE(gen[961]),

			.O(gen[1054]),
			.E(gen[1056]),

			.SO(gen[1149]),
			.S(gen[1150]),
			.SE(gen[1151]),

			.SELF(gen[1055]),
			.cell_state(gen[1055])
		); 

/******************* CELL 1056 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1056 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[960]),
			.N(gen[961]),
			.NE(gen[962]),

			.O(gen[1055]),
			.E(gen[1057]),

			.SO(gen[1150]),
			.S(gen[1151]),
			.SE(gen[1152]),

			.SELF(gen[1056]),
			.cell_state(gen[1056])
		); 

/******************* CELL 1057 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1057 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[961]),
			.N(gen[962]),
			.NE(gen[963]),

			.O(gen[1056]),
			.E(gen[1058]),

			.SO(gen[1151]),
			.S(gen[1152]),
			.SE(gen[1153]),

			.SELF(gen[1057]),
			.cell_state(gen[1057])
		); 

/******************* CELL 1058 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1058 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[962]),
			.N(gen[963]),
			.NE(gen[964]),

			.O(gen[1057]),
			.E(gen[1059]),

			.SO(gen[1152]),
			.S(gen[1153]),
			.SE(gen[1154]),

			.SELF(gen[1058]),
			.cell_state(gen[1058])
		); 

/******************* CELL 1059 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1059 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[963]),
			.N(gen[964]),
			.NE(gen[965]),

			.O(gen[1058]),
			.E(gen[1060]),

			.SO(gen[1153]),
			.S(gen[1154]),
			.SE(gen[1155]),

			.SELF(gen[1059]),
			.cell_state(gen[1059])
		); 

/******************* CELL 1060 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1060 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[964]),
			.N(gen[965]),
			.NE(gen[966]),

			.O(gen[1059]),
			.E(gen[1061]),

			.SO(gen[1154]),
			.S(gen[1155]),
			.SE(gen[1156]),

			.SELF(gen[1060]),
			.cell_state(gen[1060])
		); 

/******************* CELL 1061 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1061 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[965]),
			.N(gen[966]),
			.NE(gen[967]),

			.O(gen[1060]),
			.E(gen[1062]),

			.SO(gen[1155]),
			.S(gen[1156]),
			.SE(gen[1157]),

			.SELF(gen[1061]),
			.cell_state(gen[1061])
		); 

/******************* CELL 1062 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1062 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[966]),
			.N(gen[967]),
			.NE(gen[968]),

			.O(gen[1061]),
			.E(gen[1063]),

			.SO(gen[1156]),
			.S(gen[1157]),
			.SE(gen[1158]),

			.SELF(gen[1062]),
			.cell_state(gen[1062])
		); 

/******************* CELL 1063 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1063 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[967]),
			.N(gen[968]),
			.NE(gen[969]),

			.O(gen[1062]),
			.E(gen[1064]),

			.SO(gen[1157]),
			.S(gen[1158]),
			.SE(gen[1159]),

			.SELF(gen[1063]),
			.cell_state(gen[1063])
		); 

/******************* CELL 1064 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1064 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[968]),
			.N(gen[969]),
			.NE(gen[970]),

			.O(gen[1063]),
			.E(gen[1065]),

			.SO(gen[1158]),
			.S(gen[1159]),
			.SE(gen[1160]),

			.SELF(gen[1064]),
			.cell_state(gen[1064])
		); 

/******************* CELL 1065 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1065 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[969]),
			.N(gen[970]),
			.NE(gen[971]),

			.O(gen[1064]),
			.E(gen[1066]),

			.SO(gen[1159]),
			.S(gen[1160]),
			.SE(gen[1161]),

			.SELF(gen[1065]),
			.cell_state(gen[1065])
		); 

/******************* CELL 1066 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1066 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[970]),
			.N(gen[971]),
			.NE(gen[972]),

			.O(gen[1065]),
			.E(gen[1067]),

			.SO(gen[1160]),
			.S(gen[1161]),
			.SE(gen[1162]),

			.SELF(gen[1066]),
			.cell_state(gen[1066])
		); 

/******************* CELL 1067 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1067 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[971]),
			.N(gen[972]),
			.NE(gen[973]),

			.O(gen[1066]),
			.E(gen[1068]),

			.SO(gen[1161]),
			.S(gen[1162]),
			.SE(gen[1163]),

			.SELF(gen[1067]),
			.cell_state(gen[1067])
		); 

/******************* CELL 1068 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1068 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[972]),
			.N(gen[973]),
			.NE(gen[974]),

			.O(gen[1067]),
			.E(gen[1069]),

			.SO(gen[1162]),
			.S(gen[1163]),
			.SE(gen[1164]),

			.SELF(gen[1068]),
			.cell_state(gen[1068])
		); 

/******************* CELL 1069 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1069 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[973]),
			.N(gen[974]),
			.NE(gen[975]),

			.O(gen[1068]),
			.E(gen[1070]),

			.SO(gen[1163]),
			.S(gen[1164]),
			.SE(gen[1165]),

			.SELF(gen[1069]),
			.cell_state(gen[1069])
		); 

/******************* CELL 1070 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1070 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[974]),
			.N(gen[975]),
			.NE(gen[976]),

			.O(gen[1069]),
			.E(gen[1071]),

			.SO(gen[1164]),
			.S(gen[1165]),
			.SE(gen[1166]),

			.SELF(gen[1070]),
			.cell_state(gen[1070])
		); 

/******************* CELL 1071 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1071 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[975]),
			.N(gen[976]),
			.NE(gen[977]),

			.O(gen[1070]),
			.E(gen[1072]),

			.SO(gen[1165]),
			.S(gen[1166]),
			.SE(gen[1167]),

			.SELF(gen[1071]),
			.cell_state(gen[1071])
		); 

/******************* CELL 1072 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1072 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[976]),
			.N(gen[977]),
			.NE(gen[978]),

			.O(gen[1071]),
			.E(gen[1073]),

			.SO(gen[1166]),
			.S(gen[1167]),
			.SE(gen[1168]),

			.SELF(gen[1072]),
			.cell_state(gen[1072])
		); 

/******************* CELL 1073 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1073 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[977]),
			.N(gen[978]),
			.NE(gen[979]),

			.O(gen[1072]),
			.E(gen[1074]),

			.SO(gen[1167]),
			.S(gen[1168]),
			.SE(gen[1169]),

			.SELF(gen[1073]),
			.cell_state(gen[1073])
		); 

/******************* CELL 1074 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1074 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[978]),
			.N(gen[979]),
			.NE(gen[980]),

			.O(gen[1073]),
			.E(gen[1075]),

			.SO(gen[1168]),
			.S(gen[1169]),
			.SE(gen[1170]),

			.SELF(gen[1074]),
			.cell_state(gen[1074])
		); 

/******************* CELL 1075 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1075 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[979]),
			.N(gen[980]),
			.NE(gen[981]),

			.O(gen[1074]),
			.E(gen[1076]),

			.SO(gen[1169]),
			.S(gen[1170]),
			.SE(gen[1171]),

			.SELF(gen[1075]),
			.cell_state(gen[1075])
		); 

/******************* CELL 1076 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1076 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[980]),
			.N(gen[981]),
			.NE(gen[982]),

			.O(gen[1075]),
			.E(gen[1077]),

			.SO(gen[1170]),
			.S(gen[1171]),
			.SE(gen[1172]),

			.SELF(gen[1076]),
			.cell_state(gen[1076])
		); 

/******************* CELL 1077 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1077 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[981]),
			.N(gen[982]),
			.NE(gen[983]),

			.O(gen[1076]),
			.E(gen[1078]),

			.SO(gen[1171]),
			.S(gen[1172]),
			.SE(gen[1173]),

			.SELF(gen[1077]),
			.cell_state(gen[1077])
		); 

/******************* CELL 1078 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1078 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[982]),
			.N(gen[983]),
			.NE(gen[984]),

			.O(gen[1077]),
			.E(gen[1079]),

			.SO(gen[1172]),
			.S(gen[1173]),
			.SE(gen[1174]),

			.SELF(gen[1078]),
			.cell_state(gen[1078])
		); 

/******************* CELL 1079 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1079 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[983]),
			.N(gen[984]),
			.NE(gen[985]),

			.O(gen[1078]),
			.E(gen[1080]),

			.SO(gen[1173]),
			.S(gen[1174]),
			.SE(gen[1175]),

			.SELF(gen[1079]),
			.cell_state(gen[1079])
		); 

/******************* CELL 1080 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1080 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[984]),
			.N(gen[985]),
			.NE(gen[986]),

			.O(gen[1079]),
			.E(gen[1081]),

			.SO(gen[1174]),
			.S(gen[1175]),
			.SE(gen[1176]),

			.SELF(gen[1080]),
			.cell_state(gen[1080])
		); 

/******************* CELL 1081 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1081 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[985]),
			.N(gen[986]),
			.NE(gen[987]),

			.O(gen[1080]),
			.E(gen[1082]),

			.SO(gen[1175]),
			.S(gen[1176]),
			.SE(gen[1177]),

			.SELF(gen[1081]),
			.cell_state(gen[1081])
		); 

/******************* CELL 1082 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1082 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[986]),
			.N(gen[987]),
			.NE(gen[988]),

			.O(gen[1081]),
			.E(gen[1083]),

			.SO(gen[1176]),
			.S(gen[1177]),
			.SE(gen[1178]),

			.SELF(gen[1082]),
			.cell_state(gen[1082])
		); 

/******************* CELL 1083 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1083 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[987]),
			.N(gen[988]),
			.NE(gen[989]),

			.O(gen[1082]),
			.E(gen[1084]),

			.SO(gen[1177]),
			.S(gen[1178]),
			.SE(gen[1179]),

			.SELF(gen[1083]),
			.cell_state(gen[1083])
		); 

/******************* CELL 1084 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1084 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[988]),
			.N(gen[989]),
			.NE(gen[990]),

			.O(gen[1083]),
			.E(gen[1085]),

			.SO(gen[1178]),
			.S(gen[1179]),
			.SE(gen[1180]),

			.SELF(gen[1084]),
			.cell_state(gen[1084])
		); 

/******************* CELL 1085 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1085 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[989]),
			.N(gen[990]),
			.NE(gen[991]),

			.O(gen[1084]),
			.E(gen[1086]),

			.SO(gen[1179]),
			.S(gen[1180]),
			.SE(gen[1181]),

			.SELF(gen[1085]),
			.cell_state(gen[1085])
		); 

/******************* CELL 1086 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1086 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[990]),
			.N(gen[991]),
			.NE(gen[992]),

			.O(gen[1085]),
			.E(gen[1087]),

			.SO(gen[1180]),
			.S(gen[1181]),
			.SE(gen[1182]),

			.SELF(gen[1086]),
			.cell_state(gen[1086])
		); 

/******************* CELL 1087 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1087 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[991]),
			.N(gen[992]),
			.NE(gen[993]),

			.O(gen[1086]),
			.E(gen[1088]),

			.SO(gen[1181]),
			.S(gen[1182]),
			.SE(gen[1183]),

			.SELF(gen[1087]),
			.cell_state(gen[1087])
		); 

/******************* CELL 1088 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1088 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[992]),
			.N(gen[993]),
			.NE(gen[994]),

			.O(gen[1087]),
			.E(gen[1089]),

			.SO(gen[1182]),
			.S(gen[1183]),
			.SE(gen[1184]),

			.SELF(gen[1088]),
			.cell_state(gen[1088])
		); 

/******************* CELL 1089 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1089 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[993]),
			.N(gen[994]),
			.NE(gen[995]),

			.O(gen[1088]),
			.E(gen[1090]),

			.SO(gen[1183]),
			.S(gen[1184]),
			.SE(gen[1185]),

			.SELF(gen[1089]),
			.cell_state(gen[1089])
		); 

/******************* CELL 1090 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1090 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[994]),
			.N(gen[995]),
			.NE(gen[996]),

			.O(gen[1089]),
			.E(gen[1091]),

			.SO(gen[1184]),
			.S(gen[1185]),
			.SE(gen[1186]),

			.SELF(gen[1090]),
			.cell_state(gen[1090])
		); 

/******************* CELL 1091 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1091 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[995]),
			.N(gen[996]),
			.NE(gen[997]),

			.O(gen[1090]),
			.E(gen[1092]),

			.SO(gen[1185]),
			.S(gen[1186]),
			.SE(gen[1187]),

			.SELF(gen[1091]),
			.cell_state(gen[1091])
		); 

/******************* CELL 1092 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1092 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[996]),
			.N(gen[997]),
			.NE(gen[998]),

			.O(gen[1091]),
			.E(gen[1093]),

			.SO(gen[1186]),
			.S(gen[1187]),
			.SE(gen[1188]),

			.SELF(gen[1092]),
			.cell_state(gen[1092])
		); 

/******************* CELL 1093 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1093 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[997]),
			.N(gen[998]),
			.NE(gen[999]),

			.O(gen[1092]),
			.E(gen[1094]),

			.SO(gen[1187]),
			.S(gen[1188]),
			.SE(gen[1189]),

			.SELF(gen[1093]),
			.cell_state(gen[1093])
		); 

/******************* CELL 1094 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1094 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[998]),
			.N(gen[999]),
			.NE(gen[1000]),

			.O(gen[1093]),
			.E(gen[1095]),

			.SO(gen[1188]),
			.S(gen[1189]),
			.SE(gen[1190]),

			.SELF(gen[1094]),
			.cell_state(gen[1094])
		); 

/******************* CELL 1095 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1095 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[999]),
			.N(gen[1000]),
			.NE(gen[1001]),

			.O(gen[1094]),
			.E(gen[1096]),

			.SO(gen[1189]),
			.S(gen[1190]),
			.SE(gen[1191]),

			.SELF(gen[1095]),
			.cell_state(gen[1095])
		); 

/******************* CELL 1096 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1096 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1000]),
			.N(gen[1001]),
			.NE(gen[1002]),

			.O(gen[1095]),
			.E(gen[1097]),

			.SO(gen[1190]),
			.S(gen[1191]),
			.SE(gen[1192]),

			.SELF(gen[1096]),
			.cell_state(gen[1096])
		); 

/******************* CELL 1097 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1097 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1001]),
			.N(gen[1002]),
			.NE(gen[1003]),

			.O(gen[1096]),
			.E(gen[1098]),

			.SO(gen[1191]),
			.S(gen[1192]),
			.SE(gen[1193]),

			.SELF(gen[1097]),
			.cell_state(gen[1097])
		); 

/******************* CELL 1098 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1098 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1002]),
			.N(gen[1003]),
			.NE(gen[1004]),

			.O(gen[1097]),
			.E(gen[1099]),

			.SO(gen[1192]),
			.S(gen[1193]),
			.SE(gen[1194]),

			.SELF(gen[1098]),
			.cell_state(gen[1098])
		); 

/******************* CELL 1099 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1099 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1003]),
			.N(gen[1004]),
			.NE(gen[1005]),

			.O(gen[1098]),
			.E(gen[1100]),

			.SO(gen[1193]),
			.S(gen[1194]),
			.SE(gen[1195]),

			.SELF(gen[1099]),
			.cell_state(gen[1099])
		); 

/******************* CELL 1100 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1100 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1004]),
			.N(gen[1005]),
			.NE(gen[1006]),

			.O(gen[1099]),
			.E(gen[1101]),

			.SO(gen[1194]),
			.S(gen[1195]),
			.SE(gen[1196]),

			.SELF(gen[1100]),
			.cell_state(gen[1100])
		); 

/******************* CELL 1101 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1101 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1005]),
			.N(gen[1006]),
			.NE(gen[1007]),

			.O(gen[1100]),
			.E(gen[1102]),

			.SO(gen[1195]),
			.S(gen[1196]),
			.SE(gen[1197]),

			.SELF(gen[1101]),
			.cell_state(gen[1101])
		); 

/******************* CELL 1102 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1102 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1006]),
			.N(gen[1007]),
			.NE(gen[1008]),

			.O(gen[1101]),
			.E(gen[1103]),

			.SO(gen[1196]),
			.S(gen[1197]),
			.SE(gen[1198]),

			.SELF(gen[1102]),
			.cell_state(gen[1102])
		); 

/******************* CELL 1103 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1103 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1007]),
			.N(gen[1008]),
			.NE(gen[1009]),

			.O(gen[1102]),
			.E(gen[1104]),

			.SO(gen[1197]),
			.S(gen[1198]),
			.SE(gen[1199]),

			.SELF(gen[1103]),
			.cell_state(gen[1103])
		); 

/******************* CELL 1104 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1104 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1008]),
			.N(gen[1009]),
			.NE(gen[1010]),

			.O(gen[1103]),
			.E(gen[1105]),

			.SO(gen[1198]),
			.S(gen[1199]),
			.SE(gen[1200]),

			.SELF(gen[1104]),
			.cell_state(gen[1104])
		); 

/******************* CELL 1105 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1105 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1009]),
			.N(gen[1010]),
			.NE(gen[1011]),

			.O(gen[1104]),
			.E(gen[1106]),

			.SO(gen[1199]),
			.S(gen[1200]),
			.SE(gen[1201]),

			.SELF(gen[1105]),
			.cell_state(gen[1105])
		); 

/******************* CELL 1106 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1106 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1010]),
			.N(gen[1011]),
			.NE(gen[1012]),

			.O(gen[1105]),
			.E(gen[1107]),

			.SO(gen[1200]),
			.S(gen[1201]),
			.SE(gen[1202]),

			.SELF(gen[1106]),
			.cell_state(gen[1106])
		); 

/******************* CELL 1107 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1107 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1011]),
			.N(gen[1012]),
			.NE(gen[1013]),

			.O(gen[1106]),
			.E(gen[1108]),

			.SO(gen[1201]),
			.S(gen[1202]),
			.SE(gen[1203]),

			.SELF(gen[1107]),
			.cell_state(gen[1107])
		); 

/******************* CELL 1108 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1108 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1012]),
			.N(gen[1013]),
			.NE(gen[1014]),

			.O(gen[1107]),
			.E(gen[1109]),

			.SO(gen[1202]),
			.S(gen[1203]),
			.SE(gen[1204]),

			.SELF(gen[1108]),
			.cell_state(gen[1108])
		); 

/******************* CELL 1109 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1109 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1013]),
			.N(gen[1014]),
			.NE(gen[1015]),

			.O(gen[1108]),
			.E(gen[1110]),

			.SO(gen[1203]),
			.S(gen[1204]),
			.SE(gen[1205]),

			.SELF(gen[1109]),
			.cell_state(gen[1109])
		); 

/******************* CELL 1110 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1110 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1014]),
			.N(gen[1015]),
			.NE(gen[1016]),

			.O(gen[1109]),
			.E(gen[1111]),

			.SO(gen[1204]),
			.S(gen[1205]),
			.SE(gen[1206]),

			.SELF(gen[1110]),
			.cell_state(gen[1110])
		); 

/******************* CELL 1111 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1111 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1015]),
			.N(gen[1016]),
			.NE(gen[1017]),

			.O(gen[1110]),
			.E(gen[1112]),

			.SO(gen[1205]),
			.S(gen[1206]),
			.SE(gen[1207]),

			.SELF(gen[1111]),
			.cell_state(gen[1111])
		); 

/******************* CELL 1112 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1112 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1016]),
			.N(gen[1017]),
			.NE(gen[1018]),

			.O(gen[1111]),
			.E(gen[1113]),

			.SO(gen[1206]),
			.S(gen[1207]),
			.SE(gen[1208]),

			.SELF(gen[1112]),
			.cell_state(gen[1112])
		); 

/******************* CELL 1113 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1113 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1017]),
			.N(gen[1018]),
			.NE(gen[1019]),

			.O(gen[1112]),
			.E(gen[1114]),

			.SO(gen[1207]),
			.S(gen[1208]),
			.SE(gen[1209]),

			.SELF(gen[1113]),
			.cell_state(gen[1113])
		); 

/******************* CELL 1114 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1114 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1018]),
			.N(gen[1019]),
			.NE(gen[1020]),

			.O(gen[1113]),
			.E(gen[1115]),

			.SO(gen[1208]),
			.S(gen[1209]),
			.SE(gen[1210]),

			.SELF(gen[1114]),
			.cell_state(gen[1114])
		); 

/******************* CELL 1115 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1115 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1019]),
			.N(gen[1020]),
			.NE(gen[1021]),

			.O(gen[1114]),
			.E(gen[1116]),

			.SO(gen[1209]),
			.S(gen[1210]),
			.SE(gen[1211]),

			.SELF(gen[1115]),
			.cell_state(gen[1115])
		); 

/******************* CELL 1116 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1116 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1020]),
			.N(gen[1021]),
			.NE(gen[1022]),

			.O(gen[1115]),
			.E(gen[1117]),

			.SO(gen[1210]),
			.S(gen[1211]),
			.SE(gen[1212]),

			.SELF(gen[1116]),
			.cell_state(gen[1116])
		); 

/******************* CELL 1117 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1117 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1021]),
			.N(gen[1022]),
			.NE(gen[1023]),

			.O(gen[1116]),
			.E(gen[1118]),

			.SO(gen[1211]),
			.S(gen[1212]),
			.SE(gen[1213]),

			.SELF(gen[1117]),
			.cell_state(gen[1117])
		); 

/******************* CELL 1118 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1118 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1022]),
			.N(gen[1023]),
			.NE(gen[1024]),

			.O(gen[1117]),
			.E(gen[1119]),

			.SO(gen[1212]),
			.S(gen[1213]),
			.SE(gen[1214]),

			.SELF(gen[1118]),
			.cell_state(gen[1118])
		); 

/******************* CELL 1119 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1119 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1023]),
			.N(gen[1024]),
			.NE(gen[1025]),

			.O(gen[1118]),
			.E(gen[1120]),

			.SO(gen[1213]),
			.S(gen[1214]),
			.SE(gen[1215]),

			.SELF(gen[1119]),
			.cell_state(gen[1119])
		); 

/******************* CELL 1120 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1120 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1024]),
			.N(gen[1025]),
			.NE(gen[1026]),

			.O(gen[1119]),
			.E(gen[1121]),

			.SO(gen[1214]),
			.S(gen[1215]),
			.SE(gen[1216]),

			.SELF(gen[1120]),
			.cell_state(gen[1120])
		); 

/******************* CELL 1121 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1121 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1025]),
			.N(gen[1026]),
			.NE(gen[1027]),

			.O(gen[1120]),
			.E(gen[1122]),

			.SO(gen[1215]),
			.S(gen[1216]),
			.SE(gen[1217]),

			.SELF(gen[1121]),
			.cell_state(gen[1121])
		); 

/******************* CELL 1122 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1122 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1026]),
			.N(gen[1027]),
			.NE(gen[1028]),

			.O(gen[1121]),
			.E(gen[1123]),

			.SO(gen[1216]),
			.S(gen[1217]),
			.SE(gen[1218]),

			.SELF(gen[1122]),
			.cell_state(gen[1122])
		); 

/******************* CELL 1123 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1123 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1027]),
			.N(gen[1028]),
			.NE(gen[1029]),

			.O(gen[1122]),
			.E(gen[1124]),

			.SO(gen[1217]),
			.S(gen[1218]),
			.SE(gen[1219]),

			.SELF(gen[1123]),
			.cell_state(gen[1123])
		); 

/******************* CELL 1124 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1124 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1028]),
			.N(gen[1029]),
			.NE(gen[1030]),

			.O(gen[1123]),
			.E(gen[1125]),

			.SO(gen[1218]),
			.S(gen[1219]),
			.SE(gen[1220]),

			.SELF(gen[1124]),
			.cell_state(gen[1124])
		); 

/******************* CELL 1125 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1125 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1029]),
			.N(gen[1030]),
			.NE(gen[1031]),

			.O(gen[1124]),
			.E(gen[1126]),

			.SO(gen[1219]),
			.S(gen[1220]),
			.SE(gen[1221]),

			.SELF(gen[1125]),
			.cell_state(gen[1125])
		); 

/******************* CELL 1126 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1126 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1030]),
			.N(gen[1031]),
			.NE(gen[1032]),

			.O(gen[1125]),
			.E(gen[1127]),

			.SO(gen[1220]),
			.S(gen[1221]),
			.SE(gen[1222]),

			.SELF(gen[1126]),
			.cell_state(gen[1126])
		); 

/******************* CELL 1127 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1127 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1031]),
			.N(gen[1032]),
			.NE(gen[1033]),

			.O(gen[1126]),
			.E(gen[1128]),

			.SO(gen[1221]),
			.S(gen[1222]),
			.SE(gen[1223]),

			.SELF(gen[1127]),
			.cell_state(gen[1127])
		); 

/******************* CELL 1128 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1128 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1032]),
			.N(gen[1033]),
			.NE(gen[1034]),

			.O(gen[1127]),
			.E(gen[1129]),

			.SO(gen[1222]),
			.S(gen[1223]),
			.SE(gen[1224]),

			.SELF(gen[1128]),
			.cell_state(gen[1128])
		); 

/******************* CELL 1129 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1129 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1033]),
			.N(gen[1034]),
			.NE(gen[1035]),

			.O(gen[1128]),
			.E(gen[1130]),

			.SO(gen[1223]),
			.S(gen[1224]),
			.SE(gen[1225]),

			.SELF(gen[1129]),
			.cell_state(gen[1129])
		); 

/******************* CELL 1130 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1130 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1034]),
			.N(gen[1035]),
			.NE(gen[1036]),

			.O(gen[1129]),
			.E(gen[1131]),

			.SO(gen[1224]),
			.S(gen[1225]),
			.SE(gen[1226]),

			.SELF(gen[1130]),
			.cell_state(gen[1130])
		); 

/******************* CELL 1131 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1131 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1035]),
			.N(gen[1036]),
			.NE(gen[1037]),

			.O(gen[1130]),
			.E(gen[1132]),

			.SO(gen[1225]),
			.S(gen[1226]),
			.SE(gen[1227]),

			.SELF(gen[1131]),
			.cell_state(gen[1131])
		); 

/******************* CELL 1132 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1132 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1036]),
			.N(gen[1037]),
			.NE(gen[1038]),

			.O(gen[1131]),
			.E(gen[1133]),

			.SO(gen[1226]),
			.S(gen[1227]),
			.SE(gen[1228]),

			.SELF(gen[1132]),
			.cell_state(gen[1132])
		); 

/******************* CELL 1133 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1133 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1037]),
			.N(gen[1038]),
			.NE(gen[1039]),

			.O(gen[1132]),
			.E(gen[1134]),

			.SO(gen[1227]),
			.S(gen[1228]),
			.SE(gen[1229]),

			.SELF(gen[1133]),
			.cell_state(gen[1133])
		); 

/******************* CELL 1134 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1134 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1038]),
			.N(gen[1039]),
			.NE(gen[1040]),

			.O(gen[1133]),
			.E(gen[1135]),

			.SO(gen[1228]),
			.S(gen[1229]),
			.SE(gen[1230]),

			.SELF(gen[1134]),
			.cell_state(gen[1134])
		); 

/******************* CELL 1135 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1135 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1039]),
			.N(gen[1040]),
			.NE(gen[1041]),

			.O(gen[1134]),
			.E(gen[1136]),

			.SO(gen[1229]),
			.S(gen[1230]),
			.SE(gen[1231]),

			.SELF(gen[1135]),
			.cell_state(gen[1135])
		); 

/******************* CELL 1136 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1136 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1040]),
			.N(gen[1041]),
			.NE(gen[1042]),

			.O(gen[1135]),
			.E(gen[1137]),

			.SO(gen[1230]),
			.S(gen[1231]),
			.SE(gen[1232]),

			.SELF(gen[1136]),
			.cell_state(gen[1136])
		); 

/******************* CELL 1137 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1137 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1041]),
			.N(gen[1042]),
			.NE(gen[1043]),

			.O(gen[1136]),
			.E(gen[1138]),

			.SO(gen[1231]),
			.S(gen[1232]),
			.SE(gen[1233]),

			.SELF(gen[1137]),
			.cell_state(gen[1137])
		); 

/******************* CELL 1138 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1138 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1042]),
			.N(gen[1043]),
			.NE(gen[1044]),

			.O(gen[1137]),
			.E(gen[1139]),

			.SO(gen[1232]),
			.S(gen[1233]),
			.SE(gen[1234]),

			.SELF(gen[1138]),
			.cell_state(gen[1138])
		); 

/******************* CELL 1139 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1139 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1043]),
			.N(gen[1044]),
			.NE(gen[1043]),

			.O(gen[1138]),
			.E(gen[1138]),

			.SO(gen[1233]),
			.S(gen[1234]),
			.SE(gen[1233]),

			.SELF(gen[1139]),
			.cell_state(gen[1139])
		); 

/******************* CELL 1140 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1140 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1046]),
			.N(gen[1045]),
			.NE(gen[1046]),

			.O(gen[1141]),
			.E(gen[1141]),

			.SO(gen[1236]),
			.S(gen[1235]),
			.SE(gen[1236]),

			.SELF(gen[1140]),
			.cell_state(gen[1140])
		); 

/******************* CELL 1141 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1141 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1045]),
			.N(gen[1046]),
			.NE(gen[1047]),

			.O(gen[1140]),
			.E(gen[1142]),

			.SO(gen[1235]),
			.S(gen[1236]),
			.SE(gen[1237]),

			.SELF(gen[1141]),
			.cell_state(gen[1141])
		); 

/******************* CELL 1142 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1142 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1046]),
			.N(gen[1047]),
			.NE(gen[1048]),

			.O(gen[1141]),
			.E(gen[1143]),

			.SO(gen[1236]),
			.S(gen[1237]),
			.SE(gen[1238]),

			.SELF(gen[1142]),
			.cell_state(gen[1142])
		); 

/******************* CELL 1143 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1143 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1047]),
			.N(gen[1048]),
			.NE(gen[1049]),

			.O(gen[1142]),
			.E(gen[1144]),

			.SO(gen[1237]),
			.S(gen[1238]),
			.SE(gen[1239]),

			.SELF(gen[1143]),
			.cell_state(gen[1143])
		); 

/******************* CELL 1144 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1144 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1048]),
			.N(gen[1049]),
			.NE(gen[1050]),

			.O(gen[1143]),
			.E(gen[1145]),

			.SO(gen[1238]),
			.S(gen[1239]),
			.SE(gen[1240]),

			.SELF(gen[1144]),
			.cell_state(gen[1144])
		); 

/******************* CELL 1145 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1145 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1049]),
			.N(gen[1050]),
			.NE(gen[1051]),

			.O(gen[1144]),
			.E(gen[1146]),

			.SO(gen[1239]),
			.S(gen[1240]),
			.SE(gen[1241]),

			.SELF(gen[1145]),
			.cell_state(gen[1145])
		); 

/******************* CELL 1146 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1146 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1050]),
			.N(gen[1051]),
			.NE(gen[1052]),

			.O(gen[1145]),
			.E(gen[1147]),

			.SO(gen[1240]),
			.S(gen[1241]),
			.SE(gen[1242]),

			.SELF(gen[1146]),
			.cell_state(gen[1146])
		); 

/******************* CELL 1147 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1147 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1051]),
			.N(gen[1052]),
			.NE(gen[1053]),

			.O(gen[1146]),
			.E(gen[1148]),

			.SO(gen[1241]),
			.S(gen[1242]),
			.SE(gen[1243]),

			.SELF(gen[1147]),
			.cell_state(gen[1147])
		); 

/******************* CELL 1148 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1148 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1052]),
			.N(gen[1053]),
			.NE(gen[1054]),

			.O(gen[1147]),
			.E(gen[1149]),

			.SO(gen[1242]),
			.S(gen[1243]),
			.SE(gen[1244]),

			.SELF(gen[1148]),
			.cell_state(gen[1148])
		); 

/******************* CELL 1149 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1149 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1053]),
			.N(gen[1054]),
			.NE(gen[1055]),

			.O(gen[1148]),
			.E(gen[1150]),

			.SO(gen[1243]),
			.S(gen[1244]),
			.SE(gen[1245]),

			.SELF(gen[1149]),
			.cell_state(gen[1149])
		); 

/******************* CELL 1150 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1150 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1054]),
			.N(gen[1055]),
			.NE(gen[1056]),

			.O(gen[1149]),
			.E(gen[1151]),

			.SO(gen[1244]),
			.S(gen[1245]),
			.SE(gen[1246]),

			.SELF(gen[1150]),
			.cell_state(gen[1150])
		); 

/******************* CELL 1151 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1151 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1055]),
			.N(gen[1056]),
			.NE(gen[1057]),

			.O(gen[1150]),
			.E(gen[1152]),

			.SO(gen[1245]),
			.S(gen[1246]),
			.SE(gen[1247]),

			.SELF(gen[1151]),
			.cell_state(gen[1151])
		); 

/******************* CELL 1152 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1152 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1056]),
			.N(gen[1057]),
			.NE(gen[1058]),

			.O(gen[1151]),
			.E(gen[1153]),

			.SO(gen[1246]),
			.S(gen[1247]),
			.SE(gen[1248]),

			.SELF(gen[1152]),
			.cell_state(gen[1152])
		); 

/******************* CELL 1153 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1153 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1057]),
			.N(gen[1058]),
			.NE(gen[1059]),

			.O(gen[1152]),
			.E(gen[1154]),

			.SO(gen[1247]),
			.S(gen[1248]),
			.SE(gen[1249]),

			.SELF(gen[1153]),
			.cell_state(gen[1153])
		); 

/******************* CELL 1154 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1154 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1058]),
			.N(gen[1059]),
			.NE(gen[1060]),

			.O(gen[1153]),
			.E(gen[1155]),

			.SO(gen[1248]),
			.S(gen[1249]),
			.SE(gen[1250]),

			.SELF(gen[1154]),
			.cell_state(gen[1154])
		); 

/******************* CELL 1155 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1155 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1059]),
			.N(gen[1060]),
			.NE(gen[1061]),

			.O(gen[1154]),
			.E(gen[1156]),

			.SO(gen[1249]),
			.S(gen[1250]),
			.SE(gen[1251]),

			.SELF(gen[1155]),
			.cell_state(gen[1155])
		); 

/******************* CELL 1156 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1156 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1060]),
			.N(gen[1061]),
			.NE(gen[1062]),

			.O(gen[1155]),
			.E(gen[1157]),

			.SO(gen[1250]),
			.S(gen[1251]),
			.SE(gen[1252]),

			.SELF(gen[1156]),
			.cell_state(gen[1156])
		); 

/******************* CELL 1157 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1157 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1061]),
			.N(gen[1062]),
			.NE(gen[1063]),

			.O(gen[1156]),
			.E(gen[1158]),

			.SO(gen[1251]),
			.S(gen[1252]),
			.SE(gen[1253]),

			.SELF(gen[1157]),
			.cell_state(gen[1157])
		); 

/******************* CELL 1158 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1158 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1062]),
			.N(gen[1063]),
			.NE(gen[1064]),

			.O(gen[1157]),
			.E(gen[1159]),

			.SO(gen[1252]),
			.S(gen[1253]),
			.SE(gen[1254]),

			.SELF(gen[1158]),
			.cell_state(gen[1158])
		); 

/******************* CELL 1159 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1159 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1063]),
			.N(gen[1064]),
			.NE(gen[1065]),

			.O(gen[1158]),
			.E(gen[1160]),

			.SO(gen[1253]),
			.S(gen[1254]),
			.SE(gen[1255]),

			.SELF(gen[1159]),
			.cell_state(gen[1159])
		); 

/******************* CELL 1160 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1160 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1064]),
			.N(gen[1065]),
			.NE(gen[1066]),

			.O(gen[1159]),
			.E(gen[1161]),

			.SO(gen[1254]),
			.S(gen[1255]),
			.SE(gen[1256]),

			.SELF(gen[1160]),
			.cell_state(gen[1160])
		); 

/******************* CELL 1161 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1161 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1065]),
			.N(gen[1066]),
			.NE(gen[1067]),

			.O(gen[1160]),
			.E(gen[1162]),

			.SO(gen[1255]),
			.S(gen[1256]),
			.SE(gen[1257]),

			.SELF(gen[1161]),
			.cell_state(gen[1161])
		); 

/******************* CELL 1162 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1162 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1066]),
			.N(gen[1067]),
			.NE(gen[1068]),

			.O(gen[1161]),
			.E(gen[1163]),

			.SO(gen[1256]),
			.S(gen[1257]),
			.SE(gen[1258]),

			.SELF(gen[1162]),
			.cell_state(gen[1162])
		); 

/******************* CELL 1163 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1163 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1067]),
			.N(gen[1068]),
			.NE(gen[1069]),

			.O(gen[1162]),
			.E(gen[1164]),

			.SO(gen[1257]),
			.S(gen[1258]),
			.SE(gen[1259]),

			.SELF(gen[1163]),
			.cell_state(gen[1163])
		); 

/******************* CELL 1164 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1164 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1068]),
			.N(gen[1069]),
			.NE(gen[1070]),

			.O(gen[1163]),
			.E(gen[1165]),

			.SO(gen[1258]),
			.S(gen[1259]),
			.SE(gen[1260]),

			.SELF(gen[1164]),
			.cell_state(gen[1164])
		); 

/******************* CELL 1165 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1165 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1069]),
			.N(gen[1070]),
			.NE(gen[1071]),

			.O(gen[1164]),
			.E(gen[1166]),

			.SO(gen[1259]),
			.S(gen[1260]),
			.SE(gen[1261]),

			.SELF(gen[1165]),
			.cell_state(gen[1165])
		); 

/******************* CELL 1166 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1166 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1070]),
			.N(gen[1071]),
			.NE(gen[1072]),

			.O(gen[1165]),
			.E(gen[1167]),

			.SO(gen[1260]),
			.S(gen[1261]),
			.SE(gen[1262]),

			.SELF(gen[1166]),
			.cell_state(gen[1166])
		); 

/******************* CELL 1167 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1167 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1071]),
			.N(gen[1072]),
			.NE(gen[1073]),

			.O(gen[1166]),
			.E(gen[1168]),

			.SO(gen[1261]),
			.S(gen[1262]),
			.SE(gen[1263]),

			.SELF(gen[1167]),
			.cell_state(gen[1167])
		); 

/******************* CELL 1168 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1168 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1072]),
			.N(gen[1073]),
			.NE(gen[1074]),

			.O(gen[1167]),
			.E(gen[1169]),

			.SO(gen[1262]),
			.S(gen[1263]),
			.SE(gen[1264]),

			.SELF(gen[1168]),
			.cell_state(gen[1168])
		); 

/******************* CELL 1169 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1169 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1073]),
			.N(gen[1074]),
			.NE(gen[1075]),

			.O(gen[1168]),
			.E(gen[1170]),

			.SO(gen[1263]),
			.S(gen[1264]),
			.SE(gen[1265]),

			.SELF(gen[1169]),
			.cell_state(gen[1169])
		); 

/******************* CELL 1170 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1170 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1074]),
			.N(gen[1075]),
			.NE(gen[1076]),

			.O(gen[1169]),
			.E(gen[1171]),

			.SO(gen[1264]),
			.S(gen[1265]),
			.SE(gen[1266]),

			.SELF(gen[1170]),
			.cell_state(gen[1170])
		); 

/******************* CELL 1171 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1171 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1075]),
			.N(gen[1076]),
			.NE(gen[1077]),

			.O(gen[1170]),
			.E(gen[1172]),

			.SO(gen[1265]),
			.S(gen[1266]),
			.SE(gen[1267]),

			.SELF(gen[1171]),
			.cell_state(gen[1171])
		); 

/******************* CELL 1172 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1172 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1076]),
			.N(gen[1077]),
			.NE(gen[1078]),

			.O(gen[1171]),
			.E(gen[1173]),

			.SO(gen[1266]),
			.S(gen[1267]),
			.SE(gen[1268]),

			.SELF(gen[1172]),
			.cell_state(gen[1172])
		); 

/******************* CELL 1173 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1173 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1077]),
			.N(gen[1078]),
			.NE(gen[1079]),

			.O(gen[1172]),
			.E(gen[1174]),

			.SO(gen[1267]),
			.S(gen[1268]),
			.SE(gen[1269]),

			.SELF(gen[1173]),
			.cell_state(gen[1173])
		); 

/******************* CELL 1174 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1174 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1078]),
			.N(gen[1079]),
			.NE(gen[1080]),

			.O(gen[1173]),
			.E(gen[1175]),

			.SO(gen[1268]),
			.S(gen[1269]),
			.SE(gen[1270]),

			.SELF(gen[1174]),
			.cell_state(gen[1174])
		); 

/******************* CELL 1175 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1175 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1079]),
			.N(gen[1080]),
			.NE(gen[1081]),

			.O(gen[1174]),
			.E(gen[1176]),

			.SO(gen[1269]),
			.S(gen[1270]),
			.SE(gen[1271]),

			.SELF(gen[1175]),
			.cell_state(gen[1175])
		); 

/******************* CELL 1176 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1176 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1080]),
			.N(gen[1081]),
			.NE(gen[1082]),

			.O(gen[1175]),
			.E(gen[1177]),

			.SO(gen[1270]),
			.S(gen[1271]),
			.SE(gen[1272]),

			.SELF(gen[1176]),
			.cell_state(gen[1176])
		); 

/******************* CELL 1177 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1177 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1081]),
			.N(gen[1082]),
			.NE(gen[1083]),

			.O(gen[1176]),
			.E(gen[1178]),

			.SO(gen[1271]),
			.S(gen[1272]),
			.SE(gen[1273]),

			.SELF(gen[1177]),
			.cell_state(gen[1177])
		); 

/******************* CELL 1178 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1178 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1082]),
			.N(gen[1083]),
			.NE(gen[1084]),

			.O(gen[1177]),
			.E(gen[1179]),

			.SO(gen[1272]),
			.S(gen[1273]),
			.SE(gen[1274]),

			.SELF(gen[1178]),
			.cell_state(gen[1178])
		); 

/******************* CELL 1179 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1179 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1083]),
			.N(gen[1084]),
			.NE(gen[1085]),

			.O(gen[1178]),
			.E(gen[1180]),

			.SO(gen[1273]),
			.S(gen[1274]),
			.SE(gen[1275]),

			.SELF(gen[1179]),
			.cell_state(gen[1179])
		); 

/******************* CELL 1180 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1180 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1084]),
			.N(gen[1085]),
			.NE(gen[1086]),

			.O(gen[1179]),
			.E(gen[1181]),

			.SO(gen[1274]),
			.S(gen[1275]),
			.SE(gen[1276]),

			.SELF(gen[1180]),
			.cell_state(gen[1180])
		); 

/******************* CELL 1181 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1181 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1085]),
			.N(gen[1086]),
			.NE(gen[1087]),

			.O(gen[1180]),
			.E(gen[1182]),

			.SO(gen[1275]),
			.S(gen[1276]),
			.SE(gen[1277]),

			.SELF(gen[1181]),
			.cell_state(gen[1181])
		); 

/******************* CELL 1182 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1182 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1086]),
			.N(gen[1087]),
			.NE(gen[1088]),

			.O(gen[1181]),
			.E(gen[1183]),

			.SO(gen[1276]),
			.S(gen[1277]),
			.SE(gen[1278]),

			.SELF(gen[1182]),
			.cell_state(gen[1182])
		); 

/******************* CELL 1183 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1183 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1087]),
			.N(gen[1088]),
			.NE(gen[1089]),

			.O(gen[1182]),
			.E(gen[1184]),

			.SO(gen[1277]),
			.S(gen[1278]),
			.SE(gen[1279]),

			.SELF(gen[1183]),
			.cell_state(gen[1183])
		); 

/******************* CELL 1184 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1184 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1088]),
			.N(gen[1089]),
			.NE(gen[1090]),

			.O(gen[1183]),
			.E(gen[1185]),

			.SO(gen[1278]),
			.S(gen[1279]),
			.SE(gen[1280]),

			.SELF(gen[1184]),
			.cell_state(gen[1184])
		); 

/******************* CELL 1185 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1185 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1089]),
			.N(gen[1090]),
			.NE(gen[1091]),

			.O(gen[1184]),
			.E(gen[1186]),

			.SO(gen[1279]),
			.S(gen[1280]),
			.SE(gen[1281]),

			.SELF(gen[1185]),
			.cell_state(gen[1185])
		); 

/******************* CELL 1186 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1186 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1090]),
			.N(gen[1091]),
			.NE(gen[1092]),

			.O(gen[1185]),
			.E(gen[1187]),

			.SO(gen[1280]),
			.S(gen[1281]),
			.SE(gen[1282]),

			.SELF(gen[1186]),
			.cell_state(gen[1186])
		); 

/******************* CELL 1187 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1187 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1091]),
			.N(gen[1092]),
			.NE(gen[1093]),

			.O(gen[1186]),
			.E(gen[1188]),

			.SO(gen[1281]),
			.S(gen[1282]),
			.SE(gen[1283]),

			.SELF(gen[1187]),
			.cell_state(gen[1187])
		); 

/******************* CELL 1188 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1188 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1092]),
			.N(gen[1093]),
			.NE(gen[1094]),

			.O(gen[1187]),
			.E(gen[1189]),

			.SO(gen[1282]),
			.S(gen[1283]),
			.SE(gen[1284]),

			.SELF(gen[1188]),
			.cell_state(gen[1188])
		); 

/******************* CELL 1189 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1189 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1093]),
			.N(gen[1094]),
			.NE(gen[1095]),

			.O(gen[1188]),
			.E(gen[1190]),

			.SO(gen[1283]),
			.S(gen[1284]),
			.SE(gen[1285]),

			.SELF(gen[1189]),
			.cell_state(gen[1189])
		); 

/******************* CELL 1190 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1190 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1094]),
			.N(gen[1095]),
			.NE(gen[1096]),

			.O(gen[1189]),
			.E(gen[1191]),

			.SO(gen[1284]),
			.S(gen[1285]),
			.SE(gen[1286]),

			.SELF(gen[1190]),
			.cell_state(gen[1190])
		); 

/******************* CELL 1191 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1191 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1095]),
			.N(gen[1096]),
			.NE(gen[1097]),

			.O(gen[1190]),
			.E(gen[1192]),

			.SO(gen[1285]),
			.S(gen[1286]),
			.SE(gen[1287]),

			.SELF(gen[1191]),
			.cell_state(gen[1191])
		); 

/******************* CELL 1192 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1192 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1096]),
			.N(gen[1097]),
			.NE(gen[1098]),

			.O(gen[1191]),
			.E(gen[1193]),

			.SO(gen[1286]),
			.S(gen[1287]),
			.SE(gen[1288]),

			.SELF(gen[1192]),
			.cell_state(gen[1192])
		); 

/******************* CELL 1193 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1193 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1097]),
			.N(gen[1098]),
			.NE(gen[1099]),

			.O(gen[1192]),
			.E(gen[1194]),

			.SO(gen[1287]),
			.S(gen[1288]),
			.SE(gen[1289]),

			.SELF(gen[1193]),
			.cell_state(gen[1193])
		); 

/******************* CELL 1194 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1194 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1098]),
			.N(gen[1099]),
			.NE(gen[1100]),

			.O(gen[1193]),
			.E(gen[1195]),

			.SO(gen[1288]),
			.S(gen[1289]),
			.SE(gen[1290]),

			.SELF(gen[1194]),
			.cell_state(gen[1194])
		); 

/******************* CELL 1195 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1195 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1099]),
			.N(gen[1100]),
			.NE(gen[1101]),

			.O(gen[1194]),
			.E(gen[1196]),

			.SO(gen[1289]),
			.S(gen[1290]),
			.SE(gen[1291]),

			.SELF(gen[1195]),
			.cell_state(gen[1195])
		); 

/******************* CELL 1196 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1196 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1100]),
			.N(gen[1101]),
			.NE(gen[1102]),

			.O(gen[1195]),
			.E(gen[1197]),

			.SO(gen[1290]),
			.S(gen[1291]),
			.SE(gen[1292]),

			.SELF(gen[1196]),
			.cell_state(gen[1196])
		); 

/******************* CELL 1197 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1197 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1101]),
			.N(gen[1102]),
			.NE(gen[1103]),

			.O(gen[1196]),
			.E(gen[1198]),

			.SO(gen[1291]),
			.S(gen[1292]),
			.SE(gen[1293]),

			.SELF(gen[1197]),
			.cell_state(gen[1197])
		); 

/******************* CELL 1198 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1198 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1102]),
			.N(gen[1103]),
			.NE(gen[1104]),

			.O(gen[1197]),
			.E(gen[1199]),

			.SO(gen[1292]),
			.S(gen[1293]),
			.SE(gen[1294]),

			.SELF(gen[1198]),
			.cell_state(gen[1198])
		); 

/******************* CELL 1199 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1199 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1103]),
			.N(gen[1104]),
			.NE(gen[1105]),

			.O(gen[1198]),
			.E(gen[1200]),

			.SO(gen[1293]),
			.S(gen[1294]),
			.SE(gen[1295]),

			.SELF(gen[1199]),
			.cell_state(gen[1199])
		); 

/******************* CELL 1200 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1200 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1104]),
			.N(gen[1105]),
			.NE(gen[1106]),

			.O(gen[1199]),
			.E(gen[1201]),

			.SO(gen[1294]),
			.S(gen[1295]),
			.SE(gen[1296]),

			.SELF(gen[1200]),
			.cell_state(gen[1200])
		); 

/******************* CELL 1201 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1201 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1105]),
			.N(gen[1106]),
			.NE(gen[1107]),

			.O(gen[1200]),
			.E(gen[1202]),

			.SO(gen[1295]),
			.S(gen[1296]),
			.SE(gen[1297]),

			.SELF(gen[1201]),
			.cell_state(gen[1201])
		); 

/******************* CELL 1202 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1202 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1106]),
			.N(gen[1107]),
			.NE(gen[1108]),

			.O(gen[1201]),
			.E(gen[1203]),

			.SO(gen[1296]),
			.S(gen[1297]),
			.SE(gen[1298]),

			.SELF(gen[1202]),
			.cell_state(gen[1202])
		); 

/******************* CELL 1203 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1203 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1107]),
			.N(gen[1108]),
			.NE(gen[1109]),

			.O(gen[1202]),
			.E(gen[1204]),

			.SO(gen[1297]),
			.S(gen[1298]),
			.SE(gen[1299]),

			.SELF(gen[1203]),
			.cell_state(gen[1203])
		); 

/******************* CELL 1204 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1204 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1108]),
			.N(gen[1109]),
			.NE(gen[1110]),

			.O(gen[1203]),
			.E(gen[1205]),

			.SO(gen[1298]),
			.S(gen[1299]),
			.SE(gen[1300]),

			.SELF(gen[1204]),
			.cell_state(gen[1204])
		); 

/******************* CELL 1205 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1205 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1109]),
			.N(gen[1110]),
			.NE(gen[1111]),

			.O(gen[1204]),
			.E(gen[1206]),

			.SO(gen[1299]),
			.S(gen[1300]),
			.SE(gen[1301]),

			.SELF(gen[1205]),
			.cell_state(gen[1205])
		); 

/******************* CELL 1206 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1206 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1110]),
			.N(gen[1111]),
			.NE(gen[1112]),

			.O(gen[1205]),
			.E(gen[1207]),

			.SO(gen[1300]),
			.S(gen[1301]),
			.SE(gen[1302]),

			.SELF(gen[1206]),
			.cell_state(gen[1206])
		); 

/******************* CELL 1207 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1207 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1111]),
			.N(gen[1112]),
			.NE(gen[1113]),

			.O(gen[1206]),
			.E(gen[1208]),

			.SO(gen[1301]),
			.S(gen[1302]),
			.SE(gen[1303]),

			.SELF(gen[1207]),
			.cell_state(gen[1207])
		); 

/******************* CELL 1208 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1208 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1112]),
			.N(gen[1113]),
			.NE(gen[1114]),

			.O(gen[1207]),
			.E(gen[1209]),

			.SO(gen[1302]),
			.S(gen[1303]),
			.SE(gen[1304]),

			.SELF(gen[1208]),
			.cell_state(gen[1208])
		); 

/******************* CELL 1209 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1209 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1113]),
			.N(gen[1114]),
			.NE(gen[1115]),

			.O(gen[1208]),
			.E(gen[1210]),

			.SO(gen[1303]),
			.S(gen[1304]),
			.SE(gen[1305]),

			.SELF(gen[1209]),
			.cell_state(gen[1209])
		); 

/******************* CELL 1210 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1210 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1114]),
			.N(gen[1115]),
			.NE(gen[1116]),

			.O(gen[1209]),
			.E(gen[1211]),

			.SO(gen[1304]),
			.S(gen[1305]),
			.SE(gen[1306]),

			.SELF(gen[1210]),
			.cell_state(gen[1210])
		); 

/******************* CELL 1211 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1211 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1115]),
			.N(gen[1116]),
			.NE(gen[1117]),

			.O(gen[1210]),
			.E(gen[1212]),

			.SO(gen[1305]),
			.S(gen[1306]),
			.SE(gen[1307]),

			.SELF(gen[1211]),
			.cell_state(gen[1211])
		); 

/******************* CELL 1212 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1212 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1116]),
			.N(gen[1117]),
			.NE(gen[1118]),

			.O(gen[1211]),
			.E(gen[1213]),

			.SO(gen[1306]),
			.S(gen[1307]),
			.SE(gen[1308]),

			.SELF(gen[1212]),
			.cell_state(gen[1212])
		); 

/******************* CELL 1213 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1213 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1117]),
			.N(gen[1118]),
			.NE(gen[1119]),

			.O(gen[1212]),
			.E(gen[1214]),

			.SO(gen[1307]),
			.S(gen[1308]),
			.SE(gen[1309]),

			.SELF(gen[1213]),
			.cell_state(gen[1213])
		); 

/******************* CELL 1214 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1214 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1118]),
			.N(gen[1119]),
			.NE(gen[1120]),

			.O(gen[1213]),
			.E(gen[1215]),

			.SO(gen[1308]),
			.S(gen[1309]),
			.SE(gen[1310]),

			.SELF(gen[1214]),
			.cell_state(gen[1214])
		); 

/******************* CELL 1215 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1215 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1119]),
			.N(gen[1120]),
			.NE(gen[1121]),

			.O(gen[1214]),
			.E(gen[1216]),

			.SO(gen[1309]),
			.S(gen[1310]),
			.SE(gen[1311]),

			.SELF(gen[1215]),
			.cell_state(gen[1215])
		); 

/******************* CELL 1216 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1216 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1120]),
			.N(gen[1121]),
			.NE(gen[1122]),

			.O(gen[1215]),
			.E(gen[1217]),

			.SO(gen[1310]),
			.S(gen[1311]),
			.SE(gen[1312]),

			.SELF(gen[1216]),
			.cell_state(gen[1216])
		); 

/******************* CELL 1217 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1217 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1121]),
			.N(gen[1122]),
			.NE(gen[1123]),

			.O(gen[1216]),
			.E(gen[1218]),

			.SO(gen[1311]),
			.S(gen[1312]),
			.SE(gen[1313]),

			.SELF(gen[1217]),
			.cell_state(gen[1217])
		); 

/******************* CELL 1218 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1218 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1122]),
			.N(gen[1123]),
			.NE(gen[1124]),

			.O(gen[1217]),
			.E(gen[1219]),

			.SO(gen[1312]),
			.S(gen[1313]),
			.SE(gen[1314]),

			.SELF(gen[1218]),
			.cell_state(gen[1218])
		); 

/******************* CELL 1219 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1219 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1123]),
			.N(gen[1124]),
			.NE(gen[1125]),

			.O(gen[1218]),
			.E(gen[1220]),

			.SO(gen[1313]),
			.S(gen[1314]),
			.SE(gen[1315]),

			.SELF(gen[1219]),
			.cell_state(gen[1219])
		); 

/******************* CELL 1220 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1220 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1124]),
			.N(gen[1125]),
			.NE(gen[1126]),

			.O(gen[1219]),
			.E(gen[1221]),

			.SO(gen[1314]),
			.S(gen[1315]),
			.SE(gen[1316]),

			.SELF(gen[1220]),
			.cell_state(gen[1220])
		); 

/******************* CELL 1221 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1221 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1125]),
			.N(gen[1126]),
			.NE(gen[1127]),

			.O(gen[1220]),
			.E(gen[1222]),

			.SO(gen[1315]),
			.S(gen[1316]),
			.SE(gen[1317]),

			.SELF(gen[1221]),
			.cell_state(gen[1221])
		); 

/******************* CELL 1222 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1222 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1126]),
			.N(gen[1127]),
			.NE(gen[1128]),

			.O(gen[1221]),
			.E(gen[1223]),

			.SO(gen[1316]),
			.S(gen[1317]),
			.SE(gen[1318]),

			.SELF(gen[1222]),
			.cell_state(gen[1222])
		); 

/******************* CELL 1223 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1223 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1127]),
			.N(gen[1128]),
			.NE(gen[1129]),

			.O(gen[1222]),
			.E(gen[1224]),

			.SO(gen[1317]),
			.S(gen[1318]),
			.SE(gen[1319]),

			.SELF(gen[1223]),
			.cell_state(gen[1223])
		); 

/******************* CELL 1224 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1224 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1128]),
			.N(gen[1129]),
			.NE(gen[1130]),

			.O(gen[1223]),
			.E(gen[1225]),

			.SO(gen[1318]),
			.S(gen[1319]),
			.SE(gen[1320]),

			.SELF(gen[1224]),
			.cell_state(gen[1224])
		); 

/******************* CELL 1225 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1225 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1129]),
			.N(gen[1130]),
			.NE(gen[1131]),

			.O(gen[1224]),
			.E(gen[1226]),

			.SO(gen[1319]),
			.S(gen[1320]),
			.SE(gen[1321]),

			.SELF(gen[1225]),
			.cell_state(gen[1225])
		); 

/******************* CELL 1226 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1226 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1130]),
			.N(gen[1131]),
			.NE(gen[1132]),

			.O(gen[1225]),
			.E(gen[1227]),

			.SO(gen[1320]),
			.S(gen[1321]),
			.SE(gen[1322]),

			.SELF(gen[1226]),
			.cell_state(gen[1226])
		); 

/******************* CELL 1227 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1227 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1131]),
			.N(gen[1132]),
			.NE(gen[1133]),

			.O(gen[1226]),
			.E(gen[1228]),

			.SO(gen[1321]),
			.S(gen[1322]),
			.SE(gen[1323]),

			.SELF(gen[1227]),
			.cell_state(gen[1227])
		); 

/******************* CELL 1228 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1228 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1132]),
			.N(gen[1133]),
			.NE(gen[1134]),

			.O(gen[1227]),
			.E(gen[1229]),

			.SO(gen[1322]),
			.S(gen[1323]),
			.SE(gen[1324]),

			.SELF(gen[1228]),
			.cell_state(gen[1228])
		); 

/******************* CELL 1229 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1229 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1133]),
			.N(gen[1134]),
			.NE(gen[1135]),

			.O(gen[1228]),
			.E(gen[1230]),

			.SO(gen[1323]),
			.S(gen[1324]),
			.SE(gen[1325]),

			.SELF(gen[1229]),
			.cell_state(gen[1229])
		); 

/******************* CELL 1230 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1230 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1134]),
			.N(gen[1135]),
			.NE(gen[1136]),

			.O(gen[1229]),
			.E(gen[1231]),

			.SO(gen[1324]),
			.S(gen[1325]),
			.SE(gen[1326]),

			.SELF(gen[1230]),
			.cell_state(gen[1230])
		); 

/******************* CELL 1231 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1231 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1135]),
			.N(gen[1136]),
			.NE(gen[1137]),

			.O(gen[1230]),
			.E(gen[1232]),

			.SO(gen[1325]),
			.S(gen[1326]),
			.SE(gen[1327]),

			.SELF(gen[1231]),
			.cell_state(gen[1231])
		); 

/******************* CELL 1232 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1232 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1136]),
			.N(gen[1137]),
			.NE(gen[1138]),

			.O(gen[1231]),
			.E(gen[1233]),

			.SO(gen[1326]),
			.S(gen[1327]),
			.SE(gen[1328]),

			.SELF(gen[1232]),
			.cell_state(gen[1232])
		); 

/******************* CELL 1233 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1233 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1137]),
			.N(gen[1138]),
			.NE(gen[1139]),

			.O(gen[1232]),
			.E(gen[1234]),

			.SO(gen[1327]),
			.S(gen[1328]),
			.SE(gen[1329]),

			.SELF(gen[1233]),
			.cell_state(gen[1233])
		); 

/******************* CELL 1234 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1234 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1138]),
			.N(gen[1139]),
			.NE(gen[1138]),

			.O(gen[1233]),
			.E(gen[1233]),

			.SO(gen[1328]),
			.S(gen[1329]),
			.SE(gen[1328]),

			.SELF(gen[1234]),
			.cell_state(gen[1234])
		); 

/******************* CELL 1235 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1235 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1141]),
			.N(gen[1140]),
			.NE(gen[1141]),

			.O(gen[1236]),
			.E(gen[1236]),

			.SO(gen[1331]),
			.S(gen[1330]),
			.SE(gen[1331]),

			.SELF(gen[1235]),
			.cell_state(gen[1235])
		); 

/******************* CELL 1236 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1236 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1140]),
			.N(gen[1141]),
			.NE(gen[1142]),

			.O(gen[1235]),
			.E(gen[1237]),

			.SO(gen[1330]),
			.S(gen[1331]),
			.SE(gen[1332]),

			.SELF(gen[1236]),
			.cell_state(gen[1236])
		); 

/******************* CELL 1237 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1237 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1141]),
			.N(gen[1142]),
			.NE(gen[1143]),

			.O(gen[1236]),
			.E(gen[1238]),

			.SO(gen[1331]),
			.S(gen[1332]),
			.SE(gen[1333]),

			.SELF(gen[1237]),
			.cell_state(gen[1237])
		); 

/******************* CELL 1238 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1238 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1142]),
			.N(gen[1143]),
			.NE(gen[1144]),

			.O(gen[1237]),
			.E(gen[1239]),

			.SO(gen[1332]),
			.S(gen[1333]),
			.SE(gen[1334]),

			.SELF(gen[1238]),
			.cell_state(gen[1238])
		); 

/******************* CELL 1239 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1239 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1143]),
			.N(gen[1144]),
			.NE(gen[1145]),

			.O(gen[1238]),
			.E(gen[1240]),

			.SO(gen[1333]),
			.S(gen[1334]),
			.SE(gen[1335]),

			.SELF(gen[1239]),
			.cell_state(gen[1239])
		); 

/******************* CELL 1240 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1240 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1144]),
			.N(gen[1145]),
			.NE(gen[1146]),

			.O(gen[1239]),
			.E(gen[1241]),

			.SO(gen[1334]),
			.S(gen[1335]),
			.SE(gen[1336]),

			.SELF(gen[1240]),
			.cell_state(gen[1240])
		); 

/******************* CELL 1241 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1241 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1145]),
			.N(gen[1146]),
			.NE(gen[1147]),

			.O(gen[1240]),
			.E(gen[1242]),

			.SO(gen[1335]),
			.S(gen[1336]),
			.SE(gen[1337]),

			.SELF(gen[1241]),
			.cell_state(gen[1241])
		); 

/******************* CELL 1242 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1242 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1146]),
			.N(gen[1147]),
			.NE(gen[1148]),

			.O(gen[1241]),
			.E(gen[1243]),

			.SO(gen[1336]),
			.S(gen[1337]),
			.SE(gen[1338]),

			.SELF(gen[1242]),
			.cell_state(gen[1242])
		); 

/******************* CELL 1243 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1243 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1147]),
			.N(gen[1148]),
			.NE(gen[1149]),

			.O(gen[1242]),
			.E(gen[1244]),

			.SO(gen[1337]),
			.S(gen[1338]),
			.SE(gen[1339]),

			.SELF(gen[1243]),
			.cell_state(gen[1243])
		); 

/******************* CELL 1244 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1244 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1148]),
			.N(gen[1149]),
			.NE(gen[1150]),

			.O(gen[1243]),
			.E(gen[1245]),

			.SO(gen[1338]),
			.S(gen[1339]),
			.SE(gen[1340]),

			.SELF(gen[1244]),
			.cell_state(gen[1244])
		); 

/******************* CELL 1245 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1245 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1149]),
			.N(gen[1150]),
			.NE(gen[1151]),

			.O(gen[1244]),
			.E(gen[1246]),

			.SO(gen[1339]),
			.S(gen[1340]),
			.SE(gen[1341]),

			.SELF(gen[1245]),
			.cell_state(gen[1245])
		); 

/******************* CELL 1246 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1246 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1150]),
			.N(gen[1151]),
			.NE(gen[1152]),

			.O(gen[1245]),
			.E(gen[1247]),

			.SO(gen[1340]),
			.S(gen[1341]),
			.SE(gen[1342]),

			.SELF(gen[1246]),
			.cell_state(gen[1246])
		); 

/******************* CELL 1247 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1247 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1151]),
			.N(gen[1152]),
			.NE(gen[1153]),

			.O(gen[1246]),
			.E(gen[1248]),

			.SO(gen[1341]),
			.S(gen[1342]),
			.SE(gen[1343]),

			.SELF(gen[1247]),
			.cell_state(gen[1247])
		); 

/******************* CELL 1248 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1248 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1152]),
			.N(gen[1153]),
			.NE(gen[1154]),

			.O(gen[1247]),
			.E(gen[1249]),

			.SO(gen[1342]),
			.S(gen[1343]),
			.SE(gen[1344]),

			.SELF(gen[1248]),
			.cell_state(gen[1248])
		); 

/******************* CELL 1249 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1249 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1153]),
			.N(gen[1154]),
			.NE(gen[1155]),

			.O(gen[1248]),
			.E(gen[1250]),

			.SO(gen[1343]),
			.S(gen[1344]),
			.SE(gen[1345]),

			.SELF(gen[1249]),
			.cell_state(gen[1249])
		); 

/******************* CELL 1250 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1250 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1154]),
			.N(gen[1155]),
			.NE(gen[1156]),

			.O(gen[1249]),
			.E(gen[1251]),

			.SO(gen[1344]),
			.S(gen[1345]),
			.SE(gen[1346]),

			.SELF(gen[1250]),
			.cell_state(gen[1250])
		); 

/******************* CELL 1251 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1251 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1155]),
			.N(gen[1156]),
			.NE(gen[1157]),

			.O(gen[1250]),
			.E(gen[1252]),

			.SO(gen[1345]),
			.S(gen[1346]),
			.SE(gen[1347]),

			.SELF(gen[1251]),
			.cell_state(gen[1251])
		); 

/******************* CELL 1252 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1252 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1156]),
			.N(gen[1157]),
			.NE(gen[1158]),

			.O(gen[1251]),
			.E(gen[1253]),

			.SO(gen[1346]),
			.S(gen[1347]),
			.SE(gen[1348]),

			.SELF(gen[1252]),
			.cell_state(gen[1252])
		); 

/******************* CELL 1253 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1253 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1157]),
			.N(gen[1158]),
			.NE(gen[1159]),

			.O(gen[1252]),
			.E(gen[1254]),

			.SO(gen[1347]),
			.S(gen[1348]),
			.SE(gen[1349]),

			.SELF(gen[1253]),
			.cell_state(gen[1253])
		); 

/******************* CELL 1254 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1254 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1158]),
			.N(gen[1159]),
			.NE(gen[1160]),

			.O(gen[1253]),
			.E(gen[1255]),

			.SO(gen[1348]),
			.S(gen[1349]),
			.SE(gen[1350]),

			.SELF(gen[1254]),
			.cell_state(gen[1254])
		); 

/******************* CELL 1255 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1255 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1159]),
			.N(gen[1160]),
			.NE(gen[1161]),

			.O(gen[1254]),
			.E(gen[1256]),

			.SO(gen[1349]),
			.S(gen[1350]),
			.SE(gen[1351]),

			.SELF(gen[1255]),
			.cell_state(gen[1255])
		); 

/******************* CELL 1256 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1256 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1160]),
			.N(gen[1161]),
			.NE(gen[1162]),

			.O(gen[1255]),
			.E(gen[1257]),

			.SO(gen[1350]),
			.S(gen[1351]),
			.SE(gen[1352]),

			.SELF(gen[1256]),
			.cell_state(gen[1256])
		); 

/******************* CELL 1257 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1257 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1161]),
			.N(gen[1162]),
			.NE(gen[1163]),

			.O(gen[1256]),
			.E(gen[1258]),

			.SO(gen[1351]),
			.S(gen[1352]),
			.SE(gen[1353]),

			.SELF(gen[1257]),
			.cell_state(gen[1257])
		); 

/******************* CELL 1258 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1258 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1162]),
			.N(gen[1163]),
			.NE(gen[1164]),

			.O(gen[1257]),
			.E(gen[1259]),

			.SO(gen[1352]),
			.S(gen[1353]),
			.SE(gen[1354]),

			.SELF(gen[1258]),
			.cell_state(gen[1258])
		); 

/******************* CELL 1259 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1259 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1163]),
			.N(gen[1164]),
			.NE(gen[1165]),

			.O(gen[1258]),
			.E(gen[1260]),

			.SO(gen[1353]),
			.S(gen[1354]),
			.SE(gen[1355]),

			.SELF(gen[1259]),
			.cell_state(gen[1259])
		); 

/******************* CELL 1260 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1260 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1164]),
			.N(gen[1165]),
			.NE(gen[1166]),

			.O(gen[1259]),
			.E(gen[1261]),

			.SO(gen[1354]),
			.S(gen[1355]),
			.SE(gen[1356]),

			.SELF(gen[1260]),
			.cell_state(gen[1260])
		); 

/******************* CELL 1261 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1261 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1165]),
			.N(gen[1166]),
			.NE(gen[1167]),

			.O(gen[1260]),
			.E(gen[1262]),

			.SO(gen[1355]),
			.S(gen[1356]),
			.SE(gen[1357]),

			.SELF(gen[1261]),
			.cell_state(gen[1261])
		); 

/******************* CELL 1262 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1262 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1166]),
			.N(gen[1167]),
			.NE(gen[1168]),

			.O(gen[1261]),
			.E(gen[1263]),

			.SO(gen[1356]),
			.S(gen[1357]),
			.SE(gen[1358]),

			.SELF(gen[1262]),
			.cell_state(gen[1262])
		); 

/******************* CELL 1263 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1263 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1167]),
			.N(gen[1168]),
			.NE(gen[1169]),

			.O(gen[1262]),
			.E(gen[1264]),

			.SO(gen[1357]),
			.S(gen[1358]),
			.SE(gen[1359]),

			.SELF(gen[1263]),
			.cell_state(gen[1263])
		); 

/******************* CELL 1264 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1264 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1168]),
			.N(gen[1169]),
			.NE(gen[1170]),

			.O(gen[1263]),
			.E(gen[1265]),

			.SO(gen[1358]),
			.S(gen[1359]),
			.SE(gen[1360]),

			.SELF(gen[1264]),
			.cell_state(gen[1264])
		); 

/******************* CELL 1265 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1265 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1169]),
			.N(gen[1170]),
			.NE(gen[1171]),

			.O(gen[1264]),
			.E(gen[1266]),

			.SO(gen[1359]),
			.S(gen[1360]),
			.SE(gen[1361]),

			.SELF(gen[1265]),
			.cell_state(gen[1265])
		); 

/******************* CELL 1266 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1266 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1170]),
			.N(gen[1171]),
			.NE(gen[1172]),

			.O(gen[1265]),
			.E(gen[1267]),

			.SO(gen[1360]),
			.S(gen[1361]),
			.SE(gen[1362]),

			.SELF(gen[1266]),
			.cell_state(gen[1266])
		); 

/******************* CELL 1267 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1267 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1171]),
			.N(gen[1172]),
			.NE(gen[1173]),

			.O(gen[1266]),
			.E(gen[1268]),

			.SO(gen[1361]),
			.S(gen[1362]),
			.SE(gen[1363]),

			.SELF(gen[1267]),
			.cell_state(gen[1267])
		); 

/******************* CELL 1268 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1268 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1172]),
			.N(gen[1173]),
			.NE(gen[1174]),

			.O(gen[1267]),
			.E(gen[1269]),

			.SO(gen[1362]),
			.S(gen[1363]),
			.SE(gen[1364]),

			.SELF(gen[1268]),
			.cell_state(gen[1268])
		); 

/******************* CELL 1269 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1269 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1173]),
			.N(gen[1174]),
			.NE(gen[1175]),

			.O(gen[1268]),
			.E(gen[1270]),

			.SO(gen[1363]),
			.S(gen[1364]),
			.SE(gen[1365]),

			.SELF(gen[1269]),
			.cell_state(gen[1269])
		); 

/******************* CELL 1270 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1270 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1174]),
			.N(gen[1175]),
			.NE(gen[1176]),

			.O(gen[1269]),
			.E(gen[1271]),

			.SO(gen[1364]),
			.S(gen[1365]),
			.SE(gen[1366]),

			.SELF(gen[1270]),
			.cell_state(gen[1270])
		); 

/******************* CELL 1271 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1271 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1175]),
			.N(gen[1176]),
			.NE(gen[1177]),

			.O(gen[1270]),
			.E(gen[1272]),

			.SO(gen[1365]),
			.S(gen[1366]),
			.SE(gen[1367]),

			.SELF(gen[1271]),
			.cell_state(gen[1271])
		); 

/******************* CELL 1272 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1272 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1176]),
			.N(gen[1177]),
			.NE(gen[1178]),

			.O(gen[1271]),
			.E(gen[1273]),

			.SO(gen[1366]),
			.S(gen[1367]),
			.SE(gen[1368]),

			.SELF(gen[1272]),
			.cell_state(gen[1272])
		); 

/******************* CELL 1273 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1273 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1177]),
			.N(gen[1178]),
			.NE(gen[1179]),

			.O(gen[1272]),
			.E(gen[1274]),

			.SO(gen[1367]),
			.S(gen[1368]),
			.SE(gen[1369]),

			.SELF(gen[1273]),
			.cell_state(gen[1273])
		); 

/******************* CELL 1274 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1274 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1178]),
			.N(gen[1179]),
			.NE(gen[1180]),

			.O(gen[1273]),
			.E(gen[1275]),

			.SO(gen[1368]),
			.S(gen[1369]),
			.SE(gen[1370]),

			.SELF(gen[1274]),
			.cell_state(gen[1274])
		); 

/******************* CELL 1275 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1275 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1179]),
			.N(gen[1180]),
			.NE(gen[1181]),

			.O(gen[1274]),
			.E(gen[1276]),

			.SO(gen[1369]),
			.S(gen[1370]),
			.SE(gen[1371]),

			.SELF(gen[1275]),
			.cell_state(gen[1275])
		); 

/******************* CELL 1276 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1276 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1180]),
			.N(gen[1181]),
			.NE(gen[1182]),

			.O(gen[1275]),
			.E(gen[1277]),

			.SO(gen[1370]),
			.S(gen[1371]),
			.SE(gen[1372]),

			.SELF(gen[1276]),
			.cell_state(gen[1276])
		); 

/******************* CELL 1277 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1277 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1181]),
			.N(gen[1182]),
			.NE(gen[1183]),

			.O(gen[1276]),
			.E(gen[1278]),

			.SO(gen[1371]),
			.S(gen[1372]),
			.SE(gen[1373]),

			.SELF(gen[1277]),
			.cell_state(gen[1277])
		); 

/******************* CELL 1278 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1278 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1182]),
			.N(gen[1183]),
			.NE(gen[1184]),

			.O(gen[1277]),
			.E(gen[1279]),

			.SO(gen[1372]),
			.S(gen[1373]),
			.SE(gen[1374]),

			.SELF(gen[1278]),
			.cell_state(gen[1278])
		); 

/******************* CELL 1279 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1279 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1183]),
			.N(gen[1184]),
			.NE(gen[1185]),

			.O(gen[1278]),
			.E(gen[1280]),

			.SO(gen[1373]),
			.S(gen[1374]),
			.SE(gen[1375]),

			.SELF(gen[1279]),
			.cell_state(gen[1279])
		); 

/******************* CELL 1280 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1280 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1184]),
			.N(gen[1185]),
			.NE(gen[1186]),

			.O(gen[1279]),
			.E(gen[1281]),

			.SO(gen[1374]),
			.S(gen[1375]),
			.SE(gen[1376]),

			.SELF(gen[1280]),
			.cell_state(gen[1280])
		); 

/******************* CELL 1281 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1281 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1185]),
			.N(gen[1186]),
			.NE(gen[1187]),

			.O(gen[1280]),
			.E(gen[1282]),

			.SO(gen[1375]),
			.S(gen[1376]),
			.SE(gen[1377]),

			.SELF(gen[1281]),
			.cell_state(gen[1281])
		); 

/******************* CELL 1282 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1282 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1186]),
			.N(gen[1187]),
			.NE(gen[1188]),

			.O(gen[1281]),
			.E(gen[1283]),

			.SO(gen[1376]),
			.S(gen[1377]),
			.SE(gen[1378]),

			.SELF(gen[1282]),
			.cell_state(gen[1282])
		); 

/******************* CELL 1283 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1283 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1187]),
			.N(gen[1188]),
			.NE(gen[1189]),

			.O(gen[1282]),
			.E(gen[1284]),

			.SO(gen[1377]),
			.S(gen[1378]),
			.SE(gen[1379]),

			.SELF(gen[1283]),
			.cell_state(gen[1283])
		); 

/******************* CELL 1284 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1284 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1188]),
			.N(gen[1189]),
			.NE(gen[1190]),

			.O(gen[1283]),
			.E(gen[1285]),

			.SO(gen[1378]),
			.S(gen[1379]),
			.SE(gen[1380]),

			.SELF(gen[1284]),
			.cell_state(gen[1284])
		); 

/******************* CELL 1285 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1285 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1189]),
			.N(gen[1190]),
			.NE(gen[1191]),

			.O(gen[1284]),
			.E(gen[1286]),

			.SO(gen[1379]),
			.S(gen[1380]),
			.SE(gen[1381]),

			.SELF(gen[1285]),
			.cell_state(gen[1285])
		); 

/******************* CELL 1286 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1286 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1190]),
			.N(gen[1191]),
			.NE(gen[1192]),

			.O(gen[1285]),
			.E(gen[1287]),

			.SO(gen[1380]),
			.S(gen[1381]),
			.SE(gen[1382]),

			.SELF(gen[1286]),
			.cell_state(gen[1286])
		); 

/******************* CELL 1287 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1287 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1191]),
			.N(gen[1192]),
			.NE(gen[1193]),

			.O(gen[1286]),
			.E(gen[1288]),

			.SO(gen[1381]),
			.S(gen[1382]),
			.SE(gen[1383]),

			.SELF(gen[1287]),
			.cell_state(gen[1287])
		); 

/******************* CELL 1288 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1288 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1192]),
			.N(gen[1193]),
			.NE(gen[1194]),

			.O(gen[1287]),
			.E(gen[1289]),

			.SO(gen[1382]),
			.S(gen[1383]),
			.SE(gen[1384]),

			.SELF(gen[1288]),
			.cell_state(gen[1288])
		); 

/******************* CELL 1289 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1289 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1193]),
			.N(gen[1194]),
			.NE(gen[1195]),

			.O(gen[1288]),
			.E(gen[1290]),

			.SO(gen[1383]),
			.S(gen[1384]),
			.SE(gen[1385]),

			.SELF(gen[1289]),
			.cell_state(gen[1289])
		); 

/******************* CELL 1290 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1290 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1194]),
			.N(gen[1195]),
			.NE(gen[1196]),

			.O(gen[1289]),
			.E(gen[1291]),

			.SO(gen[1384]),
			.S(gen[1385]),
			.SE(gen[1386]),

			.SELF(gen[1290]),
			.cell_state(gen[1290])
		); 

/******************* CELL 1291 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1291 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1195]),
			.N(gen[1196]),
			.NE(gen[1197]),

			.O(gen[1290]),
			.E(gen[1292]),

			.SO(gen[1385]),
			.S(gen[1386]),
			.SE(gen[1387]),

			.SELF(gen[1291]),
			.cell_state(gen[1291])
		); 

/******************* CELL 1292 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1292 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1196]),
			.N(gen[1197]),
			.NE(gen[1198]),

			.O(gen[1291]),
			.E(gen[1293]),

			.SO(gen[1386]),
			.S(gen[1387]),
			.SE(gen[1388]),

			.SELF(gen[1292]),
			.cell_state(gen[1292])
		); 

/******************* CELL 1293 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1293 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1197]),
			.N(gen[1198]),
			.NE(gen[1199]),

			.O(gen[1292]),
			.E(gen[1294]),

			.SO(gen[1387]),
			.S(gen[1388]),
			.SE(gen[1389]),

			.SELF(gen[1293]),
			.cell_state(gen[1293])
		); 

/******************* CELL 1294 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1294 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1198]),
			.N(gen[1199]),
			.NE(gen[1200]),

			.O(gen[1293]),
			.E(gen[1295]),

			.SO(gen[1388]),
			.S(gen[1389]),
			.SE(gen[1390]),

			.SELF(gen[1294]),
			.cell_state(gen[1294])
		); 

/******************* CELL 1295 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1295 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1199]),
			.N(gen[1200]),
			.NE(gen[1201]),

			.O(gen[1294]),
			.E(gen[1296]),

			.SO(gen[1389]),
			.S(gen[1390]),
			.SE(gen[1391]),

			.SELF(gen[1295]),
			.cell_state(gen[1295])
		); 

/******************* CELL 1296 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1296 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1200]),
			.N(gen[1201]),
			.NE(gen[1202]),

			.O(gen[1295]),
			.E(gen[1297]),

			.SO(gen[1390]),
			.S(gen[1391]),
			.SE(gen[1392]),

			.SELF(gen[1296]),
			.cell_state(gen[1296])
		); 

/******************* CELL 1297 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1297 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1201]),
			.N(gen[1202]),
			.NE(gen[1203]),

			.O(gen[1296]),
			.E(gen[1298]),

			.SO(gen[1391]),
			.S(gen[1392]),
			.SE(gen[1393]),

			.SELF(gen[1297]),
			.cell_state(gen[1297])
		); 

/******************* CELL 1298 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1298 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1202]),
			.N(gen[1203]),
			.NE(gen[1204]),

			.O(gen[1297]),
			.E(gen[1299]),

			.SO(gen[1392]),
			.S(gen[1393]),
			.SE(gen[1394]),

			.SELF(gen[1298]),
			.cell_state(gen[1298])
		); 

/******************* CELL 1299 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1299 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1203]),
			.N(gen[1204]),
			.NE(gen[1205]),

			.O(gen[1298]),
			.E(gen[1300]),

			.SO(gen[1393]),
			.S(gen[1394]),
			.SE(gen[1395]),

			.SELF(gen[1299]),
			.cell_state(gen[1299])
		); 

/******************* CELL 1300 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1300 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1204]),
			.N(gen[1205]),
			.NE(gen[1206]),

			.O(gen[1299]),
			.E(gen[1301]),

			.SO(gen[1394]),
			.S(gen[1395]),
			.SE(gen[1396]),

			.SELF(gen[1300]),
			.cell_state(gen[1300])
		); 

/******************* CELL 1301 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1301 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1205]),
			.N(gen[1206]),
			.NE(gen[1207]),

			.O(gen[1300]),
			.E(gen[1302]),

			.SO(gen[1395]),
			.S(gen[1396]),
			.SE(gen[1397]),

			.SELF(gen[1301]),
			.cell_state(gen[1301])
		); 

/******************* CELL 1302 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1302 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1206]),
			.N(gen[1207]),
			.NE(gen[1208]),

			.O(gen[1301]),
			.E(gen[1303]),

			.SO(gen[1396]),
			.S(gen[1397]),
			.SE(gen[1398]),

			.SELF(gen[1302]),
			.cell_state(gen[1302])
		); 

/******************* CELL 1303 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1303 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1207]),
			.N(gen[1208]),
			.NE(gen[1209]),

			.O(gen[1302]),
			.E(gen[1304]),

			.SO(gen[1397]),
			.S(gen[1398]),
			.SE(gen[1399]),

			.SELF(gen[1303]),
			.cell_state(gen[1303])
		); 

/******************* CELL 1304 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1304 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1208]),
			.N(gen[1209]),
			.NE(gen[1210]),

			.O(gen[1303]),
			.E(gen[1305]),

			.SO(gen[1398]),
			.S(gen[1399]),
			.SE(gen[1400]),

			.SELF(gen[1304]),
			.cell_state(gen[1304])
		); 

/******************* CELL 1305 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1305 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1209]),
			.N(gen[1210]),
			.NE(gen[1211]),

			.O(gen[1304]),
			.E(gen[1306]),

			.SO(gen[1399]),
			.S(gen[1400]),
			.SE(gen[1401]),

			.SELF(gen[1305]),
			.cell_state(gen[1305])
		); 

/******************* CELL 1306 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1306 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1210]),
			.N(gen[1211]),
			.NE(gen[1212]),

			.O(gen[1305]),
			.E(gen[1307]),

			.SO(gen[1400]),
			.S(gen[1401]),
			.SE(gen[1402]),

			.SELF(gen[1306]),
			.cell_state(gen[1306])
		); 

/******************* CELL 1307 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1307 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1211]),
			.N(gen[1212]),
			.NE(gen[1213]),

			.O(gen[1306]),
			.E(gen[1308]),

			.SO(gen[1401]),
			.S(gen[1402]),
			.SE(gen[1403]),

			.SELF(gen[1307]),
			.cell_state(gen[1307])
		); 

/******************* CELL 1308 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1308 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1212]),
			.N(gen[1213]),
			.NE(gen[1214]),

			.O(gen[1307]),
			.E(gen[1309]),

			.SO(gen[1402]),
			.S(gen[1403]),
			.SE(gen[1404]),

			.SELF(gen[1308]),
			.cell_state(gen[1308])
		); 

/******************* CELL 1309 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1309 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1213]),
			.N(gen[1214]),
			.NE(gen[1215]),

			.O(gen[1308]),
			.E(gen[1310]),

			.SO(gen[1403]),
			.S(gen[1404]),
			.SE(gen[1405]),

			.SELF(gen[1309]),
			.cell_state(gen[1309])
		); 

/******************* CELL 1310 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1310 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1214]),
			.N(gen[1215]),
			.NE(gen[1216]),

			.O(gen[1309]),
			.E(gen[1311]),

			.SO(gen[1404]),
			.S(gen[1405]),
			.SE(gen[1406]),

			.SELF(gen[1310]),
			.cell_state(gen[1310])
		); 

/******************* CELL 1311 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1311 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1215]),
			.N(gen[1216]),
			.NE(gen[1217]),

			.O(gen[1310]),
			.E(gen[1312]),

			.SO(gen[1405]),
			.S(gen[1406]),
			.SE(gen[1407]),

			.SELF(gen[1311]),
			.cell_state(gen[1311])
		); 

/******************* CELL 1312 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1312 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1216]),
			.N(gen[1217]),
			.NE(gen[1218]),

			.O(gen[1311]),
			.E(gen[1313]),

			.SO(gen[1406]),
			.S(gen[1407]),
			.SE(gen[1408]),

			.SELF(gen[1312]),
			.cell_state(gen[1312])
		); 

/******************* CELL 1313 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1313 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1217]),
			.N(gen[1218]),
			.NE(gen[1219]),

			.O(gen[1312]),
			.E(gen[1314]),

			.SO(gen[1407]),
			.S(gen[1408]),
			.SE(gen[1409]),

			.SELF(gen[1313]),
			.cell_state(gen[1313])
		); 

/******************* CELL 1314 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1314 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1218]),
			.N(gen[1219]),
			.NE(gen[1220]),

			.O(gen[1313]),
			.E(gen[1315]),

			.SO(gen[1408]),
			.S(gen[1409]),
			.SE(gen[1410]),

			.SELF(gen[1314]),
			.cell_state(gen[1314])
		); 

/******************* CELL 1315 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1315 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1219]),
			.N(gen[1220]),
			.NE(gen[1221]),

			.O(gen[1314]),
			.E(gen[1316]),

			.SO(gen[1409]),
			.S(gen[1410]),
			.SE(gen[1411]),

			.SELF(gen[1315]),
			.cell_state(gen[1315])
		); 

/******************* CELL 1316 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1316 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1220]),
			.N(gen[1221]),
			.NE(gen[1222]),

			.O(gen[1315]),
			.E(gen[1317]),

			.SO(gen[1410]),
			.S(gen[1411]),
			.SE(gen[1412]),

			.SELF(gen[1316]),
			.cell_state(gen[1316])
		); 

/******************* CELL 1317 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1317 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1221]),
			.N(gen[1222]),
			.NE(gen[1223]),

			.O(gen[1316]),
			.E(gen[1318]),

			.SO(gen[1411]),
			.S(gen[1412]),
			.SE(gen[1413]),

			.SELF(gen[1317]),
			.cell_state(gen[1317])
		); 

/******************* CELL 1318 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1318 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1222]),
			.N(gen[1223]),
			.NE(gen[1224]),

			.O(gen[1317]),
			.E(gen[1319]),

			.SO(gen[1412]),
			.S(gen[1413]),
			.SE(gen[1414]),

			.SELF(gen[1318]),
			.cell_state(gen[1318])
		); 

/******************* CELL 1319 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1319 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1223]),
			.N(gen[1224]),
			.NE(gen[1225]),

			.O(gen[1318]),
			.E(gen[1320]),

			.SO(gen[1413]),
			.S(gen[1414]),
			.SE(gen[1415]),

			.SELF(gen[1319]),
			.cell_state(gen[1319])
		); 

/******************* CELL 1320 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1320 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1224]),
			.N(gen[1225]),
			.NE(gen[1226]),

			.O(gen[1319]),
			.E(gen[1321]),

			.SO(gen[1414]),
			.S(gen[1415]),
			.SE(gen[1416]),

			.SELF(gen[1320]),
			.cell_state(gen[1320])
		); 

/******************* CELL 1321 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1321 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1225]),
			.N(gen[1226]),
			.NE(gen[1227]),

			.O(gen[1320]),
			.E(gen[1322]),

			.SO(gen[1415]),
			.S(gen[1416]),
			.SE(gen[1417]),

			.SELF(gen[1321]),
			.cell_state(gen[1321])
		); 

/******************* CELL 1322 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1322 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1226]),
			.N(gen[1227]),
			.NE(gen[1228]),

			.O(gen[1321]),
			.E(gen[1323]),

			.SO(gen[1416]),
			.S(gen[1417]),
			.SE(gen[1418]),

			.SELF(gen[1322]),
			.cell_state(gen[1322])
		); 

/******************* CELL 1323 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1323 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1227]),
			.N(gen[1228]),
			.NE(gen[1229]),

			.O(gen[1322]),
			.E(gen[1324]),

			.SO(gen[1417]),
			.S(gen[1418]),
			.SE(gen[1419]),

			.SELF(gen[1323]),
			.cell_state(gen[1323])
		); 

/******************* CELL 1324 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1324 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1228]),
			.N(gen[1229]),
			.NE(gen[1230]),

			.O(gen[1323]),
			.E(gen[1325]),

			.SO(gen[1418]),
			.S(gen[1419]),
			.SE(gen[1420]),

			.SELF(gen[1324]),
			.cell_state(gen[1324])
		); 

/******************* CELL 1325 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1325 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1229]),
			.N(gen[1230]),
			.NE(gen[1231]),

			.O(gen[1324]),
			.E(gen[1326]),

			.SO(gen[1419]),
			.S(gen[1420]),
			.SE(gen[1421]),

			.SELF(gen[1325]),
			.cell_state(gen[1325])
		); 

/******************* CELL 1326 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1326 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1230]),
			.N(gen[1231]),
			.NE(gen[1232]),

			.O(gen[1325]),
			.E(gen[1327]),

			.SO(gen[1420]),
			.S(gen[1421]),
			.SE(gen[1422]),

			.SELF(gen[1326]),
			.cell_state(gen[1326])
		); 

/******************* CELL 1327 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1327 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1231]),
			.N(gen[1232]),
			.NE(gen[1233]),

			.O(gen[1326]),
			.E(gen[1328]),

			.SO(gen[1421]),
			.S(gen[1422]),
			.SE(gen[1423]),

			.SELF(gen[1327]),
			.cell_state(gen[1327])
		); 

/******************* CELL 1328 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1328 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1232]),
			.N(gen[1233]),
			.NE(gen[1234]),

			.O(gen[1327]),
			.E(gen[1329]),

			.SO(gen[1422]),
			.S(gen[1423]),
			.SE(gen[1424]),

			.SELF(gen[1328]),
			.cell_state(gen[1328])
		); 

/******************* CELL 1329 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1329 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1233]),
			.N(gen[1234]),
			.NE(gen[1233]),

			.O(gen[1328]),
			.E(gen[1328]),

			.SO(gen[1423]),
			.S(gen[1424]),
			.SE(gen[1423]),

			.SELF(gen[1329]),
			.cell_state(gen[1329])
		); 

/******************* CELL 1330 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1330 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1236]),
			.N(gen[1235]),
			.NE(gen[1236]),

			.O(gen[1331]),
			.E(gen[1331]),

			.SO(gen[1426]),
			.S(gen[1425]),
			.SE(gen[1426]),

			.SELF(gen[1330]),
			.cell_state(gen[1330])
		); 

/******************* CELL 1331 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1331 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1235]),
			.N(gen[1236]),
			.NE(gen[1237]),

			.O(gen[1330]),
			.E(gen[1332]),

			.SO(gen[1425]),
			.S(gen[1426]),
			.SE(gen[1427]),

			.SELF(gen[1331]),
			.cell_state(gen[1331])
		); 

/******************* CELL 1332 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1332 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1236]),
			.N(gen[1237]),
			.NE(gen[1238]),

			.O(gen[1331]),
			.E(gen[1333]),

			.SO(gen[1426]),
			.S(gen[1427]),
			.SE(gen[1428]),

			.SELF(gen[1332]),
			.cell_state(gen[1332])
		); 

/******************* CELL 1333 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1333 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1237]),
			.N(gen[1238]),
			.NE(gen[1239]),

			.O(gen[1332]),
			.E(gen[1334]),

			.SO(gen[1427]),
			.S(gen[1428]),
			.SE(gen[1429]),

			.SELF(gen[1333]),
			.cell_state(gen[1333])
		); 

/******************* CELL 1334 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1334 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1238]),
			.N(gen[1239]),
			.NE(gen[1240]),

			.O(gen[1333]),
			.E(gen[1335]),

			.SO(gen[1428]),
			.S(gen[1429]),
			.SE(gen[1430]),

			.SELF(gen[1334]),
			.cell_state(gen[1334])
		); 

/******************* CELL 1335 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1335 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1239]),
			.N(gen[1240]),
			.NE(gen[1241]),

			.O(gen[1334]),
			.E(gen[1336]),

			.SO(gen[1429]),
			.S(gen[1430]),
			.SE(gen[1431]),

			.SELF(gen[1335]),
			.cell_state(gen[1335])
		); 

/******************* CELL 1336 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1336 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1240]),
			.N(gen[1241]),
			.NE(gen[1242]),

			.O(gen[1335]),
			.E(gen[1337]),

			.SO(gen[1430]),
			.S(gen[1431]),
			.SE(gen[1432]),

			.SELF(gen[1336]),
			.cell_state(gen[1336])
		); 

/******************* CELL 1337 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1337 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1241]),
			.N(gen[1242]),
			.NE(gen[1243]),

			.O(gen[1336]),
			.E(gen[1338]),

			.SO(gen[1431]),
			.S(gen[1432]),
			.SE(gen[1433]),

			.SELF(gen[1337]),
			.cell_state(gen[1337])
		); 

/******************* CELL 1338 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1338 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1242]),
			.N(gen[1243]),
			.NE(gen[1244]),

			.O(gen[1337]),
			.E(gen[1339]),

			.SO(gen[1432]),
			.S(gen[1433]),
			.SE(gen[1434]),

			.SELF(gen[1338]),
			.cell_state(gen[1338])
		); 

/******************* CELL 1339 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1339 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1243]),
			.N(gen[1244]),
			.NE(gen[1245]),

			.O(gen[1338]),
			.E(gen[1340]),

			.SO(gen[1433]),
			.S(gen[1434]),
			.SE(gen[1435]),

			.SELF(gen[1339]),
			.cell_state(gen[1339])
		); 

/******************* CELL 1340 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1340 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1244]),
			.N(gen[1245]),
			.NE(gen[1246]),

			.O(gen[1339]),
			.E(gen[1341]),

			.SO(gen[1434]),
			.S(gen[1435]),
			.SE(gen[1436]),

			.SELF(gen[1340]),
			.cell_state(gen[1340])
		); 

/******************* CELL 1341 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1341 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1245]),
			.N(gen[1246]),
			.NE(gen[1247]),

			.O(gen[1340]),
			.E(gen[1342]),

			.SO(gen[1435]),
			.S(gen[1436]),
			.SE(gen[1437]),

			.SELF(gen[1341]),
			.cell_state(gen[1341])
		); 

/******************* CELL 1342 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1342 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1246]),
			.N(gen[1247]),
			.NE(gen[1248]),

			.O(gen[1341]),
			.E(gen[1343]),

			.SO(gen[1436]),
			.S(gen[1437]),
			.SE(gen[1438]),

			.SELF(gen[1342]),
			.cell_state(gen[1342])
		); 

/******************* CELL 1343 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1343 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1247]),
			.N(gen[1248]),
			.NE(gen[1249]),

			.O(gen[1342]),
			.E(gen[1344]),

			.SO(gen[1437]),
			.S(gen[1438]),
			.SE(gen[1439]),

			.SELF(gen[1343]),
			.cell_state(gen[1343])
		); 

/******************* CELL 1344 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1344 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1248]),
			.N(gen[1249]),
			.NE(gen[1250]),

			.O(gen[1343]),
			.E(gen[1345]),

			.SO(gen[1438]),
			.S(gen[1439]),
			.SE(gen[1440]),

			.SELF(gen[1344]),
			.cell_state(gen[1344])
		); 

/******************* CELL 1345 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1345 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1249]),
			.N(gen[1250]),
			.NE(gen[1251]),

			.O(gen[1344]),
			.E(gen[1346]),

			.SO(gen[1439]),
			.S(gen[1440]),
			.SE(gen[1441]),

			.SELF(gen[1345]),
			.cell_state(gen[1345])
		); 

/******************* CELL 1346 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1346 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1250]),
			.N(gen[1251]),
			.NE(gen[1252]),

			.O(gen[1345]),
			.E(gen[1347]),

			.SO(gen[1440]),
			.S(gen[1441]),
			.SE(gen[1442]),

			.SELF(gen[1346]),
			.cell_state(gen[1346])
		); 

/******************* CELL 1347 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1347 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1251]),
			.N(gen[1252]),
			.NE(gen[1253]),

			.O(gen[1346]),
			.E(gen[1348]),

			.SO(gen[1441]),
			.S(gen[1442]),
			.SE(gen[1443]),

			.SELF(gen[1347]),
			.cell_state(gen[1347])
		); 

/******************* CELL 1348 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1348 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1252]),
			.N(gen[1253]),
			.NE(gen[1254]),

			.O(gen[1347]),
			.E(gen[1349]),

			.SO(gen[1442]),
			.S(gen[1443]),
			.SE(gen[1444]),

			.SELF(gen[1348]),
			.cell_state(gen[1348])
		); 

/******************* CELL 1349 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1349 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1253]),
			.N(gen[1254]),
			.NE(gen[1255]),

			.O(gen[1348]),
			.E(gen[1350]),

			.SO(gen[1443]),
			.S(gen[1444]),
			.SE(gen[1445]),

			.SELF(gen[1349]),
			.cell_state(gen[1349])
		); 

/******************* CELL 1350 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1350 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1254]),
			.N(gen[1255]),
			.NE(gen[1256]),

			.O(gen[1349]),
			.E(gen[1351]),

			.SO(gen[1444]),
			.S(gen[1445]),
			.SE(gen[1446]),

			.SELF(gen[1350]),
			.cell_state(gen[1350])
		); 

/******************* CELL 1351 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1351 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1255]),
			.N(gen[1256]),
			.NE(gen[1257]),

			.O(gen[1350]),
			.E(gen[1352]),

			.SO(gen[1445]),
			.S(gen[1446]),
			.SE(gen[1447]),

			.SELF(gen[1351]),
			.cell_state(gen[1351])
		); 

/******************* CELL 1352 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1352 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1256]),
			.N(gen[1257]),
			.NE(gen[1258]),

			.O(gen[1351]),
			.E(gen[1353]),

			.SO(gen[1446]),
			.S(gen[1447]),
			.SE(gen[1448]),

			.SELF(gen[1352]),
			.cell_state(gen[1352])
		); 

/******************* CELL 1353 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1353 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1257]),
			.N(gen[1258]),
			.NE(gen[1259]),

			.O(gen[1352]),
			.E(gen[1354]),

			.SO(gen[1447]),
			.S(gen[1448]),
			.SE(gen[1449]),

			.SELF(gen[1353]),
			.cell_state(gen[1353])
		); 

/******************* CELL 1354 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1354 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1258]),
			.N(gen[1259]),
			.NE(gen[1260]),

			.O(gen[1353]),
			.E(gen[1355]),

			.SO(gen[1448]),
			.S(gen[1449]),
			.SE(gen[1450]),

			.SELF(gen[1354]),
			.cell_state(gen[1354])
		); 

/******************* CELL 1355 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1355 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1259]),
			.N(gen[1260]),
			.NE(gen[1261]),

			.O(gen[1354]),
			.E(gen[1356]),

			.SO(gen[1449]),
			.S(gen[1450]),
			.SE(gen[1451]),

			.SELF(gen[1355]),
			.cell_state(gen[1355])
		); 

/******************* CELL 1356 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1356 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1260]),
			.N(gen[1261]),
			.NE(gen[1262]),

			.O(gen[1355]),
			.E(gen[1357]),

			.SO(gen[1450]),
			.S(gen[1451]),
			.SE(gen[1452]),

			.SELF(gen[1356]),
			.cell_state(gen[1356])
		); 

/******************* CELL 1357 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1357 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1261]),
			.N(gen[1262]),
			.NE(gen[1263]),

			.O(gen[1356]),
			.E(gen[1358]),

			.SO(gen[1451]),
			.S(gen[1452]),
			.SE(gen[1453]),

			.SELF(gen[1357]),
			.cell_state(gen[1357])
		); 

/******************* CELL 1358 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1358 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1262]),
			.N(gen[1263]),
			.NE(gen[1264]),

			.O(gen[1357]),
			.E(gen[1359]),

			.SO(gen[1452]),
			.S(gen[1453]),
			.SE(gen[1454]),

			.SELF(gen[1358]),
			.cell_state(gen[1358])
		); 

/******************* CELL 1359 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1359 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1263]),
			.N(gen[1264]),
			.NE(gen[1265]),

			.O(gen[1358]),
			.E(gen[1360]),

			.SO(gen[1453]),
			.S(gen[1454]),
			.SE(gen[1455]),

			.SELF(gen[1359]),
			.cell_state(gen[1359])
		); 

/******************* CELL 1360 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1360 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1264]),
			.N(gen[1265]),
			.NE(gen[1266]),

			.O(gen[1359]),
			.E(gen[1361]),

			.SO(gen[1454]),
			.S(gen[1455]),
			.SE(gen[1456]),

			.SELF(gen[1360]),
			.cell_state(gen[1360])
		); 

/******************* CELL 1361 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1361 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1265]),
			.N(gen[1266]),
			.NE(gen[1267]),

			.O(gen[1360]),
			.E(gen[1362]),

			.SO(gen[1455]),
			.S(gen[1456]),
			.SE(gen[1457]),

			.SELF(gen[1361]),
			.cell_state(gen[1361])
		); 

/******************* CELL 1362 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1362 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1266]),
			.N(gen[1267]),
			.NE(gen[1268]),

			.O(gen[1361]),
			.E(gen[1363]),

			.SO(gen[1456]),
			.S(gen[1457]),
			.SE(gen[1458]),

			.SELF(gen[1362]),
			.cell_state(gen[1362])
		); 

/******************* CELL 1363 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1363 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1267]),
			.N(gen[1268]),
			.NE(gen[1269]),

			.O(gen[1362]),
			.E(gen[1364]),

			.SO(gen[1457]),
			.S(gen[1458]),
			.SE(gen[1459]),

			.SELF(gen[1363]),
			.cell_state(gen[1363])
		); 

/******************* CELL 1364 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1364 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1268]),
			.N(gen[1269]),
			.NE(gen[1270]),

			.O(gen[1363]),
			.E(gen[1365]),

			.SO(gen[1458]),
			.S(gen[1459]),
			.SE(gen[1460]),

			.SELF(gen[1364]),
			.cell_state(gen[1364])
		); 

/******************* CELL 1365 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1365 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1269]),
			.N(gen[1270]),
			.NE(gen[1271]),

			.O(gen[1364]),
			.E(gen[1366]),

			.SO(gen[1459]),
			.S(gen[1460]),
			.SE(gen[1461]),

			.SELF(gen[1365]),
			.cell_state(gen[1365])
		); 

/******************* CELL 1366 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1366 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1270]),
			.N(gen[1271]),
			.NE(gen[1272]),

			.O(gen[1365]),
			.E(gen[1367]),

			.SO(gen[1460]),
			.S(gen[1461]),
			.SE(gen[1462]),

			.SELF(gen[1366]),
			.cell_state(gen[1366])
		); 

/******************* CELL 1367 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1367 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1271]),
			.N(gen[1272]),
			.NE(gen[1273]),

			.O(gen[1366]),
			.E(gen[1368]),

			.SO(gen[1461]),
			.S(gen[1462]),
			.SE(gen[1463]),

			.SELF(gen[1367]),
			.cell_state(gen[1367])
		); 

/******************* CELL 1368 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1368 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1272]),
			.N(gen[1273]),
			.NE(gen[1274]),

			.O(gen[1367]),
			.E(gen[1369]),

			.SO(gen[1462]),
			.S(gen[1463]),
			.SE(gen[1464]),

			.SELF(gen[1368]),
			.cell_state(gen[1368])
		); 

/******************* CELL 1369 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1369 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1273]),
			.N(gen[1274]),
			.NE(gen[1275]),

			.O(gen[1368]),
			.E(gen[1370]),

			.SO(gen[1463]),
			.S(gen[1464]),
			.SE(gen[1465]),

			.SELF(gen[1369]),
			.cell_state(gen[1369])
		); 

/******************* CELL 1370 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1370 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1274]),
			.N(gen[1275]),
			.NE(gen[1276]),

			.O(gen[1369]),
			.E(gen[1371]),

			.SO(gen[1464]),
			.S(gen[1465]),
			.SE(gen[1466]),

			.SELF(gen[1370]),
			.cell_state(gen[1370])
		); 

/******************* CELL 1371 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1371 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1275]),
			.N(gen[1276]),
			.NE(gen[1277]),

			.O(gen[1370]),
			.E(gen[1372]),

			.SO(gen[1465]),
			.S(gen[1466]),
			.SE(gen[1467]),

			.SELF(gen[1371]),
			.cell_state(gen[1371])
		); 

/******************* CELL 1372 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1372 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1276]),
			.N(gen[1277]),
			.NE(gen[1278]),

			.O(gen[1371]),
			.E(gen[1373]),

			.SO(gen[1466]),
			.S(gen[1467]),
			.SE(gen[1468]),

			.SELF(gen[1372]),
			.cell_state(gen[1372])
		); 

/******************* CELL 1373 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1373 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1277]),
			.N(gen[1278]),
			.NE(gen[1279]),

			.O(gen[1372]),
			.E(gen[1374]),

			.SO(gen[1467]),
			.S(gen[1468]),
			.SE(gen[1469]),

			.SELF(gen[1373]),
			.cell_state(gen[1373])
		); 

/******************* CELL 1374 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1374 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1278]),
			.N(gen[1279]),
			.NE(gen[1280]),

			.O(gen[1373]),
			.E(gen[1375]),

			.SO(gen[1468]),
			.S(gen[1469]),
			.SE(gen[1470]),

			.SELF(gen[1374]),
			.cell_state(gen[1374])
		); 

/******************* CELL 1375 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1375 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1279]),
			.N(gen[1280]),
			.NE(gen[1281]),

			.O(gen[1374]),
			.E(gen[1376]),

			.SO(gen[1469]),
			.S(gen[1470]),
			.SE(gen[1471]),

			.SELF(gen[1375]),
			.cell_state(gen[1375])
		); 

/******************* CELL 1376 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1376 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1280]),
			.N(gen[1281]),
			.NE(gen[1282]),

			.O(gen[1375]),
			.E(gen[1377]),

			.SO(gen[1470]),
			.S(gen[1471]),
			.SE(gen[1472]),

			.SELF(gen[1376]),
			.cell_state(gen[1376])
		); 

/******************* CELL 1377 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1377 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1281]),
			.N(gen[1282]),
			.NE(gen[1283]),

			.O(gen[1376]),
			.E(gen[1378]),

			.SO(gen[1471]),
			.S(gen[1472]),
			.SE(gen[1473]),

			.SELF(gen[1377]),
			.cell_state(gen[1377])
		); 

/******************* CELL 1378 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1378 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1282]),
			.N(gen[1283]),
			.NE(gen[1284]),

			.O(gen[1377]),
			.E(gen[1379]),

			.SO(gen[1472]),
			.S(gen[1473]),
			.SE(gen[1474]),

			.SELF(gen[1378]),
			.cell_state(gen[1378])
		); 

/******************* CELL 1379 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1379 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1283]),
			.N(gen[1284]),
			.NE(gen[1285]),

			.O(gen[1378]),
			.E(gen[1380]),

			.SO(gen[1473]),
			.S(gen[1474]),
			.SE(gen[1475]),

			.SELF(gen[1379]),
			.cell_state(gen[1379])
		); 

/******************* CELL 1380 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1380 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1284]),
			.N(gen[1285]),
			.NE(gen[1286]),

			.O(gen[1379]),
			.E(gen[1381]),

			.SO(gen[1474]),
			.S(gen[1475]),
			.SE(gen[1476]),

			.SELF(gen[1380]),
			.cell_state(gen[1380])
		); 

/******************* CELL 1381 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1381 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1285]),
			.N(gen[1286]),
			.NE(gen[1287]),

			.O(gen[1380]),
			.E(gen[1382]),

			.SO(gen[1475]),
			.S(gen[1476]),
			.SE(gen[1477]),

			.SELF(gen[1381]),
			.cell_state(gen[1381])
		); 

/******************* CELL 1382 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1382 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1286]),
			.N(gen[1287]),
			.NE(gen[1288]),

			.O(gen[1381]),
			.E(gen[1383]),

			.SO(gen[1476]),
			.S(gen[1477]),
			.SE(gen[1478]),

			.SELF(gen[1382]),
			.cell_state(gen[1382])
		); 

/******************* CELL 1383 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1383 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1287]),
			.N(gen[1288]),
			.NE(gen[1289]),

			.O(gen[1382]),
			.E(gen[1384]),

			.SO(gen[1477]),
			.S(gen[1478]),
			.SE(gen[1479]),

			.SELF(gen[1383]),
			.cell_state(gen[1383])
		); 

/******************* CELL 1384 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1384 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1288]),
			.N(gen[1289]),
			.NE(gen[1290]),

			.O(gen[1383]),
			.E(gen[1385]),

			.SO(gen[1478]),
			.S(gen[1479]),
			.SE(gen[1480]),

			.SELF(gen[1384]),
			.cell_state(gen[1384])
		); 

/******************* CELL 1385 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1385 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1289]),
			.N(gen[1290]),
			.NE(gen[1291]),

			.O(gen[1384]),
			.E(gen[1386]),

			.SO(gen[1479]),
			.S(gen[1480]),
			.SE(gen[1481]),

			.SELF(gen[1385]),
			.cell_state(gen[1385])
		); 

/******************* CELL 1386 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1386 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1290]),
			.N(gen[1291]),
			.NE(gen[1292]),

			.O(gen[1385]),
			.E(gen[1387]),

			.SO(gen[1480]),
			.S(gen[1481]),
			.SE(gen[1482]),

			.SELF(gen[1386]),
			.cell_state(gen[1386])
		); 

/******************* CELL 1387 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1387 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1291]),
			.N(gen[1292]),
			.NE(gen[1293]),

			.O(gen[1386]),
			.E(gen[1388]),

			.SO(gen[1481]),
			.S(gen[1482]),
			.SE(gen[1483]),

			.SELF(gen[1387]),
			.cell_state(gen[1387])
		); 

/******************* CELL 1388 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1388 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1292]),
			.N(gen[1293]),
			.NE(gen[1294]),

			.O(gen[1387]),
			.E(gen[1389]),

			.SO(gen[1482]),
			.S(gen[1483]),
			.SE(gen[1484]),

			.SELF(gen[1388]),
			.cell_state(gen[1388])
		); 

/******************* CELL 1389 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1389 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1293]),
			.N(gen[1294]),
			.NE(gen[1295]),

			.O(gen[1388]),
			.E(gen[1390]),

			.SO(gen[1483]),
			.S(gen[1484]),
			.SE(gen[1485]),

			.SELF(gen[1389]),
			.cell_state(gen[1389])
		); 

/******************* CELL 1390 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1390 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1294]),
			.N(gen[1295]),
			.NE(gen[1296]),

			.O(gen[1389]),
			.E(gen[1391]),

			.SO(gen[1484]),
			.S(gen[1485]),
			.SE(gen[1486]),

			.SELF(gen[1390]),
			.cell_state(gen[1390])
		); 

/******************* CELL 1391 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1391 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1295]),
			.N(gen[1296]),
			.NE(gen[1297]),

			.O(gen[1390]),
			.E(gen[1392]),

			.SO(gen[1485]),
			.S(gen[1486]),
			.SE(gen[1487]),

			.SELF(gen[1391]),
			.cell_state(gen[1391])
		); 

/******************* CELL 1392 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1392 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1296]),
			.N(gen[1297]),
			.NE(gen[1298]),

			.O(gen[1391]),
			.E(gen[1393]),

			.SO(gen[1486]),
			.S(gen[1487]),
			.SE(gen[1488]),

			.SELF(gen[1392]),
			.cell_state(gen[1392])
		); 

/******************* CELL 1393 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1393 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1297]),
			.N(gen[1298]),
			.NE(gen[1299]),

			.O(gen[1392]),
			.E(gen[1394]),

			.SO(gen[1487]),
			.S(gen[1488]),
			.SE(gen[1489]),

			.SELF(gen[1393]),
			.cell_state(gen[1393])
		); 

/******************* CELL 1394 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1394 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1298]),
			.N(gen[1299]),
			.NE(gen[1300]),

			.O(gen[1393]),
			.E(gen[1395]),

			.SO(gen[1488]),
			.S(gen[1489]),
			.SE(gen[1490]),

			.SELF(gen[1394]),
			.cell_state(gen[1394])
		); 

/******************* CELL 1395 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1395 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1299]),
			.N(gen[1300]),
			.NE(gen[1301]),

			.O(gen[1394]),
			.E(gen[1396]),

			.SO(gen[1489]),
			.S(gen[1490]),
			.SE(gen[1491]),

			.SELF(gen[1395]),
			.cell_state(gen[1395])
		); 

/******************* CELL 1396 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1396 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1300]),
			.N(gen[1301]),
			.NE(gen[1302]),

			.O(gen[1395]),
			.E(gen[1397]),

			.SO(gen[1490]),
			.S(gen[1491]),
			.SE(gen[1492]),

			.SELF(gen[1396]),
			.cell_state(gen[1396])
		); 

/******************* CELL 1397 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1397 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1301]),
			.N(gen[1302]),
			.NE(gen[1303]),

			.O(gen[1396]),
			.E(gen[1398]),

			.SO(gen[1491]),
			.S(gen[1492]),
			.SE(gen[1493]),

			.SELF(gen[1397]),
			.cell_state(gen[1397])
		); 

/******************* CELL 1398 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1398 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1302]),
			.N(gen[1303]),
			.NE(gen[1304]),

			.O(gen[1397]),
			.E(gen[1399]),

			.SO(gen[1492]),
			.S(gen[1493]),
			.SE(gen[1494]),

			.SELF(gen[1398]),
			.cell_state(gen[1398])
		); 

/******************* CELL 1399 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1399 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1303]),
			.N(gen[1304]),
			.NE(gen[1305]),

			.O(gen[1398]),
			.E(gen[1400]),

			.SO(gen[1493]),
			.S(gen[1494]),
			.SE(gen[1495]),

			.SELF(gen[1399]),
			.cell_state(gen[1399])
		); 

/******************* CELL 1400 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1400 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1304]),
			.N(gen[1305]),
			.NE(gen[1306]),

			.O(gen[1399]),
			.E(gen[1401]),

			.SO(gen[1494]),
			.S(gen[1495]),
			.SE(gen[1496]),

			.SELF(gen[1400]),
			.cell_state(gen[1400])
		); 

/******************* CELL 1401 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1401 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1305]),
			.N(gen[1306]),
			.NE(gen[1307]),

			.O(gen[1400]),
			.E(gen[1402]),

			.SO(gen[1495]),
			.S(gen[1496]),
			.SE(gen[1497]),

			.SELF(gen[1401]),
			.cell_state(gen[1401])
		); 

/******************* CELL 1402 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1402 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1306]),
			.N(gen[1307]),
			.NE(gen[1308]),

			.O(gen[1401]),
			.E(gen[1403]),

			.SO(gen[1496]),
			.S(gen[1497]),
			.SE(gen[1498]),

			.SELF(gen[1402]),
			.cell_state(gen[1402])
		); 

/******************* CELL 1403 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1403 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1307]),
			.N(gen[1308]),
			.NE(gen[1309]),

			.O(gen[1402]),
			.E(gen[1404]),

			.SO(gen[1497]),
			.S(gen[1498]),
			.SE(gen[1499]),

			.SELF(gen[1403]),
			.cell_state(gen[1403])
		); 

/******************* CELL 1404 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1404 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1308]),
			.N(gen[1309]),
			.NE(gen[1310]),

			.O(gen[1403]),
			.E(gen[1405]),

			.SO(gen[1498]),
			.S(gen[1499]),
			.SE(gen[1500]),

			.SELF(gen[1404]),
			.cell_state(gen[1404])
		); 

/******************* CELL 1405 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1405 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1309]),
			.N(gen[1310]),
			.NE(gen[1311]),

			.O(gen[1404]),
			.E(gen[1406]),

			.SO(gen[1499]),
			.S(gen[1500]),
			.SE(gen[1501]),

			.SELF(gen[1405]),
			.cell_state(gen[1405])
		); 

/******************* CELL 1406 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1406 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1310]),
			.N(gen[1311]),
			.NE(gen[1312]),

			.O(gen[1405]),
			.E(gen[1407]),

			.SO(gen[1500]),
			.S(gen[1501]),
			.SE(gen[1502]),

			.SELF(gen[1406]),
			.cell_state(gen[1406])
		); 

/******************* CELL 1407 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1407 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1311]),
			.N(gen[1312]),
			.NE(gen[1313]),

			.O(gen[1406]),
			.E(gen[1408]),

			.SO(gen[1501]),
			.S(gen[1502]),
			.SE(gen[1503]),

			.SELF(gen[1407]),
			.cell_state(gen[1407])
		); 

/******************* CELL 1408 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1408 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1312]),
			.N(gen[1313]),
			.NE(gen[1314]),

			.O(gen[1407]),
			.E(gen[1409]),

			.SO(gen[1502]),
			.S(gen[1503]),
			.SE(gen[1504]),

			.SELF(gen[1408]),
			.cell_state(gen[1408])
		); 

/******************* CELL 1409 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1409 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1313]),
			.N(gen[1314]),
			.NE(gen[1315]),

			.O(gen[1408]),
			.E(gen[1410]),

			.SO(gen[1503]),
			.S(gen[1504]),
			.SE(gen[1505]),

			.SELF(gen[1409]),
			.cell_state(gen[1409])
		); 

/******************* CELL 1410 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1410 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1314]),
			.N(gen[1315]),
			.NE(gen[1316]),

			.O(gen[1409]),
			.E(gen[1411]),

			.SO(gen[1504]),
			.S(gen[1505]),
			.SE(gen[1506]),

			.SELF(gen[1410]),
			.cell_state(gen[1410])
		); 

/******************* CELL 1411 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1411 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1315]),
			.N(gen[1316]),
			.NE(gen[1317]),

			.O(gen[1410]),
			.E(gen[1412]),

			.SO(gen[1505]),
			.S(gen[1506]),
			.SE(gen[1507]),

			.SELF(gen[1411]),
			.cell_state(gen[1411])
		); 

/******************* CELL 1412 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1412 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1316]),
			.N(gen[1317]),
			.NE(gen[1318]),

			.O(gen[1411]),
			.E(gen[1413]),

			.SO(gen[1506]),
			.S(gen[1507]),
			.SE(gen[1508]),

			.SELF(gen[1412]),
			.cell_state(gen[1412])
		); 

/******************* CELL 1413 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1413 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1317]),
			.N(gen[1318]),
			.NE(gen[1319]),

			.O(gen[1412]),
			.E(gen[1414]),

			.SO(gen[1507]),
			.S(gen[1508]),
			.SE(gen[1509]),

			.SELF(gen[1413]),
			.cell_state(gen[1413])
		); 

/******************* CELL 1414 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1414 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1318]),
			.N(gen[1319]),
			.NE(gen[1320]),

			.O(gen[1413]),
			.E(gen[1415]),

			.SO(gen[1508]),
			.S(gen[1509]),
			.SE(gen[1510]),

			.SELF(gen[1414]),
			.cell_state(gen[1414])
		); 

/******************* CELL 1415 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1415 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1319]),
			.N(gen[1320]),
			.NE(gen[1321]),

			.O(gen[1414]),
			.E(gen[1416]),

			.SO(gen[1509]),
			.S(gen[1510]),
			.SE(gen[1511]),

			.SELF(gen[1415]),
			.cell_state(gen[1415])
		); 

/******************* CELL 1416 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1416 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1320]),
			.N(gen[1321]),
			.NE(gen[1322]),

			.O(gen[1415]),
			.E(gen[1417]),

			.SO(gen[1510]),
			.S(gen[1511]),
			.SE(gen[1512]),

			.SELF(gen[1416]),
			.cell_state(gen[1416])
		); 

/******************* CELL 1417 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1417 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1321]),
			.N(gen[1322]),
			.NE(gen[1323]),

			.O(gen[1416]),
			.E(gen[1418]),

			.SO(gen[1511]),
			.S(gen[1512]),
			.SE(gen[1513]),

			.SELF(gen[1417]),
			.cell_state(gen[1417])
		); 

/******************* CELL 1418 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1418 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1322]),
			.N(gen[1323]),
			.NE(gen[1324]),

			.O(gen[1417]),
			.E(gen[1419]),

			.SO(gen[1512]),
			.S(gen[1513]),
			.SE(gen[1514]),

			.SELF(gen[1418]),
			.cell_state(gen[1418])
		); 

/******************* CELL 1419 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1419 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1323]),
			.N(gen[1324]),
			.NE(gen[1325]),

			.O(gen[1418]),
			.E(gen[1420]),

			.SO(gen[1513]),
			.S(gen[1514]),
			.SE(gen[1515]),

			.SELF(gen[1419]),
			.cell_state(gen[1419])
		); 

/******************* CELL 1420 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1420 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1324]),
			.N(gen[1325]),
			.NE(gen[1326]),

			.O(gen[1419]),
			.E(gen[1421]),

			.SO(gen[1514]),
			.S(gen[1515]),
			.SE(gen[1516]),

			.SELF(gen[1420]),
			.cell_state(gen[1420])
		); 

/******************* CELL 1421 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1421 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1325]),
			.N(gen[1326]),
			.NE(gen[1327]),

			.O(gen[1420]),
			.E(gen[1422]),

			.SO(gen[1515]),
			.S(gen[1516]),
			.SE(gen[1517]),

			.SELF(gen[1421]),
			.cell_state(gen[1421])
		); 

/******************* CELL 1422 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1422 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1326]),
			.N(gen[1327]),
			.NE(gen[1328]),

			.O(gen[1421]),
			.E(gen[1423]),

			.SO(gen[1516]),
			.S(gen[1517]),
			.SE(gen[1518]),

			.SELF(gen[1422]),
			.cell_state(gen[1422])
		); 

/******************* CELL 1423 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1423 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1327]),
			.N(gen[1328]),
			.NE(gen[1329]),

			.O(gen[1422]),
			.E(gen[1424]),

			.SO(gen[1517]),
			.S(gen[1518]),
			.SE(gen[1519]),

			.SELF(gen[1423]),
			.cell_state(gen[1423])
		); 

/******************* CELL 1424 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1424 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1328]),
			.N(gen[1329]),
			.NE(gen[1328]),

			.O(gen[1423]),
			.E(gen[1423]),

			.SO(gen[1518]),
			.S(gen[1519]),
			.SE(gen[1518]),

			.SELF(gen[1424]),
			.cell_state(gen[1424])
		); 

/******************* CELL 1425 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1425 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1331]),
			.N(gen[1330]),
			.NE(gen[1331]),

			.O(gen[1426]),
			.E(gen[1426]),

			.SO(gen[1521]),
			.S(gen[1520]),
			.SE(gen[1521]),

			.SELF(gen[1425]),
			.cell_state(gen[1425])
		); 

/******************* CELL 1426 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1426 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1330]),
			.N(gen[1331]),
			.NE(gen[1332]),

			.O(gen[1425]),
			.E(gen[1427]),

			.SO(gen[1520]),
			.S(gen[1521]),
			.SE(gen[1522]),

			.SELF(gen[1426]),
			.cell_state(gen[1426])
		); 

/******************* CELL 1427 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1427 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1331]),
			.N(gen[1332]),
			.NE(gen[1333]),

			.O(gen[1426]),
			.E(gen[1428]),

			.SO(gen[1521]),
			.S(gen[1522]),
			.SE(gen[1523]),

			.SELF(gen[1427]),
			.cell_state(gen[1427])
		); 

/******************* CELL 1428 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1428 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1332]),
			.N(gen[1333]),
			.NE(gen[1334]),

			.O(gen[1427]),
			.E(gen[1429]),

			.SO(gen[1522]),
			.S(gen[1523]),
			.SE(gen[1524]),

			.SELF(gen[1428]),
			.cell_state(gen[1428])
		); 

/******************* CELL 1429 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1429 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1333]),
			.N(gen[1334]),
			.NE(gen[1335]),

			.O(gen[1428]),
			.E(gen[1430]),

			.SO(gen[1523]),
			.S(gen[1524]),
			.SE(gen[1525]),

			.SELF(gen[1429]),
			.cell_state(gen[1429])
		); 

/******************* CELL 1430 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1430 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1334]),
			.N(gen[1335]),
			.NE(gen[1336]),

			.O(gen[1429]),
			.E(gen[1431]),

			.SO(gen[1524]),
			.S(gen[1525]),
			.SE(gen[1526]),

			.SELF(gen[1430]),
			.cell_state(gen[1430])
		); 

/******************* CELL 1431 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1431 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1335]),
			.N(gen[1336]),
			.NE(gen[1337]),

			.O(gen[1430]),
			.E(gen[1432]),

			.SO(gen[1525]),
			.S(gen[1526]),
			.SE(gen[1527]),

			.SELF(gen[1431]),
			.cell_state(gen[1431])
		); 

/******************* CELL 1432 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1432 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1336]),
			.N(gen[1337]),
			.NE(gen[1338]),

			.O(gen[1431]),
			.E(gen[1433]),

			.SO(gen[1526]),
			.S(gen[1527]),
			.SE(gen[1528]),

			.SELF(gen[1432]),
			.cell_state(gen[1432])
		); 

/******************* CELL 1433 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1433 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1337]),
			.N(gen[1338]),
			.NE(gen[1339]),

			.O(gen[1432]),
			.E(gen[1434]),

			.SO(gen[1527]),
			.S(gen[1528]),
			.SE(gen[1529]),

			.SELF(gen[1433]),
			.cell_state(gen[1433])
		); 

/******************* CELL 1434 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1434 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1338]),
			.N(gen[1339]),
			.NE(gen[1340]),

			.O(gen[1433]),
			.E(gen[1435]),

			.SO(gen[1528]),
			.S(gen[1529]),
			.SE(gen[1530]),

			.SELF(gen[1434]),
			.cell_state(gen[1434])
		); 

/******************* CELL 1435 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1435 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1339]),
			.N(gen[1340]),
			.NE(gen[1341]),

			.O(gen[1434]),
			.E(gen[1436]),

			.SO(gen[1529]),
			.S(gen[1530]),
			.SE(gen[1531]),

			.SELF(gen[1435]),
			.cell_state(gen[1435])
		); 

/******************* CELL 1436 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1436 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1340]),
			.N(gen[1341]),
			.NE(gen[1342]),

			.O(gen[1435]),
			.E(gen[1437]),

			.SO(gen[1530]),
			.S(gen[1531]),
			.SE(gen[1532]),

			.SELF(gen[1436]),
			.cell_state(gen[1436])
		); 

/******************* CELL 1437 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1437 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1341]),
			.N(gen[1342]),
			.NE(gen[1343]),

			.O(gen[1436]),
			.E(gen[1438]),

			.SO(gen[1531]),
			.S(gen[1532]),
			.SE(gen[1533]),

			.SELF(gen[1437]),
			.cell_state(gen[1437])
		); 

/******************* CELL 1438 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1438 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1342]),
			.N(gen[1343]),
			.NE(gen[1344]),

			.O(gen[1437]),
			.E(gen[1439]),

			.SO(gen[1532]),
			.S(gen[1533]),
			.SE(gen[1534]),

			.SELF(gen[1438]),
			.cell_state(gen[1438])
		); 

/******************* CELL 1439 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1439 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1343]),
			.N(gen[1344]),
			.NE(gen[1345]),

			.O(gen[1438]),
			.E(gen[1440]),

			.SO(gen[1533]),
			.S(gen[1534]),
			.SE(gen[1535]),

			.SELF(gen[1439]),
			.cell_state(gen[1439])
		); 

/******************* CELL 1440 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1440 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1344]),
			.N(gen[1345]),
			.NE(gen[1346]),

			.O(gen[1439]),
			.E(gen[1441]),

			.SO(gen[1534]),
			.S(gen[1535]),
			.SE(gen[1536]),

			.SELF(gen[1440]),
			.cell_state(gen[1440])
		); 

/******************* CELL 1441 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1441 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1345]),
			.N(gen[1346]),
			.NE(gen[1347]),

			.O(gen[1440]),
			.E(gen[1442]),

			.SO(gen[1535]),
			.S(gen[1536]),
			.SE(gen[1537]),

			.SELF(gen[1441]),
			.cell_state(gen[1441])
		); 

/******************* CELL 1442 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1442 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1346]),
			.N(gen[1347]),
			.NE(gen[1348]),

			.O(gen[1441]),
			.E(gen[1443]),

			.SO(gen[1536]),
			.S(gen[1537]),
			.SE(gen[1538]),

			.SELF(gen[1442]),
			.cell_state(gen[1442])
		); 

/******************* CELL 1443 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1443 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1347]),
			.N(gen[1348]),
			.NE(gen[1349]),

			.O(gen[1442]),
			.E(gen[1444]),

			.SO(gen[1537]),
			.S(gen[1538]),
			.SE(gen[1539]),

			.SELF(gen[1443]),
			.cell_state(gen[1443])
		); 

/******************* CELL 1444 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1444 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1348]),
			.N(gen[1349]),
			.NE(gen[1350]),

			.O(gen[1443]),
			.E(gen[1445]),

			.SO(gen[1538]),
			.S(gen[1539]),
			.SE(gen[1540]),

			.SELF(gen[1444]),
			.cell_state(gen[1444])
		); 

/******************* CELL 1445 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1445 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1349]),
			.N(gen[1350]),
			.NE(gen[1351]),

			.O(gen[1444]),
			.E(gen[1446]),

			.SO(gen[1539]),
			.S(gen[1540]),
			.SE(gen[1541]),

			.SELF(gen[1445]),
			.cell_state(gen[1445])
		); 

/******************* CELL 1446 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1446 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1350]),
			.N(gen[1351]),
			.NE(gen[1352]),

			.O(gen[1445]),
			.E(gen[1447]),

			.SO(gen[1540]),
			.S(gen[1541]),
			.SE(gen[1542]),

			.SELF(gen[1446]),
			.cell_state(gen[1446])
		); 

/******************* CELL 1447 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1447 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1351]),
			.N(gen[1352]),
			.NE(gen[1353]),

			.O(gen[1446]),
			.E(gen[1448]),

			.SO(gen[1541]),
			.S(gen[1542]),
			.SE(gen[1543]),

			.SELF(gen[1447]),
			.cell_state(gen[1447])
		); 

/******************* CELL 1448 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1448 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1352]),
			.N(gen[1353]),
			.NE(gen[1354]),

			.O(gen[1447]),
			.E(gen[1449]),

			.SO(gen[1542]),
			.S(gen[1543]),
			.SE(gen[1544]),

			.SELF(gen[1448]),
			.cell_state(gen[1448])
		); 

/******************* CELL 1449 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1449 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1353]),
			.N(gen[1354]),
			.NE(gen[1355]),

			.O(gen[1448]),
			.E(gen[1450]),

			.SO(gen[1543]),
			.S(gen[1544]),
			.SE(gen[1545]),

			.SELF(gen[1449]),
			.cell_state(gen[1449])
		); 

/******************* CELL 1450 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1450 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1354]),
			.N(gen[1355]),
			.NE(gen[1356]),

			.O(gen[1449]),
			.E(gen[1451]),

			.SO(gen[1544]),
			.S(gen[1545]),
			.SE(gen[1546]),

			.SELF(gen[1450]),
			.cell_state(gen[1450])
		); 

/******************* CELL 1451 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1451 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1355]),
			.N(gen[1356]),
			.NE(gen[1357]),

			.O(gen[1450]),
			.E(gen[1452]),

			.SO(gen[1545]),
			.S(gen[1546]),
			.SE(gen[1547]),

			.SELF(gen[1451]),
			.cell_state(gen[1451])
		); 

/******************* CELL 1452 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1452 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1356]),
			.N(gen[1357]),
			.NE(gen[1358]),

			.O(gen[1451]),
			.E(gen[1453]),

			.SO(gen[1546]),
			.S(gen[1547]),
			.SE(gen[1548]),

			.SELF(gen[1452]),
			.cell_state(gen[1452])
		); 

/******************* CELL 1453 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1453 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1357]),
			.N(gen[1358]),
			.NE(gen[1359]),

			.O(gen[1452]),
			.E(gen[1454]),

			.SO(gen[1547]),
			.S(gen[1548]),
			.SE(gen[1549]),

			.SELF(gen[1453]),
			.cell_state(gen[1453])
		); 

/******************* CELL 1454 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1454 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1358]),
			.N(gen[1359]),
			.NE(gen[1360]),

			.O(gen[1453]),
			.E(gen[1455]),

			.SO(gen[1548]),
			.S(gen[1549]),
			.SE(gen[1550]),

			.SELF(gen[1454]),
			.cell_state(gen[1454])
		); 

/******************* CELL 1455 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1455 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1359]),
			.N(gen[1360]),
			.NE(gen[1361]),

			.O(gen[1454]),
			.E(gen[1456]),

			.SO(gen[1549]),
			.S(gen[1550]),
			.SE(gen[1551]),

			.SELF(gen[1455]),
			.cell_state(gen[1455])
		); 

/******************* CELL 1456 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1456 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1360]),
			.N(gen[1361]),
			.NE(gen[1362]),

			.O(gen[1455]),
			.E(gen[1457]),

			.SO(gen[1550]),
			.S(gen[1551]),
			.SE(gen[1552]),

			.SELF(gen[1456]),
			.cell_state(gen[1456])
		); 

/******************* CELL 1457 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1457 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1361]),
			.N(gen[1362]),
			.NE(gen[1363]),

			.O(gen[1456]),
			.E(gen[1458]),

			.SO(gen[1551]),
			.S(gen[1552]),
			.SE(gen[1553]),

			.SELF(gen[1457]),
			.cell_state(gen[1457])
		); 

/******************* CELL 1458 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1458 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1362]),
			.N(gen[1363]),
			.NE(gen[1364]),

			.O(gen[1457]),
			.E(gen[1459]),

			.SO(gen[1552]),
			.S(gen[1553]),
			.SE(gen[1554]),

			.SELF(gen[1458]),
			.cell_state(gen[1458])
		); 

/******************* CELL 1459 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1459 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1363]),
			.N(gen[1364]),
			.NE(gen[1365]),

			.O(gen[1458]),
			.E(gen[1460]),

			.SO(gen[1553]),
			.S(gen[1554]),
			.SE(gen[1555]),

			.SELF(gen[1459]),
			.cell_state(gen[1459])
		); 

/******************* CELL 1460 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1460 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1364]),
			.N(gen[1365]),
			.NE(gen[1366]),

			.O(gen[1459]),
			.E(gen[1461]),

			.SO(gen[1554]),
			.S(gen[1555]),
			.SE(gen[1556]),

			.SELF(gen[1460]),
			.cell_state(gen[1460])
		); 

/******************* CELL 1461 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1461 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1365]),
			.N(gen[1366]),
			.NE(gen[1367]),

			.O(gen[1460]),
			.E(gen[1462]),

			.SO(gen[1555]),
			.S(gen[1556]),
			.SE(gen[1557]),

			.SELF(gen[1461]),
			.cell_state(gen[1461])
		); 

/******************* CELL 1462 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1462 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1366]),
			.N(gen[1367]),
			.NE(gen[1368]),

			.O(gen[1461]),
			.E(gen[1463]),

			.SO(gen[1556]),
			.S(gen[1557]),
			.SE(gen[1558]),

			.SELF(gen[1462]),
			.cell_state(gen[1462])
		); 

/******************* CELL 1463 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1463 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1367]),
			.N(gen[1368]),
			.NE(gen[1369]),

			.O(gen[1462]),
			.E(gen[1464]),

			.SO(gen[1557]),
			.S(gen[1558]),
			.SE(gen[1559]),

			.SELF(gen[1463]),
			.cell_state(gen[1463])
		); 

/******************* CELL 1464 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1464 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1368]),
			.N(gen[1369]),
			.NE(gen[1370]),

			.O(gen[1463]),
			.E(gen[1465]),

			.SO(gen[1558]),
			.S(gen[1559]),
			.SE(gen[1560]),

			.SELF(gen[1464]),
			.cell_state(gen[1464])
		); 

/******************* CELL 1465 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1465 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1369]),
			.N(gen[1370]),
			.NE(gen[1371]),

			.O(gen[1464]),
			.E(gen[1466]),

			.SO(gen[1559]),
			.S(gen[1560]),
			.SE(gen[1561]),

			.SELF(gen[1465]),
			.cell_state(gen[1465])
		); 

/******************* CELL 1466 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1466 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1370]),
			.N(gen[1371]),
			.NE(gen[1372]),

			.O(gen[1465]),
			.E(gen[1467]),

			.SO(gen[1560]),
			.S(gen[1561]),
			.SE(gen[1562]),

			.SELF(gen[1466]),
			.cell_state(gen[1466])
		); 

/******************* CELL 1467 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1467 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1371]),
			.N(gen[1372]),
			.NE(gen[1373]),

			.O(gen[1466]),
			.E(gen[1468]),

			.SO(gen[1561]),
			.S(gen[1562]),
			.SE(gen[1563]),

			.SELF(gen[1467]),
			.cell_state(gen[1467])
		); 

/******************* CELL 1468 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1468 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1372]),
			.N(gen[1373]),
			.NE(gen[1374]),

			.O(gen[1467]),
			.E(gen[1469]),

			.SO(gen[1562]),
			.S(gen[1563]),
			.SE(gen[1564]),

			.SELF(gen[1468]),
			.cell_state(gen[1468])
		); 

/******************* CELL 1469 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1469 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1373]),
			.N(gen[1374]),
			.NE(gen[1375]),

			.O(gen[1468]),
			.E(gen[1470]),

			.SO(gen[1563]),
			.S(gen[1564]),
			.SE(gen[1565]),

			.SELF(gen[1469]),
			.cell_state(gen[1469])
		); 

/******************* CELL 1470 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1470 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1374]),
			.N(gen[1375]),
			.NE(gen[1376]),

			.O(gen[1469]),
			.E(gen[1471]),

			.SO(gen[1564]),
			.S(gen[1565]),
			.SE(gen[1566]),

			.SELF(gen[1470]),
			.cell_state(gen[1470])
		); 

/******************* CELL 1471 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1471 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1375]),
			.N(gen[1376]),
			.NE(gen[1377]),

			.O(gen[1470]),
			.E(gen[1472]),

			.SO(gen[1565]),
			.S(gen[1566]),
			.SE(gen[1567]),

			.SELF(gen[1471]),
			.cell_state(gen[1471])
		); 

/******************* CELL 1472 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1472 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1376]),
			.N(gen[1377]),
			.NE(gen[1378]),

			.O(gen[1471]),
			.E(gen[1473]),

			.SO(gen[1566]),
			.S(gen[1567]),
			.SE(gen[1568]),

			.SELF(gen[1472]),
			.cell_state(gen[1472])
		); 

/******************* CELL 1473 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1473 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1377]),
			.N(gen[1378]),
			.NE(gen[1379]),

			.O(gen[1472]),
			.E(gen[1474]),

			.SO(gen[1567]),
			.S(gen[1568]),
			.SE(gen[1569]),

			.SELF(gen[1473]),
			.cell_state(gen[1473])
		); 

/******************* CELL 1474 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1474 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1378]),
			.N(gen[1379]),
			.NE(gen[1380]),

			.O(gen[1473]),
			.E(gen[1475]),

			.SO(gen[1568]),
			.S(gen[1569]),
			.SE(gen[1570]),

			.SELF(gen[1474]),
			.cell_state(gen[1474])
		); 

/******************* CELL 1475 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1475 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1379]),
			.N(gen[1380]),
			.NE(gen[1381]),

			.O(gen[1474]),
			.E(gen[1476]),

			.SO(gen[1569]),
			.S(gen[1570]),
			.SE(gen[1571]),

			.SELF(gen[1475]),
			.cell_state(gen[1475])
		); 

/******************* CELL 1476 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1476 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1380]),
			.N(gen[1381]),
			.NE(gen[1382]),

			.O(gen[1475]),
			.E(gen[1477]),

			.SO(gen[1570]),
			.S(gen[1571]),
			.SE(gen[1572]),

			.SELF(gen[1476]),
			.cell_state(gen[1476])
		); 

/******************* CELL 1477 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1477 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1381]),
			.N(gen[1382]),
			.NE(gen[1383]),

			.O(gen[1476]),
			.E(gen[1478]),

			.SO(gen[1571]),
			.S(gen[1572]),
			.SE(gen[1573]),

			.SELF(gen[1477]),
			.cell_state(gen[1477])
		); 

/******************* CELL 1478 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1478 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1382]),
			.N(gen[1383]),
			.NE(gen[1384]),

			.O(gen[1477]),
			.E(gen[1479]),

			.SO(gen[1572]),
			.S(gen[1573]),
			.SE(gen[1574]),

			.SELF(gen[1478]),
			.cell_state(gen[1478])
		); 

/******************* CELL 1479 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1479 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1383]),
			.N(gen[1384]),
			.NE(gen[1385]),

			.O(gen[1478]),
			.E(gen[1480]),

			.SO(gen[1573]),
			.S(gen[1574]),
			.SE(gen[1575]),

			.SELF(gen[1479]),
			.cell_state(gen[1479])
		); 

/******************* CELL 1480 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1480 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1384]),
			.N(gen[1385]),
			.NE(gen[1386]),

			.O(gen[1479]),
			.E(gen[1481]),

			.SO(gen[1574]),
			.S(gen[1575]),
			.SE(gen[1576]),

			.SELF(gen[1480]),
			.cell_state(gen[1480])
		); 

/******************* CELL 1481 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1481 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1385]),
			.N(gen[1386]),
			.NE(gen[1387]),

			.O(gen[1480]),
			.E(gen[1482]),

			.SO(gen[1575]),
			.S(gen[1576]),
			.SE(gen[1577]),

			.SELF(gen[1481]),
			.cell_state(gen[1481])
		); 

/******************* CELL 1482 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1482 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1386]),
			.N(gen[1387]),
			.NE(gen[1388]),

			.O(gen[1481]),
			.E(gen[1483]),

			.SO(gen[1576]),
			.S(gen[1577]),
			.SE(gen[1578]),

			.SELF(gen[1482]),
			.cell_state(gen[1482])
		); 

/******************* CELL 1483 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1483 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1387]),
			.N(gen[1388]),
			.NE(gen[1389]),

			.O(gen[1482]),
			.E(gen[1484]),

			.SO(gen[1577]),
			.S(gen[1578]),
			.SE(gen[1579]),

			.SELF(gen[1483]),
			.cell_state(gen[1483])
		); 

/******************* CELL 1484 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1484 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1388]),
			.N(gen[1389]),
			.NE(gen[1390]),

			.O(gen[1483]),
			.E(gen[1485]),

			.SO(gen[1578]),
			.S(gen[1579]),
			.SE(gen[1580]),

			.SELF(gen[1484]),
			.cell_state(gen[1484])
		); 

/******************* CELL 1485 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1485 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1389]),
			.N(gen[1390]),
			.NE(gen[1391]),

			.O(gen[1484]),
			.E(gen[1486]),

			.SO(gen[1579]),
			.S(gen[1580]),
			.SE(gen[1581]),

			.SELF(gen[1485]),
			.cell_state(gen[1485])
		); 

/******************* CELL 1486 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1486 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1390]),
			.N(gen[1391]),
			.NE(gen[1392]),

			.O(gen[1485]),
			.E(gen[1487]),

			.SO(gen[1580]),
			.S(gen[1581]),
			.SE(gen[1582]),

			.SELF(gen[1486]),
			.cell_state(gen[1486])
		); 

/******************* CELL 1487 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1487 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1391]),
			.N(gen[1392]),
			.NE(gen[1393]),

			.O(gen[1486]),
			.E(gen[1488]),

			.SO(gen[1581]),
			.S(gen[1582]),
			.SE(gen[1583]),

			.SELF(gen[1487]),
			.cell_state(gen[1487])
		); 

/******************* CELL 1488 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1488 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1392]),
			.N(gen[1393]),
			.NE(gen[1394]),

			.O(gen[1487]),
			.E(gen[1489]),

			.SO(gen[1582]),
			.S(gen[1583]),
			.SE(gen[1584]),

			.SELF(gen[1488]),
			.cell_state(gen[1488])
		); 

/******************* CELL 1489 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1489 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1393]),
			.N(gen[1394]),
			.NE(gen[1395]),

			.O(gen[1488]),
			.E(gen[1490]),

			.SO(gen[1583]),
			.S(gen[1584]),
			.SE(gen[1585]),

			.SELF(gen[1489]),
			.cell_state(gen[1489])
		); 

/******************* CELL 1490 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1490 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1394]),
			.N(gen[1395]),
			.NE(gen[1396]),

			.O(gen[1489]),
			.E(gen[1491]),

			.SO(gen[1584]),
			.S(gen[1585]),
			.SE(gen[1586]),

			.SELF(gen[1490]),
			.cell_state(gen[1490])
		); 

/******************* CELL 1491 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1491 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1395]),
			.N(gen[1396]),
			.NE(gen[1397]),

			.O(gen[1490]),
			.E(gen[1492]),

			.SO(gen[1585]),
			.S(gen[1586]),
			.SE(gen[1587]),

			.SELF(gen[1491]),
			.cell_state(gen[1491])
		); 

/******************* CELL 1492 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1492 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1396]),
			.N(gen[1397]),
			.NE(gen[1398]),

			.O(gen[1491]),
			.E(gen[1493]),

			.SO(gen[1586]),
			.S(gen[1587]),
			.SE(gen[1588]),

			.SELF(gen[1492]),
			.cell_state(gen[1492])
		); 

/******************* CELL 1493 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1493 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1397]),
			.N(gen[1398]),
			.NE(gen[1399]),

			.O(gen[1492]),
			.E(gen[1494]),

			.SO(gen[1587]),
			.S(gen[1588]),
			.SE(gen[1589]),

			.SELF(gen[1493]),
			.cell_state(gen[1493])
		); 

/******************* CELL 1494 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1494 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1398]),
			.N(gen[1399]),
			.NE(gen[1400]),

			.O(gen[1493]),
			.E(gen[1495]),

			.SO(gen[1588]),
			.S(gen[1589]),
			.SE(gen[1590]),

			.SELF(gen[1494]),
			.cell_state(gen[1494])
		); 

/******************* CELL 1495 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1495 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1399]),
			.N(gen[1400]),
			.NE(gen[1401]),

			.O(gen[1494]),
			.E(gen[1496]),

			.SO(gen[1589]),
			.S(gen[1590]),
			.SE(gen[1591]),

			.SELF(gen[1495]),
			.cell_state(gen[1495])
		); 

/******************* CELL 1496 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1496 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1400]),
			.N(gen[1401]),
			.NE(gen[1402]),

			.O(gen[1495]),
			.E(gen[1497]),

			.SO(gen[1590]),
			.S(gen[1591]),
			.SE(gen[1592]),

			.SELF(gen[1496]),
			.cell_state(gen[1496])
		); 

/******************* CELL 1497 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1497 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1401]),
			.N(gen[1402]),
			.NE(gen[1403]),

			.O(gen[1496]),
			.E(gen[1498]),

			.SO(gen[1591]),
			.S(gen[1592]),
			.SE(gen[1593]),

			.SELF(gen[1497]),
			.cell_state(gen[1497])
		); 

/******************* CELL 1498 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1498 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1402]),
			.N(gen[1403]),
			.NE(gen[1404]),

			.O(gen[1497]),
			.E(gen[1499]),

			.SO(gen[1592]),
			.S(gen[1593]),
			.SE(gen[1594]),

			.SELF(gen[1498]),
			.cell_state(gen[1498])
		); 

/******************* CELL 1499 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1499 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1403]),
			.N(gen[1404]),
			.NE(gen[1405]),

			.O(gen[1498]),
			.E(gen[1500]),

			.SO(gen[1593]),
			.S(gen[1594]),
			.SE(gen[1595]),

			.SELF(gen[1499]),
			.cell_state(gen[1499])
		); 

/******************* CELL 1500 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1500 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1404]),
			.N(gen[1405]),
			.NE(gen[1406]),

			.O(gen[1499]),
			.E(gen[1501]),

			.SO(gen[1594]),
			.S(gen[1595]),
			.SE(gen[1596]),

			.SELF(gen[1500]),
			.cell_state(gen[1500])
		); 

/******************* CELL 1501 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1501 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1405]),
			.N(gen[1406]),
			.NE(gen[1407]),

			.O(gen[1500]),
			.E(gen[1502]),

			.SO(gen[1595]),
			.S(gen[1596]),
			.SE(gen[1597]),

			.SELF(gen[1501]),
			.cell_state(gen[1501])
		); 

/******************* CELL 1502 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1502 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1406]),
			.N(gen[1407]),
			.NE(gen[1408]),

			.O(gen[1501]),
			.E(gen[1503]),

			.SO(gen[1596]),
			.S(gen[1597]),
			.SE(gen[1598]),

			.SELF(gen[1502]),
			.cell_state(gen[1502])
		); 

/******************* CELL 1503 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1503 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1407]),
			.N(gen[1408]),
			.NE(gen[1409]),

			.O(gen[1502]),
			.E(gen[1504]),

			.SO(gen[1597]),
			.S(gen[1598]),
			.SE(gen[1599]),

			.SELF(gen[1503]),
			.cell_state(gen[1503])
		); 

/******************* CELL 1504 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1504 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1408]),
			.N(gen[1409]),
			.NE(gen[1410]),

			.O(gen[1503]),
			.E(gen[1505]),

			.SO(gen[1598]),
			.S(gen[1599]),
			.SE(gen[1600]),

			.SELF(gen[1504]),
			.cell_state(gen[1504])
		); 

/******************* CELL 1505 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1505 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1409]),
			.N(gen[1410]),
			.NE(gen[1411]),

			.O(gen[1504]),
			.E(gen[1506]),

			.SO(gen[1599]),
			.S(gen[1600]),
			.SE(gen[1601]),

			.SELF(gen[1505]),
			.cell_state(gen[1505])
		); 

/******************* CELL 1506 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1506 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1410]),
			.N(gen[1411]),
			.NE(gen[1412]),

			.O(gen[1505]),
			.E(gen[1507]),

			.SO(gen[1600]),
			.S(gen[1601]),
			.SE(gen[1602]),

			.SELF(gen[1506]),
			.cell_state(gen[1506])
		); 

/******************* CELL 1507 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1507 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1411]),
			.N(gen[1412]),
			.NE(gen[1413]),

			.O(gen[1506]),
			.E(gen[1508]),

			.SO(gen[1601]),
			.S(gen[1602]),
			.SE(gen[1603]),

			.SELF(gen[1507]),
			.cell_state(gen[1507])
		); 

/******************* CELL 1508 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1508 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1412]),
			.N(gen[1413]),
			.NE(gen[1414]),

			.O(gen[1507]),
			.E(gen[1509]),

			.SO(gen[1602]),
			.S(gen[1603]),
			.SE(gen[1604]),

			.SELF(gen[1508]),
			.cell_state(gen[1508])
		); 

/******************* CELL 1509 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1509 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1413]),
			.N(gen[1414]),
			.NE(gen[1415]),

			.O(gen[1508]),
			.E(gen[1510]),

			.SO(gen[1603]),
			.S(gen[1604]),
			.SE(gen[1605]),

			.SELF(gen[1509]),
			.cell_state(gen[1509])
		); 

/******************* CELL 1510 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1510 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1414]),
			.N(gen[1415]),
			.NE(gen[1416]),

			.O(gen[1509]),
			.E(gen[1511]),

			.SO(gen[1604]),
			.S(gen[1605]),
			.SE(gen[1606]),

			.SELF(gen[1510]),
			.cell_state(gen[1510])
		); 

/******************* CELL 1511 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1511 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1415]),
			.N(gen[1416]),
			.NE(gen[1417]),

			.O(gen[1510]),
			.E(gen[1512]),

			.SO(gen[1605]),
			.S(gen[1606]),
			.SE(gen[1607]),

			.SELF(gen[1511]),
			.cell_state(gen[1511])
		); 

/******************* CELL 1512 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1512 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1416]),
			.N(gen[1417]),
			.NE(gen[1418]),

			.O(gen[1511]),
			.E(gen[1513]),

			.SO(gen[1606]),
			.S(gen[1607]),
			.SE(gen[1608]),

			.SELF(gen[1512]),
			.cell_state(gen[1512])
		); 

/******************* CELL 1513 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1513 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1417]),
			.N(gen[1418]),
			.NE(gen[1419]),

			.O(gen[1512]),
			.E(gen[1514]),

			.SO(gen[1607]),
			.S(gen[1608]),
			.SE(gen[1609]),

			.SELF(gen[1513]),
			.cell_state(gen[1513])
		); 

/******************* CELL 1514 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1514 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1418]),
			.N(gen[1419]),
			.NE(gen[1420]),

			.O(gen[1513]),
			.E(gen[1515]),

			.SO(gen[1608]),
			.S(gen[1609]),
			.SE(gen[1610]),

			.SELF(gen[1514]),
			.cell_state(gen[1514])
		); 

/******************* CELL 1515 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1515 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1419]),
			.N(gen[1420]),
			.NE(gen[1421]),

			.O(gen[1514]),
			.E(gen[1516]),

			.SO(gen[1609]),
			.S(gen[1610]),
			.SE(gen[1611]),

			.SELF(gen[1515]),
			.cell_state(gen[1515])
		); 

/******************* CELL 1516 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1516 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1420]),
			.N(gen[1421]),
			.NE(gen[1422]),

			.O(gen[1515]),
			.E(gen[1517]),

			.SO(gen[1610]),
			.S(gen[1611]),
			.SE(gen[1612]),

			.SELF(gen[1516]),
			.cell_state(gen[1516])
		); 

/******************* CELL 1517 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1517 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1421]),
			.N(gen[1422]),
			.NE(gen[1423]),

			.O(gen[1516]),
			.E(gen[1518]),

			.SO(gen[1611]),
			.S(gen[1612]),
			.SE(gen[1613]),

			.SELF(gen[1517]),
			.cell_state(gen[1517])
		); 

/******************* CELL 1518 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1518 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1422]),
			.N(gen[1423]),
			.NE(gen[1424]),

			.O(gen[1517]),
			.E(gen[1519]),

			.SO(gen[1612]),
			.S(gen[1613]),
			.SE(gen[1614]),

			.SELF(gen[1518]),
			.cell_state(gen[1518])
		); 

/******************* CELL 1519 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1519 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1423]),
			.N(gen[1424]),
			.NE(gen[1423]),

			.O(gen[1518]),
			.E(gen[1518]),

			.SO(gen[1613]),
			.S(gen[1614]),
			.SE(gen[1613]),

			.SELF(gen[1519]),
			.cell_state(gen[1519])
		); 

/******************* CELL 1520 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1520 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1426]),
			.N(gen[1425]),
			.NE(gen[1426]),

			.O(gen[1521]),
			.E(gen[1521]),

			.SO(gen[1616]),
			.S(gen[1615]),
			.SE(gen[1616]),

			.SELF(gen[1520]),
			.cell_state(gen[1520])
		); 

/******************* CELL 1521 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1521 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1425]),
			.N(gen[1426]),
			.NE(gen[1427]),

			.O(gen[1520]),
			.E(gen[1522]),

			.SO(gen[1615]),
			.S(gen[1616]),
			.SE(gen[1617]),

			.SELF(gen[1521]),
			.cell_state(gen[1521])
		); 

/******************* CELL 1522 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1522 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1426]),
			.N(gen[1427]),
			.NE(gen[1428]),

			.O(gen[1521]),
			.E(gen[1523]),

			.SO(gen[1616]),
			.S(gen[1617]),
			.SE(gen[1618]),

			.SELF(gen[1522]),
			.cell_state(gen[1522])
		); 

/******************* CELL 1523 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1523 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1427]),
			.N(gen[1428]),
			.NE(gen[1429]),

			.O(gen[1522]),
			.E(gen[1524]),

			.SO(gen[1617]),
			.S(gen[1618]),
			.SE(gen[1619]),

			.SELF(gen[1523]),
			.cell_state(gen[1523])
		); 

/******************* CELL 1524 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1524 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1428]),
			.N(gen[1429]),
			.NE(gen[1430]),

			.O(gen[1523]),
			.E(gen[1525]),

			.SO(gen[1618]),
			.S(gen[1619]),
			.SE(gen[1620]),

			.SELF(gen[1524]),
			.cell_state(gen[1524])
		); 

/******************* CELL 1525 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1525 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1429]),
			.N(gen[1430]),
			.NE(gen[1431]),

			.O(gen[1524]),
			.E(gen[1526]),

			.SO(gen[1619]),
			.S(gen[1620]),
			.SE(gen[1621]),

			.SELF(gen[1525]),
			.cell_state(gen[1525])
		); 

/******************* CELL 1526 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1526 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1430]),
			.N(gen[1431]),
			.NE(gen[1432]),

			.O(gen[1525]),
			.E(gen[1527]),

			.SO(gen[1620]),
			.S(gen[1621]),
			.SE(gen[1622]),

			.SELF(gen[1526]),
			.cell_state(gen[1526])
		); 

/******************* CELL 1527 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1527 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1431]),
			.N(gen[1432]),
			.NE(gen[1433]),

			.O(gen[1526]),
			.E(gen[1528]),

			.SO(gen[1621]),
			.S(gen[1622]),
			.SE(gen[1623]),

			.SELF(gen[1527]),
			.cell_state(gen[1527])
		); 

/******************* CELL 1528 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1528 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1432]),
			.N(gen[1433]),
			.NE(gen[1434]),

			.O(gen[1527]),
			.E(gen[1529]),

			.SO(gen[1622]),
			.S(gen[1623]),
			.SE(gen[1624]),

			.SELF(gen[1528]),
			.cell_state(gen[1528])
		); 

/******************* CELL 1529 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1529 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1433]),
			.N(gen[1434]),
			.NE(gen[1435]),

			.O(gen[1528]),
			.E(gen[1530]),

			.SO(gen[1623]),
			.S(gen[1624]),
			.SE(gen[1625]),

			.SELF(gen[1529]),
			.cell_state(gen[1529])
		); 

/******************* CELL 1530 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1530 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1434]),
			.N(gen[1435]),
			.NE(gen[1436]),

			.O(gen[1529]),
			.E(gen[1531]),

			.SO(gen[1624]),
			.S(gen[1625]),
			.SE(gen[1626]),

			.SELF(gen[1530]),
			.cell_state(gen[1530])
		); 

/******************* CELL 1531 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1531 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1435]),
			.N(gen[1436]),
			.NE(gen[1437]),

			.O(gen[1530]),
			.E(gen[1532]),

			.SO(gen[1625]),
			.S(gen[1626]),
			.SE(gen[1627]),

			.SELF(gen[1531]),
			.cell_state(gen[1531])
		); 

/******************* CELL 1532 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1532 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1436]),
			.N(gen[1437]),
			.NE(gen[1438]),

			.O(gen[1531]),
			.E(gen[1533]),

			.SO(gen[1626]),
			.S(gen[1627]),
			.SE(gen[1628]),

			.SELF(gen[1532]),
			.cell_state(gen[1532])
		); 

/******************* CELL 1533 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1533 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1437]),
			.N(gen[1438]),
			.NE(gen[1439]),

			.O(gen[1532]),
			.E(gen[1534]),

			.SO(gen[1627]),
			.S(gen[1628]),
			.SE(gen[1629]),

			.SELF(gen[1533]),
			.cell_state(gen[1533])
		); 

/******************* CELL 1534 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1534 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1438]),
			.N(gen[1439]),
			.NE(gen[1440]),

			.O(gen[1533]),
			.E(gen[1535]),

			.SO(gen[1628]),
			.S(gen[1629]),
			.SE(gen[1630]),

			.SELF(gen[1534]),
			.cell_state(gen[1534])
		); 

/******************* CELL 1535 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1535 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1439]),
			.N(gen[1440]),
			.NE(gen[1441]),

			.O(gen[1534]),
			.E(gen[1536]),

			.SO(gen[1629]),
			.S(gen[1630]),
			.SE(gen[1631]),

			.SELF(gen[1535]),
			.cell_state(gen[1535])
		); 

/******************* CELL 1536 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1536 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1440]),
			.N(gen[1441]),
			.NE(gen[1442]),

			.O(gen[1535]),
			.E(gen[1537]),

			.SO(gen[1630]),
			.S(gen[1631]),
			.SE(gen[1632]),

			.SELF(gen[1536]),
			.cell_state(gen[1536])
		); 

/******************* CELL 1537 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1537 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1441]),
			.N(gen[1442]),
			.NE(gen[1443]),

			.O(gen[1536]),
			.E(gen[1538]),

			.SO(gen[1631]),
			.S(gen[1632]),
			.SE(gen[1633]),

			.SELF(gen[1537]),
			.cell_state(gen[1537])
		); 

/******************* CELL 1538 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1538 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1442]),
			.N(gen[1443]),
			.NE(gen[1444]),

			.O(gen[1537]),
			.E(gen[1539]),

			.SO(gen[1632]),
			.S(gen[1633]),
			.SE(gen[1634]),

			.SELF(gen[1538]),
			.cell_state(gen[1538])
		); 

/******************* CELL 1539 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1539 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1443]),
			.N(gen[1444]),
			.NE(gen[1445]),

			.O(gen[1538]),
			.E(gen[1540]),

			.SO(gen[1633]),
			.S(gen[1634]),
			.SE(gen[1635]),

			.SELF(gen[1539]),
			.cell_state(gen[1539])
		); 

/******************* CELL 1540 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1540 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1444]),
			.N(gen[1445]),
			.NE(gen[1446]),

			.O(gen[1539]),
			.E(gen[1541]),

			.SO(gen[1634]),
			.S(gen[1635]),
			.SE(gen[1636]),

			.SELF(gen[1540]),
			.cell_state(gen[1540])
		); 

/******************* CELL 1541 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1541 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1445]),
			.N(gen[1446]),
			.NE(gen[1447]),

			.O(gen[1540]),
			.E(gen[1542]),

			.SO(gen[1635]),
			.S(gen[1636]),
			.SE(gen[1637]),

			.SELF(gen[1541]),
			.cell_state(gen[1541])
		); 

/******************* CELL 1542 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1542 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1446]),
			.N(gen[1447]),
			.NE(gen[1448]),

			.O(gen[1541]),
			.E(gen[1543]),

			.SO(gen[1636]),
			.S(gen[1637]),
			.SE(gen[1638]),

			.SELF(gen[1542]),
			.cell_state(gen[1542])
		); 

/******************* CELL 1543 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1543 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1447]),
			.N(gen[1448]),
			.NE(gen[1449]),

			.O(gen[1542]),
			.E(gen[1544]),

			.SO(gen[1637]),
			.S(gen[1638]),
			.SE(gen[1639]),

			.SELF(gen[1543]),
			.cell_state(gen[1543])
		); 

/******************* CELL 1544 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1544 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1448]),
			.N(gen[1449]),
			.NE(gen[1450]),

			.O(gen[1543]),
			.E(gen[1545]),

			.SO(gen[1638]),
			.S(gen[1639]),
			.SE(gen[1640]),

			.SELF(gen[1544]),
			.cell_state(gen[1544])
		); 

/******************* CELL 1545 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1545 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1449]),
			.N(gen[1450]),
			.NE(gen[1451]),

			.O(gen[1544]),
			.E(gen[1546]),

			.SO(gen[1639]),
			.S(gen[1640]),
			.SE(gen[1641]),

			.SELF(gen[1545]),
			.cell_state(gen[1545])
		); 

/******************* CELL 1546 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1546 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1450]),
			.N(gen[1451]),
			.NE(gen[1452]),

			.O(gen[1545]),
			.E(gen[1547]),

			.SO(gen[1640]),
			.S(gen[1641]),
			.SE(gen[1642]),

			.SELF(gen[1546]),
			.cell_state(gen[1546])
		); 

/******************* CELL 1547 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1547 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1451]),
			.N(gen[1452]),
			.NE(gen[1453]),

			.O(gen[1546]),
			.E(gen[1548]),

			.SO(gen[1641]),
			.S(gen[1642]),
			.SE(gen[1643]),

			.SELF(gen[1547]),
			.cell_state(gen[1547])
		); 

/******************* CELL 1548 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1548 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1452]),
			.N(gen[1453]),
			.NE(gen[1454]),

			.O(gen[1547]),
			.E(gen[1549]),

			.SO(gen[1642]),
			.S(gen[1643]),
			.SE(gen[1644]),

			.SELF(gen[1548]),
			.cell_state(gen[1548])
		); 

/******************* CELL 1549 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1549 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1453]),
			.N(gen[1454]),
			.NE(gen[1455]),

			.O(gen[1548]),
			.E(gen[1550]),

			.SO(gen[1643]),
			.S(gen[1644]),
			.SE(gen[1645]),

			.SELF(gen[1549]),
			.cell_state(gen[1549])
		); 

/******************* CELL 1550 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1550 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1454]),
			.N(gen[1455]),
			.NE(gen[1456]),

			.O(gen[1549]),
			.E(gen[1551]),

			.SO(gen[1644]),
			.S(gen[1645]),
			.SE(gen[1646]),

			.SELF(gen[1550]),
			.cell_state(gen[1550])
		); 

/******************* CELL 1551 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1551 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1455]),
			.N(gen[1456]),
			.NE(gen[1457]),

			.O(gen[1550]),
			.E(gen[1552]),

			.SO(gen[1645]),
			.S(gen[1646]),
			.SE(gen[1647]),

			.SELF(gen[1551]),
			.cell_state(gen[1551])
		); 

/******************* CELL 1552 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1552 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1456]),
			.N(gen[1457]),
			.NE(gen[1458]),

			.O(gen[1551]),
			.E(gen[1553]),

			.SO(gen[1646]),
			.S(gen[1647]),
			.SE(gen[1648]),

			.SELF(gen[1552]),
			.cell_state(gen[1552])
		); 

/******************* CELL 1553 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1553 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1457]),
			.N(gen[1458]),
			.NE(gen[1459]),

			.O(gen[1552]),
			.E(gen[1554]),

			.SO(gen[1647]),
			.S(gen[1648]),
			.SE(gen[1649]),

			.SELF(gen[1553]),
			.cell_state(gen[1553])
		); 

/******************* CELL 1554 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1554 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1458]),
			.N(gen[1459]),
			.NE(gen[1460]),

			.O(gen[1553]),
			.E(gen[1555]),

			.SO(gen[1648]),
			.S(gen[1649]),
			.SE(gen[1650]),

			.SELF(gen[1554]),
			.cell_state(gen[1554])
		); 

/******************* CELL 1555 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1555 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1459]),
			.N(gen[1460]),
			.NE(gen[1461]),

			.O(gen[1554]),
			.E(gen[1556]),

			.SO(gen[1649]),
			.S(gen[1650]),
			.SE(gen[1651]),

			.SELF(gen[1555]),
			.cell_state(gen[1555])
		); 

/******************* CELL 1556 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1556 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1460]),
			.N(gen[1461]),
			.NE(gen[1462]),

			.O(gen[1555]),
			.E(gen[1557]),

			.SO(gen[1650]),
			.S(gen[1651]),
			.SE(gen[1652]),

			.SELF(gen[1556]),
			.cell_state(gen[1556])
		); 

/******************* CELL 1557 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1557 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1461]),
			.N(gen[1462]),
			.NE(gen[1463]),

			.O(gen[1556]),
			.E(gen[1558]),

			.SO(gen[1651]),
			.S(gen[1652]),
			.SE(gen[1653]),

			.SELF(gen[1557]),
			.cell_state(gen[1557])
		); 

/******************* CELL 1558 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1558 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1462]),
			.N(gen[1463]),
			.NE(gen[1464]),

			.O(gen[1557]),
			.E(gen[1559]),

			.SO(gen[1652]),
			.S(gen[1653]),
			.SE(gen[1654]),

			.SELF(gen[1558]),
			.cell_state(gen[1558])
		); 

/******************* CELL 1559 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1559 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1463]),
			.N(gen[1464]),
			.NE(gen[1465]),

			.O(gen[1558]),
			.E(gen[1560]),

			.SO(gen[1653]),
			.S(gen[1654]),
			.SE(gen[1655]),

			.SELF(gen[1559]),
			.cell_state(gen[1559])
		); 

/******************* CELL 1560 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1560 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1464]),
			.N(gen[1465]),
			.NE(gen[1466]),

			.O(gen[1559]),
			.E(gen[1561]),

			.SO(gen[1654]),
			.S(gen[1655]),
			.SE(gen[1656]),

			.SELF(gen[1560]),
			.cell_state(gen[1560])
		); 

/******************* CELL 1561 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1561 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1465]),
			.N(gen[1466]),
			.NE(gen[1467]),

			.O(gen[1560]),
			.E(gen[1562]),

			.SO(gen[1655]),
			.S(gen[1656]),
			.SE(gen[1657]),

			.SELF(gen[1561]),
			.cell_state(gen[1561])
		); 

/******************* CELL 1562 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1562 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1466]),
			.N(gen[1467]),
			.NE(gen[1468]),

			.O(gen[1561]),
			.E(gen[1563]),

			.SO(gen[1656]),
			.S(gen[1657]),
			.SE(gen[1658]),

			.SELF(gen[1562]),
			.cell_state(gen[1562])
		); 

/******************* CELL 1563 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1563 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1467]),
			.N(gen[1468]),
			.NE(gen[1469]),

			.O(gen[1562]),
			.E(gen[1564]),

			.SO(gen[1657]),
			.S(gen[1658]),
			.SE(gen[1659]),

			.SELF(gen[1563]),
			.cell_state(gen[1563])
		); 

/******************* CELL 1564 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1564 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1468]),
			.N(gen[1469]),
			.NE(gen[1470]),

			.O(gen[1563]),
			.E(gen[1565]),

			.SO(gen[1658]),
			.S(gen[1659]),
			.SE(gen[1660]),

			.SELF(gen[1564]),
			.cell_state(gen[1564])
		); 

/******************* CELL 1565 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1565 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1469]),
			.N(gen[1470]),
			.NE(gen[1471]),

			.O(gen[1564]),
			.E(gen[1566]),

			.SO(gen[1659]),
			.S(gen[1660]),
			.SE(gen[1661]),

			.SELF(gen[1565]),
			.cell_state(gen[1565])
		); 

/******************* CELL 1566 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1566 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1470]),
			.N(gen[1471]),
			.NE(gen[1472]),

			.O(gen[1565]),
			.E(gen[1567]),

			.SO(gen[1660]),
			.S(gen[1661]),
			.SE(gen[1662]),

			.SELF(gen[1566]),
			.cell_state(gen[1566])
		); 

/******************* CELL 1567 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1567 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1471]),
			.N(gen[1472]),
			.NE(gen[1473]),

			.O(gen[1566]),
			.E(gen[1568]),

			.SO(gen[1661]),
			.S(gen[1662]),
			.SE(gen[1663]),

			.SELF(gen[1567]),
			.cell_state(gen[1567])
		); 

/******************* CELL 1568 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1568 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1472]),
			.N(gen[1473]),
			.NE(gen[1474]),

			.O(gen[1567]),
			.E(gen[1569]),

			.SO(gen[1662]),
			.S(gen[1663]),
			.SE(gen[1664]),

			.SELF(gen[1568]),
			.cell_state(gen[1568])
		); 

/******************* CELL 1569 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1569 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1473]),
			.N(gen[1474]),
			.NE(gen[1475]),

			.O(gen[1568]),
			.E(gen[1570]),

			.SO(gen[1663]),
			.S(gen[1664]),
			.SE(gen[1665]),

			.SELF(gen[1569]),
			.cell_state(gen[1569])
		); 

/******************* CELL 1570 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1570 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1474]),
			.N(gen[1475]),
			.NE(gen[1476]),

			.O(gen[1569]),
			.E(gen[1571]),

			.SO(gen[1664]),
			.S(gen[1665]),
			.SE(gen[1666]),

			.SELF(gen[1570]),
			.cell_state(gen[1570])
		); 

/******************* CELL 1571 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1571 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1475]),
			.N(gen[1476]),
			.NE(gen[1477]),

			.O(gen[1570]),
			.E(gen[1572]),

			.SO(gen[1665]),
			.S(gen[1666]),
			.SE(gen[1667]),

			.SELF(gen[1571]),
			.cell_state(gen[1571])
		); 

/******************* CELL 1572 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1572 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1476]),
			.N(gen[1477]),
			.NE(gen[1478]),

			.O(gen[1571]),
			.E(gen[1573]),

			.SO(gen[1666]),
			.S(gen[1667]),
			.SE(gen[1668]),

			.SELF(gen[1572]),
			.cell_state(gen[1572])
		); 

/******************* CELL 1573 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1573 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1477]),
			.N(gen[1478]),
			.NE(gen[1479]),

			.O(gen[1572]),
			.E(gen[1574]),

			.SO(gen[1667]),
			.S(gen[1668]),
			.SE(gen[1669]),

			.SELF(gen[1573]),
			.cell_state(gen[1573])
		); 

/******************* CELL 1574 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1574 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1478]),
			.N(gen[1479]),
			.NE(gen[1480]),

			.O(gen[1573]),
			.E(gen[1575]),

			.SO(gen[1668]),
			.S(gen[1669]),
			.SE(gen[1670]),

			.SELF(gen[1574]),
			.cell_state(gen[1574])
		); 

/******************* CELL 1575 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1575 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1479]),
			.N(gen[1480]),
			.NE(gen[1481]),

			.O(gen[1574]),
			.E(gen[1576]),

			.SO(gen[1669]),
			.S(gen[1670]),
			.SE(gen[1671]),

			.SELF(gen[1575]),
			.cell_state(gen[1575])
		); 

/******************* CELL 1576 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1576 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1480]),
			.N(gen[1481]),
			.NE(gen[1482]),

			.O(gen[1575]),
			.E(gen[1577]),

			.SO(gen[1670]),
			.S(gen[1671]),
			.SE(gen[1672]),

			.SELF(gen[1576]),
			.cell_state(gen[1576])
		); 

/******************* CELL 1577 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1577 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1481]),
			.N(gen[1482]),
			.NE(gen[1483]),

			.O(gen[1576]),
			.E(gen[1578]),

			.SO(gen[1671]),
			.S(gen[1672]),
			.SE(gen[1673]),

			.SELF(gen[1577]),
			.cell_state(gen[1577])
		); 

/******************* CELL 1578 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1578 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1482]),
			.N(gen[1483]),
			.NE(gen[1484]),

			.O(gen[1577]),
			.E(gen[1579]),

			.SO(gen[1672]),
			.S(gen[1673]),
			.SE(gen[1674]),

			.SELF(gen[1578]),
			.cell_state(gen[1578])
		); 

/******************* CELL 1579 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1579 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1483]),
			.N(gen[1484]),
			.NE(gen[1485]),

			.O(gen[1578]),
			.E(gen[1580]),

			.SO(gen[1673]),
			.S(gen[1674]),
			.SE(gen[1675]),

			.SELF(gen[1579]),
			.cell_state(gen[1579])
		); 

/******************* CELL 1580 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1580 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1484]),
			.N(gen[1485]),
			.NE(gen[1486]),

			.O(gen[1579]),
			.E(gen[1581]),

			.SO(gen[1674]),
			.S(gen[1675]),
			.SE(gen[1676]),

			.SELF(gen[1580]),
			.cell_state(gen[1580])
		); 

/******************* CELL 1581 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1581 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1485]),
			.N(gen[1486]),
			.NE(gen[1487]),

			.O(gen[1580]),
			.E(gen[1582]),

			.SO(gen[1675]),
			.S(gen[1676]),
			.SE(gen[1677]),

			.SELF(gen[1581]),
			.cell_state(gen[1581])
		); 

/******************* CELL 1582 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1582 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1486]),
			.N(gen[1487]),
			.NE(gen[1488]),

			.O(gen[1581]),
			.E(gen[1583]),

			.SO(gen[1676]),
			.S(gen[1677]),
			.SE(gen[1678]),

			.SELF(gen[1582]),
			.cell_state(gen[1582])
		); 

/******************* CELL 1583 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1583 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1487]),
			.N(gen[1488]),
			.NE(gen[1489]),

			.O(gen[1582]),
			.E(gen[1584]),

			.SO(gen[1677]),
			.S(gen[1678]),
			.SE(gen[1679]),

			.SELF(gen[1583]),
			.cell_state(gen[1583])
		); 

/******************* CELL 1584 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1584 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1488]),
			.N(gen[1489]),
			.NE(gen[1490]),

			.O(gen[1583]),
			.E(gen[1585]),

			.SO(gen[1678]),
			.S(gen[1679]),
			.SE(gen[1680]),

			.SELF(gen[1584]),
			.cell_state(gen[1584])
		); 

/******************* CELL 1585 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1585 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1489]),
			.N(gen[1490]),
			.NE(gen[1491]),

			.O(gen[1584]),
			.E(gen[1586]),

			.SO(gen[1679]),
			.S(gen[1680]),
			.SE(gen[1681]),

			.SELF(gen[1585]),
			.cell_state(gen[1585])
		); 

/******************* CELL 1586 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1586 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1490]),
			.N(gen[1491]),
			.NE(gen[1492]),

			.O(gen[1585]),
			.E(gen[1587]),

			.SO(gen[1680]),
			.S(gen[1681]),
			.SE(gen[1682]),

			.SELF(gen[1586]),
			.cell_state(gen[1586])
		); 

/******************* CELL 1587 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1587 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1491]),
			.N(gen[1492]),
			.NE(gen[1493]),

			.O(gen[1586]),
			.E(gen[1588]),

			.SO(gen[1681]),
			.S(gen[1682]),
			.SE(gen[1683]),

			.SELF(gen[1587]),
			.cell_state(gen[1587])
		); 

/******************* CELL 1588 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1588 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1492]),
			.N(gen[1493]),
			.NE(gen[1494]),

			.O(gen[1587]),
			.E(gen[1589]),

			.SO(gen[1682]),
			.S(gen[1683]),
			.SE(gen[1684]),

			.SELF(gen[1588]),
			.cell_state(gen[1588])
		); 

/******************* CELL 1589 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1589 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1493]),
			.N(gen[1494]),
			.NE(gen[1495]),

			.O(gen[1588]),
			.E(gen[1590]),

			.SO(gen[1683]),
			.S(gen[1684]),
			.SE(gen[1685]),

			.SELF(gen[1589]),
			.cell_state(gen[1589])
		); 

/******************* CELL 1590 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1590 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1494]),
			.N(gen[1495]),
			.NE(gen[1496]),

			.O(gen[1589]),
			.E(gen[1591]),

			.SO(gen[1684]),
			.S(gen[1685]),
			.SE(gen[1686]),

			.SELF(gen[1590]),
			.cell_state(gen[1590])
		); 

/******************* CELL 1591 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1591 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1495]),
			.N(gen[1496]),
			.NE(gen[1497]),

			.O(gen[1590]),
			.E(gen[1592]),

			.SO(gen[1685]),
			.S(gen[1686]),
			.SE(gen[1687]),

			.SELF(gen[1591]),
			.cell_state(gen[1591])
		); 

/******************* CELL 1592 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1592 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1496]),
			.N(gen[1497]),
			.NE(gen[1498]),

			.O(gen[1591]),
			.E(gen[1593]),

			.SO(gen[1686]),
			.S(gen[1687]),
			.SE(gen[1688]),

			.SELF(gen[1592]),
			.cell_state(gen[1592])
		); 

/******************* CELL 1593 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1593 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1497]),
			.N(gen[1498]),
			.NE(gen[1499]),

			.O(gen[1592]),
			.E(gen[1594]),

			.SO(gen[1687]),
			.S(gen[1688]),
			.SE(gen[1689]),

			.SELF(gen[1593]),
			.cell_state(gen[1593])
		); 

/******************* CELL 1594 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1594 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1498]),
			.N(gen[1499]),
			.NE(gen[1500]),

			.O(gen[1593]),
			.E(gen[1595]),

			.SO(gen[1688]),
			.S(gen[1689]),
			.SE(gen[1690]),

			.SELF(gen[1594]),
			.cell_state(gen[1594])
		); 

/******************* CELL 1595 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1595 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1499]),
			.N(gen[1500]),
			.NE(gen[1501]),

			.O(gen[1594]),
			.E(gen[1596]),

			.SO(gen[1689]),
			.S(gen[1690]),
			.SE(gen[1691]),

			.SELF(gen[1595]),
			.cell_state(gen[1595])
		); 

/******************* CELL 1596 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1596 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1500]),
			.N(gen[1501]),
			.NE(gen[1502]),

			.O(gen[1595]),
			.E(gen[1597]),

			.SO(gen[1690]),
			.S(gen[1691]),
			.SE(gen[1692]),

			.SELF(gen[1596]),
			.cell_state(gen[1596])
		); 

/******************* CELL 1597 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1597 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1501]),
			.N(gen[1502]),
			.NE(gen[1503]),

			.O(gen[1596]),
			.E(gen[1598]),

			.SO(gen[1691]),
			.S(gen[1692]),
			.SE(gen[1693]),

			.SELF(gen[1597]),
			.cell_state(gen[1597])
		); 

/******************* CELL 1598 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1598 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1502]),
			.N(gen[1503]),
			.NE(gen[1504]),

			.O(gen[1597]),
			.E(gen[1599]),

			.SO(gen[1692]),
			.S(gen[1693]),
			.SE(gen[1694]),

			.SELF(gen[1598]),
			.cell_state(gen[1598])
		); 

/******************* CELL 1599 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1599 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1503]),
			.N(gen[1504]),
			.NE(gen[1505]),

			.O(gen[1598]),
			.E(gen[1600]),

			.SO(gen[1693]),
			.S(gen[1694]),
			.SE(gen[1695]),

			.SELF(gen[1599]),
			.cell_state(gen[1599])
		); 

/******************* CELL 1600 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1600 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1504]),
			.N(gen[1505]),
			.NE(gen[1506]),

			.O(gen[1599]),
			.E(gen[1601]),

			.SO(gen[1694]),
			.S(gen[1695]),
			.SE(gen[1696]),

			.SELF(gen[1600]),
			.cell_state(gen[1600])
		); 

/******************* CELL 1601 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1601 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1505]),
			.N(gen[1506]),
			.NE(gen[1507]),

			.O(gen[1600]),
			.E(gen[1602]),

			.SO(gen[1695]),
			.S(gen[1696]),
			.SE(gen[1697]),

			.SELF(gen[1601]),
			.cell_state(gen[1601])
		); 

/******************* CELL 1602 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1602 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1506]),
			.N(gen[1507]),
			.NE(gen[1508]),

			.O(gen[1601]),
			.E(gen[1603]),

			.SO(gen[1696]),
			.S(gen[1697]),
			.SE(gen[1698]),

			.SELF(gen[1602]),
			.cell_state(gen[1602])
		); 

/******************* CELL 1603 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1603 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1507]),
			.N(gen[1508]),
			.NE(gen[1509]),

			.O(gen[1602]),
			.E(gen[1604]),

			.SO(gen[1697]),
			.S(gen[1698]),
			.SE(gen[1699]),

			.SELF(gen[1603]),
			.cell_state(gen[1603])
		); 

/******************* CELL 1604 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1604 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1508]),
			.N(gen[1509]),
			.NE(gen[1510]),

			.O(gen[1603]),
			.E(gen[1605]),

			.SO(gen[1698]),
			.S(gen[1699]),
			.SE(gen[1700]),

			.SELF(gen[1604]),
			.cell_state(gen[1604])
		); 

/******************* CELL 1605 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1605 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1509]),
			.N(gen[1510]),
			.NE(gen[1511]),

			.O(gen[1604]),
			.E(gen[1606]),

			.SO(gen[1699]),
			.S(gen[1700]),
			.SE(gen[1701]),

			.SELF(gen[1605]),
			.cell_state(gen[1605])
		); 

/******************* CELL 1606 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1606 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1510]),
			.N(gen[1511]),
			.NE(gen[1512]),

			.O(gen[1605]),
			.E(gen[1607]),

			.SO(gen[1700]),
			.S(gen[1701]),
			.SE(gen[1702]),

			.SELF(gen[1606]),
			.cell_state(gen[1606])
		); 

/******************* CELL 1607 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1607 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1511]),
			.N(gen[1512]),
			.NE(gen[1513]),

			.O(gen[1606]),
			.E(gen[1608]),

			.SO(gen[1701]),
			.S(gen[1702]),
			.SE(gen[1703]),

			.SELF(gen[1607]),
			.cell_state(gen[1607])
		); 

/******************* CELL 1608 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1608 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1512]),
			.N(gen[1513]),
			.NE(gen[1514]),

			.O(gen[1607]),
			.E(gen[1609]),

			.SO(gen[1702]),
			.S(gen[1703]),
			.SE(gen[1704]),

			.SELF(gen[1608]),
			.cell_state(gen[1608])
		); 

/******************* CELL 1609 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1609 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1513]),
			.N(gen[1514]),
			.NE(gen[1515]),

			.O(gen[1608]),
			.E(gen[1610]),

			.SO(gen[1703]),
			.S(gen[1704]),
			.SE(gen[1705]),

			.SELF(gen[1609]),
			.cell_state(gen[1609])
		); 

/******************* CELL 1610 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1610 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1514]),
			.N(gen[1515]),
			.NE(gen[1516]),

			.O(gen[1609]),
			.E(gen[1611]),

			.SO(gen[1704]),
			.S(gen[1705]),
			.SE(gen[1706]),

			.SELF(gen[1610]),
			.cell_state(gen[1610])
		); 

/******************* CELL 1611 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1611 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1515]),
			.N(gen[1516]),
			.NE(gen[1517]),

			.O(gen[1610]),
			.E(gen[1612]),

			.SO(gen[1705]),
			.S(gen[1706]),
			.SE(gen[1707]),

			.SELF(gen[1611]),
			.cell_state(gen[1611])
		); 

/******************* CELL 1612 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1612 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1516]),
			.N(gen[1517]),
			.NE(gen[1518]),

			.O(gen[1611]),
			.E(gen[1613]),

			.SO(gen[1706]),
			.S(gen[1707]),
			.SE(gen[1708]),

			.SELF(gen[1612]),
			.cell_state(gen[1612])
		); 

/******************* CELL 1613 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1613 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1517]),
			.N(gen[1518]),
			.NE(gen[1519]),

			.O(gen[1612]),
			.E(gen[1614]),

			.SO(gen[1707]),
			.S(gen[1708]),
			.SE(gen[1709]),

			.SELF(gen[1613]),
			.cell_state(gen[1613])
		); 

/******************* CELL 1614 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1614 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1518]),
			.N(gen[1519]),
			.NE(gen[1518]),

			.O(gen[1613]),
			.E(gen[1613]),

			.SO(gen[1708]),
			.S(gen[1709]),
			.SE(gen[1708]),

			.SELF(gen[1614]),
			.cell_state(gen[1614])
		); 

/******************* CELL 1615 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1615 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1521]),
			.N(gen[1520]),
			.NE(gen[1521]),

			.O(gen[1616]),
			.E(gen[1616]),

			.SO(gen[1711]),
			.S(gen[1710]),
			.SE(gen[1711]),

			.SELF(gen[1615]),
			.cell_state(gen[1615])
		); 

/******************* CELL 1616 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1616 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1520]),
			.N(gen[1521]),
			.NE(gen[1522]),

			.O(gen[1615]),
			.E(gen[1617]),

			.SO(gen[1710]),
			.S(gen[1711]),
			.SE(gen[1712]),

			.SELF(gen[1616]),
			.cell_state(gen[1616])
		); 

/******************* CELL 1617 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1617 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1521]),
			.N(gen[1522]),
			.NE(gen[1523]),

			.O(gen[1616]),
			.E(gen[1618]),

			.SO(gen[1711]),
			.S(gen[1712]),
			.SE(gen[1713]),

			.SELF(gen[1617]),
			.cell_state(gen[1617])
		); 

/******************* CELL 1618 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1618 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1522]),
			.N(gen[1523]),
			.NE(gen[1524]),

			.O(gen[1617]),
			.E(gen[1619]),

			.SO(gen[1712]),
			.S(gen[1713]),
			.SE(gen[1714]),

			.SELF(gen[1618]),
			.cell_state(gen[1618])
		); 

/******************* CELL 1619 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1619 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1523]),
			.N(gen[1524]),
			.NE(gen[1525]),

			.O(gen[1618]),
			.E(gen[1620]),

			.SO(gen[1713]),
			.S(gen[1714]),
			.SE(gen[1715]),

			.SELF(gen[1619]),
			.cell_state(gen[1619])
		); 

/******************* CELL 1620 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1620 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1524]),
			.N(gen[1525]),
			.NE(gen[1526]),

			.O(gen[1619]),
			.E(gen[1621]),

			.SO(gen[1714]),
			.S(gen[1715]),
			.SE(gen[1716]),

			.SELF(gen[1620]),
			.cell_state(gen[1620])
		); 

/******************* CELL 1621 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1621 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1525]),
			.N(gen[1526]),
			.NE(gen[1527]),

			.O(gen[1620]),
			.E(gen[1622]),

			.SO(gen[1715]),
			.S(gen[1716]),
			.SE(gen[1717]),

			.SELF(gen[1621]),
			.cell_state(gen[1621])
		); 

/******************* CELL 1622 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1622 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1526]),
			.N(gen[1527]),
			.NE(gen[1528]),

			.O(gen[1621]),
			.E(gen[1623]),

			.SO(gen[1716]),
			.S(gen[1717]),
			.SE(gen[1718]),

			.SELF(gen[1622]),
			.cell_state(gen[1622])
		); 

/******************* CELL 1623 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1623 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1527]),
			.N(gen[1528]),
			.NE(gen[1529]),

			.O(gen[1622]),
			.E(gen[1624]),

			.SO(gen[1717]),
			.S(gen[1718]),
			.SE(gen[1719]),

			.SELF(gen[1623]),
			.cell_state(gen[1623])
		); 

/******************* CELL 1624 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1624 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1528]),
			.N(gen[1529]),
			.NE(gen[1530]),

			.O(gen[1623]),
			.E(gen[1625]),

			.SO(gen[1718]),
			.S(gen[1719]),
			.SE(gen[1720]),

			.SELF(gen[1624]),
			.cell_state(gen[1624])
		); 

/******************* CELL 1625 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1625 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1529]),
			.N(gen[1530]),
			.NE(gen[1531]),

			.O(gen[1624]),
			.E(gen[1626]),

			.SO(gen[1719]),
			.S(gen[1720]),
			.SE(gen[1721]),

			.SELF(gen[1625]),
			.cell_state(gen[1625])
		); 

/******************* CELL 1626 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1626 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1530]),
			.N(gen[1531]),
			.NE(gen[1532]),

			.O(gen[1625]),
			.E(gen[1627]),

			.SO(gen[1720]),
			.S(gen[1721]),
			.SE(gen[1722]),

			.SELF(gen[1626]),
			.cell_state(gen[1626])
		); 

/******************* CELL 1627 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1627 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1531]),
			.N(gen[1532]),
			.NE(gen[1533]),

			.O(gen[1626]),
			.E(gen[1628]),

			.SO(gen[1721]),
			.S(gen[1722]),
			.SE(gen[1723]),

			.SELF(gen[1627]),
			.cell_state(gen[1627])
		); 

/******************* CELL 1628 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1628 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1532]),
			.N(gen[1533]),
			.NE(gen[1534]),

			.O(gen[1627]),
			.E(gen[1629]),

			.SO(gen[1722]),
			.S(gen[1723]),
			.SE(gen[1724]),

			.SELF(gen[1628]),
			.cell_state(gen[1628])
		); 

/******************* CELL 1629 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1629 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1533]),
			.N(gen[1534]),
			.NE(gen[1535]),

			.O(gen[1628]),
			.E(gen[1630]),

			.SO(gen[1723]),
			.S(gen[1724]),
			.SE(gen[1725]),

			.SELF(gen[1629]),
			.cell_state(gen[1629])
		); 

/******************* CELL 1630 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1630 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1534]),
			.N(gen[1535]),
			.NE(gen[1536]),

			.O(gen[1629]),
			.E(gen[1631]),

			.SO(gen[1724]),
			.S(gen[1725]),
			.SE(gen[1726]),

			.SELF(gen[1630]),
			.cell_state(gen[1630])
		); 

/******************* CELL 1631 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1631 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1535]),
			.N(gen[1536]),
			.NE(gen[1537]),

			.O(gen[1630]),
			.E(gen[1632]),

			.SO(gen[1725]),
			.S(gen[1726]),
			.SE(gen[1727]),

			.SELF(gen[1631]),
			.cell_state(gen[1631])
		); 

/******************* CELL 1632 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1632 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1536]),
			.N(gen[1537]),
			.NE(gen[1538]),

			.O(gen[1631]),
			.E(gen[1633]),

			.SO(gen[1726]),
			.S(gen[1727]),
			.SE(gen[1728]),

			.SELF(gen[1632]),
			.cell_state(gen[1632])
		); 

/******************* CELL 1633 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1633 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1537]),
			.N(gen[1538]),
			.NE(gen[1539]),

			.O(gen[1632]),
			.E(gen[1634]),

			.SO(gen[1727]),
			.S(gen[1728]),
			.SE(gen[1729]),

			.SELF(gen[1633]),
			.cell_state(gen[1633])
		); 

/******************* CELL 1634 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1634 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1538]),
			.N(gen[1539]),
			.NE(gen[1540]),

			.O(gen[1633]),
			.E(gen[1635]),

			.SO(gen[1728]),
			.S(gen[1729]),
			.SE(gen[1730]),

			.SELF(gen[1634]),
			.cell_state(gen[1634])
		); 

/******************* CELL 1635 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1635 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1539]),
			.N(gen[1540]),
			.NE(gen[1541]),

			.O(gen[1634]),
			.E(gen[1636]),

			.SO(gen[1729]),
			.S(gen[1730]),
			.SE(gen[1731]),

			.SELF(gen[1635]),
			.cell_state(gen[1635])
		); 

/******************* CELL 1636 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1636 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1540]),
			.N(gen[1541]),
			.NE(gen[1542]),

			.O(gen[1635]),
			.E(gen[1637]),

			.SO(gen[1730]),
			.S(gen[1731]),
			.SE(gen[1732]),

			.SELF(gen[1636]),
			.cell_state(gen[1636])
		); 

/******************* CELL 1637 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1637 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1541]),
			.N(gen[1542]),
			.NE(gen[1543]),

			.O(gen[1636]),
			.E(gen[1638]),

			.SO(gen[1731]),
			.S(gen[1732]),
			.SE(gen[1733]),

			.SELF(gen[1637]),
			.cell_state(gen[1637])
		); 

/******************* CELL 1638 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1638 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1542]),
			.N(gen[1543]),
			.NE(gen[1544]),

			.O(gen[1637]),
			.E(gen[1639]),

			.SO(gen[1732]),
			.S(gen[1733]),
			.SE(gen[1734]),

			.SELF(gen[1638]),
			.cell_state(gen[1638])
		); 

/******************* CELL 1639 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1639 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1543]),
			.N(gen[1544]),
			.NE(gen[1545]),

			.O(gen[1638]),
			.E(gen[1640]),

			.SO(gen[1733]),
			.S(gen[1734]),
			.SE(gen[1735]),

			.SELF(gen[1639]),
			.cell_state(gen[1639])
		); 

/******************* CELL 1640 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1640 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1544]),
			.N(gen[1545]),
			.NE(gen[1546]),

			.O(gen[1639]),
			.E(gen[1641]),

			.SO(gen[1734]),
			.S(gen[1735]),
			.SE(gen[1736]),

			.SELF(gen[1640]),
			.cell_state(gen[1640])
		); 

/******************* CELL 1641 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1641 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1545]),
			.N(gen[1546]),
			.NE(gen[1547]),

			.O(gen[1640]),
			.E(gen[1642]),

			.SO(gen[1735]),
			.S(gen[1736]),
			.SE(gen[1737]),

			.SELF(gen[1641]),
			.cell_state(gen[1641])
		); 

/******************* CELL 1642 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1642 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1546]),
			.N(gen[1547]),
			.NE(gen[1548]),

			.O(gen[1641]),
			.E(gen[1643]),

			.SO(gen[1736]),
			.S(gen[1737]),
			.SE(gen[1738]),

			.SELF(gen[1642]),
			.cell_state(gen[1642])
		); 

/******************* CELL 1643 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1643 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1547]),
			.N(gen[1548]),
			.NE(gen[1549]),

			.O(gen[1642]),
			.E(gen[1644]),

			.SO(gen[1737]),
			.S(gen[1738]),
			.SE(gen[1739]),

			.SELF(gen[1643]),
			.cell_state(gen[1643])
		); 

/******************* CELL 1644 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1644 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1548]),
			.N(gen[1549]),
			.NE(gen[1550]),

			.O(gen[1643]),
			.E(gen[1645]),

			.SO(gen[1738]),
			.S(gen[1739]),
			.SE(gen[1740]),

			.SELF(gen[1644]),
			.cell_state(gen[1644])
		); 

/******************* CELL 1645 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1645 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1549]),
			.N(gen[1550]),
			.NE(gen[1551]),

			.O(gen[1644]),
			.E(gen[1646]),

			.SO(gen[1739]),
			.S(gen[1740]),
			.SE(gen[1741]),

			.SELF(gen[1645]),
			.cell_state(gen[1645])
		); 

/******************* CELL 1646 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1646 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1550]),
			.N(gen[1551]),
			.NE(gen[1552]),

			.O(gen[1645]),
			.E(gen[1647]),

			.SO(gen[1740]),
			.S(gen[1741]),
			.SE(gen[1742]),

			.SELF(gen[1646]),
			.cell_state(gen[1646])
		); 

/******************* CELL 1647 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1647 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1551]),
			.N(gen[1552]),
			.NE(gen[1553]),

			.O(gen[1646]),
			.E(gen[1648]),

			.SO(gen[1741]),
			.S(gen[1742]),
			.SE(gen[1743]),

			.SELF(gen[1647]),
			.cell_state(gen[1647])
		); 

/******************* CELL 1648 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1648 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1552]),
			.N(gen[1553]),
			.NE(gen[1554]),

			.O(gen[1647]),
			.E(gen[1649]),

			.SO(gen[1742]),
			.S(gen[1743]),
			.SE(gen[1744]),

			.SELF(gen[1648]),
			.cell_state(gen[1648])
		); 

/******************* CELL 1649 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1649 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1553]),
			.N(gen[1554]),
			.NE(gen[1555]),

			.O(gen[1648]),
			.E(gen[1650]),

			.SO(gen[1743]),
			.S(gen[1744]),
			.SE(gen[1745]),

			.SELF(gen[1649]),
			.cell_state(gen[1649])
		); 

/******************* CELL 1650 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1650 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1554]),
			.N(gen[1555]),
			.NE(gen[1556]),

			.O(gen[1649]),
			.E(gen[1651]),

			.SO(gen[1744]),
			.S(gen[1745]),
			.SE(gen[1746]),

			.SELF(gen[1650]),
			.cell_state(gen[1650])
		); 

/******************* CELL 1651 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1651 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1555]),
			.N(gen[1556]),
			.NE(gen[1557]),

			.O(gen[1650]),
			.E(gen[1652]),

			.SO(gen[1745]),
			.S(gen[1746]),
			.SE(gen[1747]),

			.SELF(gen[1651]),
			.cell_state(gen[1651])
		); 

/******************* CELL 1652 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1652 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1556]),
			.N(gen[1557]),
			.NE(gen[1558]),

			.O(gen[1651]),
			.E(gen[1653]),

			.SO(gen[1746]),
			.S(gen[1747]),
			.SE(gen[1748]),

			.SELF(gen[1652]),
			.cell_state(gen[1652])
		); 

/******************* CELL 1653 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1653 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1557]),
			.N(gen[1558]),
			.NE(gen[1559]),

			.O(gen[1652]),
			.E(gen[1654]),

			.SO(gen[1747]),
			.S(gen[1748]),
			.SE(gen[1749]),

			.SELF(gen[1653]),
			.cell_state(gen[1653])
		); 

/******************* CELL 1654 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1654 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1558]),
			.N(gen[1559]),
			.NE(gen[1560]),

			.O(gen[1653]),
			.E(gen[1655]),

			.SO(gen[1748]),
			.S(gen[1749]),
			.SE(gen[1750]),

			.SELF(gen[1654]),
			.cell_state(gen[1654])
		); 

/******************* CELL 1655 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1655 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1559]),
			.N(gen[1560]),
			.NE(gen[1561]),

			.O(gen[1654]),
			.E(gen[1656]),

			.SO(gen[1749]),
			.S(gen[1750]),
			.SE(gen[1751]),

			.SELF(gen[1655]),
			.cell_state(gen[1655])
		); 

/******************* CELL 1656 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1656 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1560]),
			.N(gen[1561]),
			.NE(gen[1562]),

			.O(gen[1655]),
			.E(gen[1657]),

			.SO(gen[1750]),
			.S(gen[1751]),
			.SE(gen[1752]),

			.SELF(gen[1656]),
			.cell_state(gen[1656])
		); 

/******************* CELL 1657 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1657 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1561]),
			.N(gen[1562]),
			.NE(gen[1563]),

			.O(gen[1656]),
			.E(gen[1658]),

			.SO(gen[1751]),
			.S(gen[1752]),
			.SE(gen[1753]),

			.SELF(gen[1657]),
			.cell_state(gen[1657])
		); 

/******************* CELL 1658 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1658 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1562]),
			.N(gen[1563]),
			.NE(gen[1564]),

			.O(gen[1657]),
			.E(gen[1659]),

			.SO(gen[1752]),
			.S(gen[1753]),
			.SE(gen[1754]),

			.SELF(gen[1658]),
			.cell_state(gen[1658])
		); 

/******************* CELL 1659 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1659 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1563]),
			.N(gen[1564]),
			.NE(gen[1565]),

			.O(gen[1658]),
			.E(gen[1660]),

			.SO(gen[1753]),
			.S(gen[1754]),
			.SE(gen[1755]),

			.SELF(gen[1659]),
			.cell_state(gen[1659])
		); 

/******************* CELL 1660 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1660 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1564]),
			.N(gen[1565]),
			.NE(gen[1566]),

			.O(gen[1659]),
			.E(gen[1661]),

			.SO(gen[1754]),
			.S(gen[1755]),
			.SE(gen[1756]),

			.SELF(gen[1660]),
			.cell_state(gen[1660])
		); 

/******************* CELL 1661 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1661 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1565]),
			.N(gen[1566]),
			.NE(gen[1567]),

			.O(gen[1660]),
			.E(gen[1662]),

			.SO(gen[1755]),
			.S(gen[1756]),
			.SE(gen[1757]),

			.SELF(gen[1661]),
			.cell_state(gen[1661])
		); 

/******************* CELL 1662 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1662 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1566]),
			.N(gen[1567]),
			.NE(gen[1568]),

			.O(gen[1661]),
			.E(gen[1663]),

			.SO(gen[1756]),
			.S(gen[1757]),
			.SE(gen[1758]),

			.SELF(gen[1662]),
			.cell_state(gen[1662])
		); 

/******************* CELL 1663 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1663 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1567]),
			.N(gen[1568]),
			.NE(gen[1569]),

			.O(gen[1662]),
			.E(gen[1664]),

			.SO(gen[1757]),
			.S(gen[1758]),
			.SE(gen[1759]),

			.SELF(gen[1663]),
			.cell_state(gen[1663])
		); 

/******************* CELL 1664 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1664 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1568]),
			.N(gen[1569]),
			.NE(gen[1570]),

			.O(gen[1663]),
			.E(gen[1665]),

			.SO(gen[1758]),
			.S(gen[1759]),
			.SE(gen[1760]),

			.SELF(gen[1664]),
			.cell_state(gen[1664])
		); 

/******************* CELL 1665 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1665 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1569]),
			.N(gen[1570]),
			.NE(gen[1571]),

			.O(gen[1664]),
			.E(gen[1666]),

			.SO(gen[1759]),
			.S(gen[1760]),
			.SE(gen[1761]),

			.SELF(gen[1665]),
			.cell_state(gen[1665])
		); 

/******************* CELL 1666 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1666 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1570]),
			.N(gen[1571]),
			.NE(gen[1572]),

			.O(gen[1665]),
			.E(gen[1667]),

			.SO(gen[1760]),
			.S(gen[1761]),
			.SE(gen[1762]),

			.SELF(gen[1666]),
			.cell_state(gen[1666])
		); 

/******************* CELL 1667 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1667 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1571]),
			.N(gen[1572]),
			.NE(gen[1573]),

			.O(gen[1666]),
			.E(gen[1668]),

			.SO(gen[1761]),
			.S(gen[1762]),
			.SE(gen[1763]),

			.SELF(gen[1667]),
			.cell_state(gen[1667])
		); 

/******************* CELL 1668 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1668 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1572]),
			.N(gen[1573]),
			.NE(gen[1574]),

			.O(gen[1667]),
			.E(gen[1669]),

			.SO(gen[1762]),
			.S(gen[1763]),
			.SE(gen[1764]),

			.SELF(gen[1668]),
			.cell_state(gen[1668])
		); 

/******************* CELL 1669 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1669 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1573]),
			.N(gen[1574]),
			.NE(gen[1575]),

			.O(gen[1668]),
			.E(gen[1670]),

			.SO(gen[1763]),
			.S(gen[1764]),
			.SE(gen[1765]),

			.SELF(gen[1669]),
			.cell_state(gen[1669])
		); 

/******************* CELL 1670 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1670 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1574]),
			.N(gen[1575]),
			.NE(gen[1576]),

			.O(gen[1669]),
			.E(gen[1671]),

			.SO(gen[1764]),
			.S(gen[1765]),
			.SE(gen[1766]),

			.SELF(gen[1670]),
			.cell_state(gen[1670])
		); 

/******************* CELL 1671 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1671 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1575]),
			.N(gen[1576]),
			.NE(gen[1577]),

			.O(gen[1670]),
			.E(gen[1672]),

			.SO(gen[1765]),
			.S(gen[1766]),
			.SE(gen[1767]),

			.SELF(gen[1671]),
			.cell_state(gen[1671])
		); 

/******************* CELL 1672 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1672 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1576]),
			.N(gen[1577]),
			.NE(gen[1578]),

			.O(gen[1671]),
			.E(gen[1673]),

			.SO(gen[1766]),
			.S(gen[1767]),
			.SE(gen[1768]),

			.SELF(gen[1672]),
			.cell_state(gen[1672])
		); 

/******************* CELL 1673 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1673 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1577]),
			.N(gen[1578]),
			.NE(gen[1579]),

			.O(gen[1672]),
			.E(gen[1674]),

			.SO(gen[1767]),
			.S(gen[1768]),
			.SE(gen[1769]),

			.SELF(gen[1673]),
			.cell_state(gen[1673])
		); 

/******************* CELL 1674 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1674 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1578]),
			.N(gen[1579]),
			.NE(gen[1580]),

			.O(gen[1673]),
			.E(gen[1675]),

			.SO(gen[1768]),
			.S(gen[1769]),
			.SE(gen[1770]),

			.SELF(gen[1674]),
			.cell_state(gen[1674])
		); 

/******************* CELL 1675 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1675 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1579]),
			.N(gen[1580]),
			.NE(gen[1581]),

			.O(gen[1674]),
			.E(gen[1676]),

			.SO(gen[1769]),
			.S(gen[1770]),
			.SE(gen[1771]),

			.SELF(gen[1675]),
			.cell_state(gen[1675])
		); 

/******************* CELL 1676 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1676 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1580]),
			.N(gen[1581]),
			.NE(gen[1582]),

			.O(gen[1675]),
			.E(gen[1677]),

			.SO(gen[1770]),
			.S(gen[1771]),
			.SE(gen[1772]),

			.SELF(gen[1676]),
			.cell_state(gen[1676])
		); 

/******************* CELL 1677 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1677 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1581]),
			.N(gen[1582]),
			.NE(gen[1583]),

			.O(gen[1676]),
			.E(gen[1678]),

			.SO(gen[1771]),
			.S(gen[1772]),
			.SE(gen[1773]),

			.SELF(gen[1677]),
			.cell_state(gen[1677])
		); 

/******************* CELL 1678 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1678 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1582]),
			.N(gen[1583]),
			.NE(gen[1584]),

			.O(gen[1677]),
			.E(gen[1679]),

			.SO(gen[1772]),
			.S(gen[1773]),
			.SE(gen[1774]),

			.SELF(gen[1678]),
			.cell_state(gen[1678])
		); 

/******************* CELL 1679 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1679 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1583]),
			.N(gen[1584]),
			.NE(gen[1585]),

			.O(gen[1678]),
			.E(gen[1680]),

			.SO(gen[1773]),
			.S(gen[1774]),
			.SE(gen[1775]),

			.SELF(gen[1679]),
			.cell_state(gen[1679])
		); 

/******************* CELL 1680 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1680 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1584]),
			.N(gen[1585]),
			.NE(gen[1586]),

			.O(gen[1679]),
			.E(gen[1681]),

			.SO(gen[1774]),
			.S(gen[1775]),
			.SE(gen[1776]),

			.SELF(gen[1680]),
			.cell_state(gen[1680])
		); 

/******************* CELL 1681 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1681 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1585]),
			.N(gen[1586]),
			.NE(gen[1587]),

			.O(gen[1680]),
			.E(gen[1682]),

			.SO(gen[1775]),
			.S(gen[1776]),
			.SE(gen[1777]),

			.SELF(gen[1681]),
			.cell_state(gen[1681])
		); 

/******************* CELL 1682 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1682 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1586]),
			.N(gen[1587]),
			.NE(gen[1588]),

			.O(gen[1681]),
			.E(gen[1683]),

			.SO(gen[1776]),
			.S(gen[1777]),
			.SE(gen[1778]),

			.SELF(gen[1682]),
			.cell_state(gen[1682])
		); 

/******************* CELL 1683 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1683 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1587]),
			.N(gen[1588]),
			.NE(gen[1589]),

			.O(gen[1682]),
			.E(gen[1684]),

			.SO(gen[1777]),
			.S(gen[1778]),
			.SE(gen[1779]),

			.SELF(gen[1683]),
			.cell_state(gen[1683])
		); 

/******************* CELL 1684 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1684 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1588]),
			.N(gen[1589]),
			.NE(gen[1590]),

			.O(gen[1683]),
			.E(gen[1685]),

			.SO(gen[1778]),
			.S(gen[1779]),
			.SE(gen[1780]),

			.SELF(gen[1684]),
			.cell_state(gen[1684])
		); 

/******************* CELL 1685 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1685 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1589]),
			.N(gen[1590]),
			.NE(gen[1591]),

			.O(gen[1684]),
			.E(gen[1686]),

			.SO(gen[1779]),
			.S(gen[1780]),
			.SE(gen[1781]),

			.SELF(gen[1685]),
			.cell_state(gen[1685])
		); 

/******************* CELL 1686 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1686 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1590]),
			.N(gen[1591]),
			.NE(gen[1592]),

			.O(gen[1685]),
			.E(gen[1687]),

			.SO(gen[1780]),
			.S(gen[1781]),
			.SE(gen[1782]),

			.SELF(gen[1686]),
			.cell_state(gen[1686])
		); 

/******************* CELL 1687 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1687 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1591]),
			.N(gen[1592]),
			.NE(gen[1593]),

			.O(gen[1686]),
			.E(gen[1688]),

			.SO(gen[1781]),
			.S(gen[1782]),
			.SE(gen[1783]),

			.SELF(gen[1687]),
			.cell_state(gen[1687])
		); 

/******************* CELL 1688 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1688 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1592]),
			.N(gen[1593]),
			.NE(gen[1594]),

			.O(gen[1687]),
			.E(gen[1689]),

			.SO(gen[1782]),
			.S(gen[1783]),
			.SE(gen[1784]),

			.SELF(gen[1688]),
			.cell_state(gen[1688])
		); 

/******************* CELL 1689 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1689 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1593]),
			.N(gen[1594]),
			.NE(gen[1595]),

			.O(gen[1688]),
			.E(gen[1690]),

			.SO(gen[1783]),
			.S(gen[1784]),
			.SE(gen[1785]),

			.SELF(gen[1689]),
			.cell_state(gen[1689])
		); 

/******************* CELL 1690 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1690 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1594]),
			.N(gen[1595]),
			.NE(gen[1596]),

			.O(gen[1689]),
			.E(gen[1691]),

			.SO(gen[1784]),
			.S(gen[1785]),
			.SE(gen[1786]),

			.SELF(gen[1690]),
			.cell_state(gen[1690])
		); 

/******************* CELL 1691 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1691 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1595]),
			.N(gen[1596]),
			.NE(gen[1597]),

			.O(gen[1690]),
			.E(gen[1692]),

			.SO(gen[1785]),
			.S(gen[1786]),
			.SE(gen[1787]),

			.SELF(gen[1691]),
			.cell_state(gen[1691])
		); 

/******************* CELL 1692 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1692 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1596]),
			.N(gen[1597]),
			.NE(gen[1598]),

			.O(gen[1691]),
			.E(gen[1693]),

			.SO(gen[1786]),
			.S(gen[1787]),
			.SE(gen[1788]),

			.SELF(gen[1692]),
			.cell_state(gen[1692])
		); 

/******************* CELL 1693 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1693 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1597]),
			.N(gen[1598]),
			.NE(gen[1599]),

			.O(gen[1692]),
			.E(gen[1694]),

			.SO(gen[1787]),
			.S(gen[1788]),
			.SE(gen[1789]),

			.SELF(gen[1693]),
			.cell_state(gen[1693])
		); 

/******************* CELL 1694 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1694 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1598]),
			.N(gen[1599]),
			.NE(gen[1600]),

			.O(gen[1693]),
			.E(gen[1695]),

			.SO(gen[1788]),
			.S(gen[1789]),
			.SE(gen[1790]),

			.SELF(gen[1694]),
			.cell_state(gen[1694])
		); 

/******************* CELL 1695 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1695 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1599]),
			.N(gen[1600]),
			.NE(gen[1601]),

			.O(gen[1694]),
			.E(gen[1696]),

			.SO(gen[1789]),
			.S(gen[1790]),
			.SE(gen[1791]),

			.SELF(gen[1695]),
			.cell_state(gen[1695])
		); 

/******************* CELL 1696 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1696 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1600]),
			.N(gen[1601]),
			.NE(gen[1602]),

			.O(gen[1695]),
			.E(gen[1697]),

			.SO(gen[1790]),
			.S(gen[1791]),
			.SE(gen[1792]),

			.SELF(gen[1696]),
			.cell_state(gen[1696])
		); 

/******************* CELL 1697 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1697 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1601]),
			.N(gen[1602]),
			.NE(gen[1603]),

			.O(gen[1696]),
			.E(gen[1698]),

			.SO(gen[1791]),
			.S(gen[1792]),
			.SE(gen[1793]),

			.SELF(gen[1697]),
			.cell_state(gen[1697])
		); 

/******************* CELL 1698 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1698 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1602]),
			.N(gen[1603]),
			.NE(gen[1604]),

			.O(gen[1697]),
			.E(gen[1699]),

			.SO(gen[1792]),
			.S(gen[1793]),
			.SE(gen[1794]),

			.SELF(gen[1698]),
			.cell_state(gen[1698])
		); 

/******************* CELL 1699 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1699 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1603]),
			.N(gen[1604]),
			.NE(gen[1605]),

			.O(gen[1698]),
			.E(gen[1700]),

			.SO(gen[1793]),
			.S(gen[1794]),
			.SE(gen[1795]),

			.SELF(gen[1699]),
			.cell_state(gen[1699])
		); 

/******************* CELL 1700 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1700 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1604]),
			.N(gen[1605]),
			.NE(gen[1606]),

			.O(gen[1699]),
			.E(gen[1701]),

			.SO(gen[1794]),
			.S(gen[1795]),
			.SE(gen[1796]),

			.SELF(gen[1700]),
			.cell_state(gen[1700])
		); 

/******************* CELL 1701 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1701 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1605]),
			.N(gen[1606]),
			.NE(gen[1607]),

			.O(gen[1700]),
			.E(gen[1702]),

			.SO(gen[1795]),
			.S(gen[1796]),
			.SE(gen[1797]),

			.SELF(gen[1701]),
			.cell_state(gen[1701])
		); 

/******************* CELL 1702 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1702 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1606]),
			.N(gen[1607]),
			.NE(gen[1608]),

			.O(gen[1701]),
			.E(gen[1703]),

			.SO(gen[1796]),
			.S(gen[1797]),
			.SE(gen[1798]),

			.SELF(gen[1702]),
			.cell_state(gen[1702])
		); 

/******************* CELL 1703 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1703 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1607]),
			.N(gen[1608]),
			.NE(gen[1609]),

			.O(gen[1702]),
			.E(gen[1704]),

			.SO(gen[1797]),
			.S(gen[1798]),
			.SE(gen[1799]),

			.SELF(gen[1703]),
			.cell_state(gen[1703])
		); 

/******************* CELL 1704 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1704 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1608]),
			.N(gen[1609]),
			.NE(gen[1610]),

			.O(gen[1703]),
			.E(gen[1705]),

			.SO(gen[1798]),
			.S(gen[1799]),
			.SE(gen[1800]),

			.SELF(gen[1704]),
			.cell_state(gen[1704])
		); 

/******************* CELL 1705 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1705 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1609]),
			.N(gen[1610]),
			.NE(gen[1611]),

			.O(gen[1704]),
			.E(gen[1706]),

			.SO(gen[1799]),
			.S(gen[1800]),
			.SE(gen[1801]),

			.SELF(gen[1705]),
			.cell_state(gen[1705])
		); 

/******************* CELL 1706 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1706 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1610]),
			.N(gen[1611]),
			.NE(gen[1612]),

			.O(gen[1705]),
			.E(gen[1707]),

			.SO(gen[1800]),
			.S(gen[1801]),
			.SE(gen[1802]),

			.SELF(gen[1706]),
			.cell_state(gen[1706])
		); 

/******************* CELL 1707 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1707 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1611]),
			.N(gen[1612]),
			.NE(gen[1613]),

			.O(gen[1706]),
			.E(gen[1708]),

			.SO(gen[1801]),
			.S(gen[1802]),
			.SE(gen[1803]),

			.SELF(gen[1707]),
			.cell_state(gen[1707])
		); 

/******************* CELL 1708 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1708 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1612]),
			.N(gen[1613]),
			.NE(gen[1614]),

			.O(gen[1707]),
			.E(gen[1709]),

			.SO(gen[1802]),
			.S(gen[1803]),
			.SE(gen[1804]),

			.SELF(gen[1708]),
			.cell_state(gen[1708])
		); 

/******************* CELL 1709 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1709 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1613]),
			.N(gen[1614]),
			.NE(gen[1613]),

			.O(gen[1708]),
			.E(gen[1708]),

			.SO(gen[1803]),
			.S(gen[1804]),
			.SE(gen[1803]),

			.SELF(gen[1709]),
			.cell_state(gen[1709])
		); 

/******************* CELL 1710 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1710 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1616]),
			.N(gen[1615]),
			.NE(gen[1616]),

			.O(gen[1711]),
			.E(gen[1711]),

			.SO(gen[1806]),
			.S(gen[1805]),
			.SE(gen[1806]),

			.SELF(gen[1710]),
			.cell_state(gen[1710])
		); 

/******************* CELL 1711 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1711 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1615]),
			.N(gen[1616]),
			.NE(gen[1617]),

			.O(gen[1710]),
			.E(gen[1712]),

			.SO(gen[1805]),
			.S(gen[1806]),
			.SE(gen[1807]),

			.SELF(gen[1711]),
			.cell_state(gen[1711])
		); 

/******************* CELL 1712 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1712 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1616]),
			.N(gen[1617]),
			.NE(gen[1618]),

			.O(gen[1711]),
			.E(gen[1713]),

			.SO(gen[1806]),
			.S(gen[1807]),
			.SE(gen[1808]),

			.SELF(gen[1712]),
			.cell_state(gen[1712])
		); 

/******************* CELL 1713 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1713 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1617]),
			.N(gen[1618]),
			.NE(gen[1619]),

			.O(gen[1712]),
			.E(gen[1714]),

			.SO(gen[1807]),
			.S(gen[1808]),
			.SE(gen[1809]),

			.SELF(gen[1713]),
			.cell_state(gen[1713])
		); 

/******************* CELL 1714 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1714 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1618]),
			.N(gen[1619]),
			.NE(gen[1620]),

			.O(gen[1713]),
			.E(gen[1715]),

			.SO(gen[1808]),
			.S(gen[1809]),
			.SE(gen[1810]),

			.SELF(gen[1714]),
			.cell_state(gen[1714])
		); 

/******************* CELL 1715 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1715 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1619]),
			.N(gen[1620]),
			.NE(gen[1621]),

			.O(gen[1714]),
			.E(gen[1716]),

			.SO(gen[1809]),
			.S(gen[1810]),
			.SE(gen[1811]),

			.SELF(gen[1715]),
			.cell_state(gen[1715])
		); 

/******************* CELL 1716 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1716 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1620]),
			.N(gen[1621]),
			.NE(gen[1622]),

			.O(gen[1715]),
			.E(gen[1717]),

			.SO(gen[1810]),
			.S(gen[1811]),
			.SE(gen[1812]),

			.SELF(gen[1716]),
			.cell_state(gen[1716])
		); 

/******************* CELL 1717 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1717 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1621]),
			.N(gen[1622]),
			.NE(gen[1623]),

			.O(gen[1716]),
			.E(gen[1718]),

			.SO(gen[1811]),
			.S(gen[1812]),
			.SE(gen[1813]),

			.SELF(gen[1717]),
			.cell_state(gen[1717])
		); 

/******************* CELL 1718 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1718 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1622]),
			.N(gen[1623]),
			.NE(gen[1624]),

			.O(gen[1717]),
			.E(gen[1719]),

			.SO(gen[1812]),
			.S(gen[1813]),
			.SE(gen[1814]),

			.SELF(gen[1718]),
			.cell_state(gen[1718])
		); 

/******************* CELL 1719 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1719 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1623]),
			.N(gen[1624]),
			.NE(gen[1625]),

			.O(gen[1718]),
			.E(gen[1720]),

			.SO(gen[1813]),
			.S(gen[1814]),
			.SE(gen[1815]),

			.SELF(gen[1719]),
			.cell_state(gen[1719])
		); 

/******************* CELL 1720 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1720 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1624]),
			.N(gen[1625]),
			.NE(gen[1626]),

			.O(gen[1719]),
			.E(gen[1721]),

			.SO(gen[1814]),
			.S(gen[1815]),
			.SE(gen[1816]),

			.SELF(gen[1720]),
			.cell_state(gen[1720])
		); 

/******************* CELL 1721 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1721 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1625]),
			.N(gen[1626]),
			.NE(gen[1627]),

			.O(gen[1720]),
			.E(gen[1722]),

			.SO(gen[1815]),
			.S(gen[1816]),
			.SE(gen[1817]),

			.SELF(gen[1721]),
			.cell_state(gen[1721])
		); 

/******************* CELL 1722 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1722 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1626]),
			.N(gen[1627]),
			.NE(gen[1628]),

			.O(gen[1721]),
			.E(gen[1723]),

			.SO(gen[1816]),
			.S(gen[1817]),
			.SE(gen[1818]),

			.SELF(gen[1722]),
			.cell_state(gen[1722])
		); 

/******************* CELL 1723 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1723 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1627]),
			.N(gen[1628]),
			.NE(gen[1629]),

			.O(gen[1722]),
			.E(gen[1724]),

			.SO(gen[1817]),
			.S(gen[1818]),
			.SE(gen[1819]),

			.SELF(gen[1723]),
			.cell_state(gen[1723])
		); 

/******************* CELL 1724 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1724 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1628]),
			.N(gen[1629]),
			.NE(gen[1630]),

			.O(gen[1723]),
			.E(gen[1725]),

			.SO(gen[1818]),
			.S(gen[1819]),
			.SE(gen[1820]),

			.SELF(gen[1724]),
			.cell_state(gen[1724])
		); 

/******************* CELL 1725 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1725 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1629]),
			.N(gen[1630]),
			.NE(gen[1631]),

			.O(gen[1724]),
			.E(gen[1726]),

			.SO(gen[1819]),
			.S(gen[1820]),
			.SE(gen[1821]),

			.SELF(gen[1725]),
			.cell_state(gen[1725])
		); 

/******************* CELL 1726 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1726 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1630]),
			.N(gen[1631]),
			.NE(gen[1632]),

			.O(gen[1725]),
			.E(gen[1727]),

			.SO(gen[1820]),
			.S(gen[1821]),
			.SE(gen[1822]),

			.SELF(gen[1726]),
			.cell_state(gen[1726])
		); 

/******************* CELL 1727 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1727 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1631]),
			.N(gen[1632]),
			.NE(gen[1633]),

			.O(gen[1726]),
			.E(gen[1728]),

			.SO(gen[1821]),
			.S(gen[1822]),
			.SE(gen[1823]),

			.SELF(gen[1727]),
			.cell_state(gen[1727])
		); 

/******************* CELL 1728 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1728 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1632]),
			.N(gen[1633]),
			.NE(gen[1634]),

			.O(gen[1727]),
			.E(gen[1729]),

			.SO(gen[1822]),
			.S(gen[1823]),
			.SE(gen[1824]),

			.SELF(gen[1728]),
			.cell_state(gen[1728])
		); 

/******************* CELL 1729 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1729 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1633]),
			.N(gen[1634]),
			.NE(gen[1635]),

			.O(gen[1728]),
			.E(gen[1730]),

			.SO(gen[1823]),
			.S(gen[1824]),
			.SE(gen[1825]),

			.SELF(gen[1729]),
			.cell_state(gen[1729])
		); 

/******************* CELL 1730 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1730 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1634]),
			.N(gen[1635]),
			.NE(gen[1636]),

			.O(gen[1729]),
			.E(gen[1731]),

			.SO(gen[1824]),
			.S(gen[1825]),
			.SE(gen[1826]),

			.SELF(gen[1730]),
			.cell_state(gen[1730])
		); 

/******************* CELL 1731 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1731 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1635]),
			.N(gen[1636]),
			.NE(gen[1637]),

			.O(gen[1730]),
			.E(gen[1732]),

			.SO(gen[1825]),
			.S(gen[1826]),
			.SE(gen[1827]),

			.SELF(gen[1731]),
			.cell_state(gen[1731])
		); 

/******************* CELL 1732 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1732 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1636]),
			.N(gen[1637]),
			.NE(gen[1638]),

			.O(gen[1731]),
			.E(gen[1733]),

			.SO(gen[1826]),
			.S(gen[1827]),
			.SE(gen[1828]),

			.SELF(gen[1732]),
			.cell_state(gen[1732])
		); 

/******************* CELL 1733 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1733 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1637]),
			.N(gen[1638]),
			.NE(gen[1639]),

			.O(gen[1732]),
			.E(gen[1734]),

			.SO(gen[1827]),
			.S(gen[1828]),
			.SE(gen[1829]),

			.SELF(gen[1733]),
			.cell_state(gen[1733])
		); 

/******************* CELL 1734 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1734 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1638]),
			.N(gen[1639]),
			.NE(gen[1640]),

			.O(gen[1733]),
			.E(gen[1735]),

			.SO(gen[1828]),
			.S(gen[1829]),
			.SE(gen[1830]),

			.SELF(gen[1734]),
			.cell_state(gen[1734])
		); 

/******************* CELL 1735 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1735 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1639]),
			.N(gen[1640]),
			.NE(gen[1641]),

			.O(gen[1734]),
			.E(gen[1736]),

			.SO(gen[1829]),
			.S(gen[1830]),
			.SE(gen[1831]),

			.SELF(gen[1735]),
			.cell_state(gen[1735])
		); 

/******************* CELL 1736 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1736 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1640]),
			.N(gen[1641]),
			.NE(gen[1642]),

			.O(gen[1735]),
			.E(gen[1737]),

			.SO(gen[1830]),
			.S(gen[1831]),
			.SE(gen[1832]),

			.SELF(gen[1736]),
			.cell_state(gen[1736])
		); 

/******************* CELL 1737 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1737 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1641]),
			.N(gen[1642]),
			.NE(gen[1643]),

			.O(gen[1736]),
			.E(gen[1738]),

			.SO(gen[1831]),
			.S(gen[1832]),
			.SE(gen[1833]),

			.SELF(gen[1737]),
			.cell_state(gen[1737])
		); 

/******************* CELL 1738 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1738 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1642]),
			.N(gen[1643]),
			.NE(gen[1644]),

			.O(gen[1737]),
			.E(gen[1739]),

			.SO(gen[1832]),
			.S(gen[1833]),
			.SE(gen[1834]),

			.SELF(gen[1738]),
			.cell_state(gen[1738])
		); 

/******************* CELL 1739 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1739 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1643]),
			.N(gen[1644]),
			.NE(gen[1645]),

			.O(gen[1738]),
			.E(gen[1740]),

			.SO(gen[1833]),
			.S(gen[1834]),
			.SE(gen[1835]),

			.SELF(gen[1739]),
			.cell_state(gen[1739])
		); 

/******************* CELL 1740 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1740 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1644]),
			.N(gen[1645]),
			.NE(gen[1646]),

			.O(gen[1739]),
			.E(gen[1741]),

			.SO(gen[1834]),
			.S(gen[1835]),
			.SE(gen[1836]),

			.SELF(gen[1740]),
			.cell_state(gen[1740])
		); 

/******************* CELL 1741 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1741 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1645]),
			.N(gen[1646]),
			.NE(gen[1647]),

			.O(gen[1740]),
			.E(gen[1742]),

			.SO(gen[1835]),
			.S(gen[1836]),
			.SE(gen[1837]),

			.SELF(gen[1741]),
			.cell_state(gen[1741])
		); 

/******************* CELL 1742 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1742 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1646]),
			.N(gen[1647]),
			.NE(gen[1648]),

			.O(gen[1741]),
			.E(gen[1743]),

			.SO(gen[1836]),
			.S(gen[1837]),
			.SE(gen[1838]),

			.SELF(gen[1742]),
			.cell_state(gen[1742])
		); 

/******************* CELL 1743 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1743 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1647]),
			.N(gen[1648]),
			.NE(gen[1649]),

			.O(gen[1742]),
			.E(gen[1744]),

			.SO(gen[1837]),
			.S(gen[1838]),
			.SE(gen[1839]),

			.SELF(gen[1743]),
			.cell_state(gen[1743])
		); 

/******************* CELL 1744 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1744 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1648]),
			.N(gen[1649]),
			.NE(gen[1650]),

			.O(gen[1743]),
			.E(gen[1745]),

			.SO(gen[1838]),
			.S(gen[1839]),
			.SE(gen[1840]),

			.SELF(gen[1744]),
			.cell_state(gen[1744])
		); 

/******************* CELL 1745 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1745 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1649]),
			.N(gen[1650]),
			.NE(gen[1651]),

			.O(gen[1744]),
			.E(gen[1746]),

			.SO(gen[1839]),
			.S(gen[1840]),
			.SE(gen[1841]),

			.SELF(gen[1745]),
			.cell_state(gen[1745])
		); 

/******************* CELL 1746 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1746 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1650]),
			.N(gen[1651]),
			.NE(gen[1652]),

			.O(gen[1745]),
			.E(gen[1747]),

			.SO(gen[1840]),
			.S(gen[1841]),
			.SE(gen[1842]),

			.SELF(gen[1746]),
			.cell_state(gen[1746])
		); 

/******************* CELL 1747 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1747 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1651]),
			.N(gen[1652]),
			.NE(gen[1653]),

			.O(gen[1746]),
			.E(gen[1748]),

			.SO(gen[1841]),
			.S(gen[1842]),
			.SE(gen[1843]),

			.SELF(gen[1747]),
			.cell_state(gen[1747])
		); 

/******************* CELL 1748 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1748 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1652]),
			.N(gen[1653]),
			.NE(gen[1654]),

			.O(gen[1747]),
			.E(gen[1749]),

			.SO(gen[1842]),
			.S(gen[1843]),
			.SE(gen[1844]),

			.SELF(gen[1748]),
			.cell_state(gen[1748])
		); 

/******************* CELL 1749 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1749 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1653]),
			.N(gen[1654]),
			.NE(gen[1655]),

			.O(gen[1748]),
			.E(gen[1750]),

			.SO(gen[1843]),
			.S(gen[1844]),
			.SE(gen[1845]),

			.SELF(gen[1749]),
			.cell_state(gen[1749])
		); 

/******************* CELL 1750 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1750 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1654]),
			.N(gen[1655]),
			.NE(gen[1656]),

			.O(gen[1749]),
			.E(gen[1751]),

			.SO(gen[1844]),
			.S(gen[1845]),
			.SE(gen[1846]),

			.SELF(gen[1750]),
			.cell_state(gen[1750])
		); 

/******************* CELL 1751 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1751 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1655]),
			.N(gen[1656]),
			.NE(gen[1657]),

			.O(gen[1750]),
			.E(gen[1752]),

			.SO(gen[1845]),
			.S(gen[1846]),
			.SE(gen[1847]),

			.SELF(gen[1751]),
			.cell_state(gen[1751])
		); 

/******************* CELL 1752 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1752 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1656]),
			.N(gen[1657]),
			.NE(gen[1658]),

			.O(gen[1751]),
			.E(gen[1753]),

			.SO(gen[1846]),
			.S(gen[1847]),
			.SE(gen[1848]),

			.SELF(gen[1752]),
			.cell_state(gen[1752])
		); 

/******************* CELL 1753 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1753 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1657]),
			.N(gen[1658]),
			.NE(gen[1659]),

			.O(gen[1752]),
			.E(gen[1754]),

			.SO(gen[1847]),
			.S(gen[1848]),
			.SE(gen[1849]),

			.SELF(gen[1753]),
			.cell_state(gen[1753])
		); 

/******************* CELL 1754 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1754 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1658]),
			.N(gen[1659]),
			.NE(gen[1660]),

			.O(gen[1753]),
			.E(gen[1755]),

			.SO(gen[1848]),
			.S(gen[1849]),
			.SE(gen[1850]),

			.SELF(gen[1754]),
			.cell_state(gen[1754])
		); 

/******************* CELL 1755 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1755 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1659]),
			.N(gen[1660]),
			.NE(gen[1661]),

			.O(gen[1754]),
			.E(gen[1756]),

			.SO(gen[1849]),
			.S(gen[1850]),
			.SE(gen[1851]),

			.SELF(gen[1755]),
			.cell_state(gen[1755])
		); 

/******************* CELL 1756 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1756 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1660]),
			.N(gen[1661]),
			.NE(gen[1662]),

			.O(gen[1755]),
			.E(gen[1757]),

			.SO(gen[1850]),
			.S(gen[1851]),
			.SE(gen[1852]),

			.SELF(gen[1756]),
			.cell_state(gen[1756])
		); 

/******************* CELL 1757 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1757 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1661]),
			.N(gen[1662]),
			.NE(gen[1663]),

			.O(gen[1756]),
			.E(gen[1758]),

			.SO(gen[1851]),
			.S(gen[1852]),
			.SE(gen[1853]),

			.SELF(gen[1757]),
			.cell_state(gen[1757])
		); 

/******************* CELL 1758 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1758 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1662]),
			.N(gen[1663]),
			.NE(gen[1664]),

			.O(gen[1757]),
			.E(gen[1759]),

			.SO(gen[1852]),
			.S(gen[1853]),
			.SE(gen[1854]),

			.SELF(gen[1758]),
			.cell_state(gen[1758])
		); 

/******************* CELL 1759 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1759 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1663]),
			.N(gen[1664]),
			.NE(gen[1665]),

			.O(gen[1758]),
			.E(gen[1760]),

			.SO(gen[1853]),
			.S(gen[1854]),
			.SE(gen[1855]),

			.SELF(gen[1759]),
			.cell_state(gen[1759])
		); 

/******************* CELL 1760 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1760 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1664]),
			.N(gen[1665]),
			.NE(gen[1666]),

			.O(gen[1759]),
			.E(gen[1761]),

			.SO(gen[1854]),
			.S(gen[1855]),
			.SE(gen[1856]),

			.SELF(gen[1760]),
			.cell_state(gen[1760])
		); 

/******************* CELL 1761 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1761 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1665]),
			.N(gen[1666]),
			.NE(gen[1667]),

			.O(gen[1760]),
			.E(gen[1762]),

			.SO(gen[1855]),
			.S(gen[1856]),
			.SE(gen[1857]),

			.SELF(gen[1761]),
			.cell_state(gen[1761])
		); 

/******************* CELL 1762 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1762 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1666]),
			.N(gen[1667]),
			.NE(gen[1668]),

			.O(gen[1761]),
			.E(gen[1763]),

			.SO(gen[1856]),
			.S(gen[1857]),
			.SE(gen[1858]),

			.SELF(gen[1762]),
			.cell_state(gen[1762])
		); 

/******************* CELL 1763 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1763 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1667]),
			.N(gen[1668]),
			.NE(gen[1669]),

			.O(gen[1762]),
			.E(gen[1764]),

			.SO(gen[1857]),
			.S(gen[1858]),
			.SE(gen[1859]),

			.SELF(gen[1763]),
			.cell_state(gen[1763])
		); 

/******************* CELL 1764 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1764 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1668]),
			.N(gen[1669]),
			.NE(gen[1670]),

			.O(gen[1763]),
			.E(gen[1765]),

			.SO(gen[1858]),
			.S(gen[1859]),
			.SE(gen[1860]),

			.SELF(gen[1764]),
			.cell_state(gen[1764])
		); 

/******************* CELL 1765 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1765 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1669]),
			.N(gen[1670]),
			.NE(gen[1671]),

			.O(gen[1764]),
			.E(gen[1766]),

			.SO(gen[1859]),
			.S(gen[1860]),
			.SE(gen[1861]),

			.SELF(gen[1765]),
			.cell_state(gen[1765])
		); 

/******************* CELL 1766 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1766 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1670]),
			.N(gen[1671]),
			.NE(gen[1672]),

			.O(gen[1765]),
			.E(gen[1767]),

			.SO(gen[1860]),
			.S(gen[1861]),
			.SE(gen[1862]),

			.SELF(gen[1766]),
			.cell_state(gen[1766])
		); 

/******************* CELL 1767 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1767 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1671]),
			.N(gen[1672]),
			.NE(gen[1673]),

			.O(gen[1766]),
			.E(gen[1768]),

			.SO(gen[1861]),
			.S(gen[1862]),
			.SE(gen[1863]),

			.SELF(gen[1767]),
			.cell_state(gen[1767])
		); 

/******************* CELL 1768 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1768 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1672]),
			.N(gen[1673]),
			.NE(gen[1674]),

			.O(gen[1767]),
			.E(gen[1769]),

			.SO(gen[1862]),
			.S(gen[1863]),
			.SE(gen[1864]),

			.SELF(gen[1768]),
			.cell_state(gen[1768])
		); 

/******************* CELL 1769 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1769 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1673]),
			.N(gen[1674]),
			.NE(gen[1675]),

			.O(gen[1768]),
			.E(gen[1770]),

			.SO(gen[1863]),
			.S(gen[1864]),
			.SE(gen[1865]),

			.SELF(gen[1769]),
			.cell_state(gen[1769])
		); 

/******************* CELL 1770 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1770 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1674]),
			.N(gen[1675]),
			.NE(gen[1676]),

			.O(gen[1769]),
			.E(gen[1771]),

			.SO(gen[1864]),
			.S(gen[1865]),
			.SE(gen[1866]),

			.SELF(gen[1770]),
			.cell_state(gen[1770])
		); 

/******************* CELL 1771 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1771 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1675]),
			.N(gen[1676]),
			.NE(gen[1677]),

			.O(gen[1770]),
			.E(gen[1772]),

			.SO(gen[1865]),
			.S(gen[1866]),
			.SE(gen[1867]),

			.SELF(gen[1771]),
			.cell_state(gen[1771])
		); 

/******************* CELL 1772 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1772 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1676]),
			.N(gen[1677]),
			.NE(gen[1678]),

			.O(gen[1771]),
			.E(gen[1773]),

			.SO(gen[1866]),
			.S(gen[1867]),
			.SE(gen[1868]),

			.SELF(gen[1772]),
			.cell_state(gen[1772])
		); 

/******************* CELL 1773 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1773 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1677]),
			.N(gen[1678]),
			.NE(gen[1679]),

			.O(gen[1772]),
			.E(gen[1774]),

			.SO(gen[1867]),
			.S(gen[1868]),
			.SE(gen[1869]),

			.SELF(gen[1773]),
			.cell_state(gen[1773])
		); 

/******************* CELL 1774 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1774 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1678]),
			.N(gen[1679]),
			.NE(gen[1680]),

			.O(gen[1773]),
			.E(gen[1775]),

			.SO(gen[1868]),
			.S(gen[1869]),
			.SE(gen[1870]),

			.SELF(gen[1774]),
			.cell_state(gen[1774])
		); 

/******************* CELL 1775 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1775 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1679]),
			.N(gen[1680]),
			.NE(gen[1681]),

			.O(gen[1774]),
			.E(gen[1776]),

			.SO(gen[1869]),
			.S(gen[1870]),
			.SE(gen[1871]),

			.SELF(gen[1775]),
			.cell_state(gen[1775])
		); 

/******************* CELL 1776 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1776 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1680]),
			.N(gen[1681]),
			.NE(gen[1682]),

			.O(gen[1775]),
			.E(gen[1777]),

			.SO(gen[1870]),
			.S(gen[1871]),
			.SE(gen[1872]),

			.SELF(gen[1776]),
			.cell_state(gen[1776])
		); 

/******************* CELL 1777 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1777 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1681]),
			.N(gen[1682]),
			.NE(gen[1683]),

			.O(gen[1776]),
			.E(gen[1778]),

			.SO(gen[1871]),
			.S(gen[1872]),
			.SE(gen[1873]),

			.SELF(gen[1777]),
			.cell_state(gen[1777])
		); 

/******************* CELL 1778 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1778 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1682]),
			.N(gen[1683]),
			.NE(gen[1684]),

			.O(gen[1777]),
			.E(gen[1779]),

			.SO(gen[1872]),
			.S(gen[1873]),
			.SE(gen[1874]),

			.SELF(gen[1778]),
			.cell_state(gen[1778])
		); 

/******************* CELL 1779 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1779 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1683]),
			.N(gen[1684]),
			.NE(gen[1685]),

			.O(gen[1778]),
			.E(gen[1780]),

			.SO(gen[1873]),
			.S(gen[1874]),
			.SE(gen[1875]),

			.SELF(gen[1779]),
			.cell_state(gen[1779])
		); 

/******************* CELL 1780 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1780 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1684]),
			.N(gen[1685]),
			.NE(gen[1686]),

			.O(gen[1779]),
			.E(gen[1781]),

			.SO(gen[1874]),
			.S(gen[1875]),
			.SE(gen[1876]),

			.SELF(gen[1780]),
			.cell_state(gen[1780])
		); 

/******************* CELL 1781 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1781 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1685]),
			.N(gen[1686]),
			.NE(gen[1687]),

			.O(gen[1780]),
			.E(gen[1782]),

			.SO(gen[1875]),
			.S(gen[1876]),
			.SE(gen[1877]),

			.SELF(gen[1781]),
			.cell_state(gen[1781])
		); 

/******************* CELL 1782 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1782 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1686]),
			.N(gen[1687]),
			.NE(gen[1688]),

			.O(gen[1781]),
			.E(gen[1783]),

			.SO(gen[1876]),
			.S(gen[1877]),
			.SE(gen[1878]),

			.SELF(gen[1782]),
			.cell_state(gen[1782])
		); 

/******************* CELL 1783 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1783 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1687]),
			.N(gen[1688]),
			.NE(gen[1689]),

			.O(gen[1782]),
			.E(gen[1784]),

			.SO(gen[1877]),
			.S(gen[1878]),
			.SE(gen[1879]),

			.SELF(gen[1783]),
			.cell_state(gen[1783])
		); 

/******************* CELL 1784 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1784 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1688]),
			.N(gen[1689]),
			.NE(gen[1690]),

			.O(gen[1783]),
			.E(gen[1785]),

			.SO(gen[1878]),
			.S(gen[1879]),
			.SE(gen[1880]),

			.SELF(gen[1784]),
			.cell_state(gen[1784])
		); 

/******************* CELL 1785 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1785 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1689]),
			.N(gen[1690]),
			.NE(gen[1691]),

			.O(gen[1784]),
			.E(gen[1786]),

			.SO(gen[1879]),
			.S(gen[1880]),
			.SE(gen[1881]),

			.SELF(gen[1785]),
			.cell_state(gen[1785])
		); 

/******************* CELL 1786 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1786 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1690]),
			.N(gen[1691]),
			.NE(gen[1692]),

			.O(gen[1785]),
			.E(gen[1787]),

			.SO(gen[1880]),
			.S(gen[1881]),
			.SE(gen[1882]),

			.SELF(gen[1786]),
			.cell_state(gen[1786])
		); 

/******************* CELL 1787 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1787 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1691]),
			.N(gen[1692]),
			.NE(gen[1693]),

			.O(gen[1786]),
			.E(gen[1788]),

			.SO(gen[1881]),
			.S(gen[1882]),
			.SE(gen[1883]),

			.SELF(gen[1787]),
			.cell_state(gen[1787])
		); 

/******************* CELL 1788 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1788 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1692]),
			.N(gen[1693]),
			.NE(gen[1694]),

			.O(gen[1787]),
			.E(gen[1789]),

			.SO(gen[1882]),
			.S(gen[1883]),
			.SE(gen[1884]),

			.SELF(gen[1788]),
			.cell_state(gen[1788])
		); 

/******************* CELL 1789 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1789 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1693]),
			.N(gen[1694]),
			.NE(gen[1695]),

			.O(gen[1788]),
			.E(gen[1790]),

			.SO(gen[1883]),
			.S(gen[1884]),
			.SE(gen[1885]),

			.SELF(gen[1789]),
			.cell_state(gen[1789])
		); 

/******************* CELL 1790 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1790 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1694]),
			.N(gen[1695]),
			.NE(gen[1696]),

			.O(gen[1789]),
			.E(gen[1791]),

			.SO(gen[1884]),
			.S(gen[1885]),
			.SE(gen[1886]),

			.SELF(gen[1790]),
			.cell_state(gen[1790])
		); 

/******************* CELL 1791 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1791 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1695]),
			.N(gen[1696]),
			.NE(gen[1697]),

			.O(gen[1790]),
			.E(gen[1792]),

			.SO(gen[1885]),
			.S(gen[1886]),
			.SE(gen[1887]),

			.SELF(gen[1791]),
			.cell_state(gen[1791])
		); 

/******************* CELL 1792 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1792 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1696]),
			.N(gen[1697]),
			.NE(gen[1698]),

			.O(gen[1791]),
			.E(gen[1793]),

			.SO(gen[1886]),
			.S(gen[1887]),
			.SE(gen[1888]),

			.SELF(gen[1792]),
			.cell_state(gen[1792])
		); 

/******************* CELL 1793 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1793 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1697]),
			.N(gen[1698]),
			.NE(gen[1699]),

			.O(gen[1792]),
			.E(gen[1794]),

			.SO(gen[1887]),
			.S(gen[1888]),
			.SE(gen[1889]),

			.SELF(gen[1793]),
			.cell_state(gen[1793])
		); 

/******************* CELL 1794 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1794 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1698]),
			.N(gen[1699]),
			.NE(gen[1700]),

			.O(gen[1793]),
			.E(gen[1795]),

			.SO(gen[1888]),
			.S(gen[1889]),
			.SE(gen[1890]),

			.SELF(gen[1794]),
			.cell_state(gen[1794])
		); 

/******************* CELL 1795 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1795 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1699]),
			.N(gen[1700]),
			.NE(gen[1701]),

			.O(gen[1794]),
			.E(gen[1796]),

			.SO(gen[1889]),
			.S(gen[1890]),
			.SE(gen[1891]),

			.SELF(gen[1795]),
			.cell_state(gen[1795])
		); 

/******************* CELL 1796 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1796 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1700]),
			.N(gen[1701]),
			.NE(gen[1702]),

			.O(gen[1795]),
			.E(gen[1797]),

			.SO(gen[1890]),
			.S(gen[1891]),
			.SE(gen[1892]),

			.SELF(gen[1796]),
			.cell_state(gen[1796])
		); 

/******************* CELL 1797 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1797 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1701]),
			.N(gen[1702]),
			.NE(gen[1703]),

			.O(gen[1796]),
			.E(gen[1798]),

			.SO(gen[1891]),
			.S(gen[1892]),
			.SE(gen[1893]),

			.SELF(gen[1797]),
			.cell_state(gen[1797])
		); 

/******************* CELL 1798 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1798 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1702]),
			.N(gen[1703]),
			.NE(gen[1704]),

			.O(gen[1797]),
			.E(gen[1799]),

			.SO(gen[1892]),
			.S(gen[1893]),
			.SE(gen[1894]),

			.SELF(gen[1798]),
			.cell_state(gen[1798])
		); 

/******************* CELL 1799 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1799 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1703]),
			.N(gen[1704]),
			.NE(gen[1705]),

			.O(gen[1798]),
			.E(gen[1800]),

			.SO(gen[1893]),
			.S(gen[1894]),
			.SE(gen[1895]),

			.SELF(gen[1799]),
			.cell_state(gen[1799])
		); 

/******************* CELL 1800 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1800 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1704]),
			.N(gen[1705]),
			.NE(gen[1706]),

			.O(gen[1799]),
			.E(gen[1801]),

			.SO(gen[1894]),
			.S(gen[1895]),
			.SE(gen[1896]),

			.SELF(gen[1800]),
			.cell_state(gen[1800])
		); 

/******************* CELL 1801 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1801 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1705]),
			.N(gen[1706]),
			.NE(gen[1707]),

			.O(gen[1800]),
			.E(gen[1802]),

			.SO(gen[1895]),
			.S(gen[1896]),
			.SE(gen[1897]),

			.SELF(gen[1801]),
			.cell_state(gen[1801])
		); 

/******************* CELL 1802 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1802 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1706]),
			.N(gen[1707]),
			.NE(gen[1708]),

			.O(gen[1801]),
			.E(gen[1803]),

			.SO(gen[1896]),
			.S(gen[1897]),
			.SE(gen[1898]),

			.SELF(gen[1802]),
			.cell_state(gen[1802])
		); 

/******************* CELL 1803 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1803 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1707]),
			.N(gen[1708]),
			.NE(gen[1709]),

			.O(gen[1802]),
			.E(gen[1804]),

			.SO(gen[1897]),
			.S(gen[1898]),
			.SE(gen[1899]),

			.SELF(gen[1803]),
			.cell_state(gen[1803])
		); 

/******************* CELL 1804 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1804 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1708]),
			.N(gen[1709]),
			.NE(gen[1708]),

			.O(gen[1803]),
			.E(gen[1803]),

			.SO(gen[1898]),
			.S(gen[1899]),
			.SE(gen[1898]),

			.SELF(gen[1804]),
			.cell_state(gen[1804])
		); 

/******************* CELL 1805 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1805 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1711]),
			.N(gen[1710]),
			.NE(gen[1711]),

			.O(gen[1806]),
			.E(gen[1806]),

			.SO(gen[1901]),
			.S(gen[1900]),
			.SE(gen[1901]),

			.SELF(gen[1805]),
			.cell_state(gen[1805])
		); 

/******************* CELL 1806 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1806 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1710]),
			.N(gen[1711]),
			.NE(gen[1712]),

			.O(gen[1805]),
			.E(gen[1807]),

			.SO(gen[1900]),
			.S(gen[1901]),
			.SE(gen[1902]),

			.SELF(gen[1806]),
			.cell_state(gen[1806])
		); 

/******************* CELL 1807 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1807 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1711]),
			.N(gen[1712]),
			.NE(gen[1713]),

			.O(gen[1806]),
			.E(gen[1808]),

			.SO(gen[1901]),
			.S(gen[1902]),
			.SE(gen[1903]),

			.SELF(gen[1807]),
			.cell_state(gen[1807])
		); 

/******************* CELL 1808 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1808 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1712]),
			.N(gen[1713]),
			.NE(gen[1714]),

			.O(gen[1807]),
			.E(gen[1809]),

			.SO(gen[1902]),
			.S(gen[1903]),
			.SE(gen[1904]),

			.SELF(gen[1808]),
			.cell_state(gen[1808])
		); 

/******************* CELL 1809 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1809 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1713]),
			.N(gen[1714]),
			.NE(gen[1715]),

			.O(gen[1808]),
			.E(gen[1810]),

			.SO(gen[1903]),
			.S(gen[1904]),
			.SE(gen[1905]),

			.SELF(gen[1809]),
			.cell_state(gen[1809])
		); 

/******************* CELL 1810 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1810 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1714]),
			.N(gen[1715]),
			.NE(gen[1716]),

			.O(gen[1809]),
			.E(gen[1811]),

			.SO(gen[1904]),
			.S(gen[1905]),
			.SE(gen[1906]),

			.SELF(gen[1810]),
			.cell_state(gen[1810])
		); 

/******************* CELL 1811 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1811 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1715]),
			.N(gen[1716]),
			.NE(gen[1717]),

			.O(gen[1810]),
			.E(gen[1812]),

			.SO(gen[1905]),
			.S(gen[1906]),
			.SE(gen[1907]),

			.SELF(gen[1811]),
			.cell_state(gen[1811])
		); 

/******************* CELL 1812 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1812 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1716]),
			.N(gen[1717]),
			.NE(gen[1718]),

			.O(gen[1811]),
			.E(gen[1813]),

			.SO(gen[1906]),
			.S(gen[1907]),
			.SE(gen[1908]),

			.SELF(gen[1812]),
			.cell_state(gen[1812])
		); 

/******************* CELL 1813 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1813 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1717]),
			.N(gen[1718]),
			.NE(gen[1719]),

			.O(gen[1812]),
			.E(gen[1814]),

			.SO(gen[1907]),
			.S(gen[1908]),
			.SE(gen[1909]),

			.SELF(gen[1813]),
			.cell_state(gen[1813])
		); 

/******************* CELL 1814 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1814 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1718]),
			.N(gen[1719]),
			.NE(gen[1720]),

			.O(gen[1813]),
			.E(gen[1815]),

			.SO(gen[1908]),
			.S(gen[1909]),
			.SE(gen[1910]),

			.SELF(gen[1814]),
			.cell_state(gen[1814])
		); 

/******************* CELL 1815 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1815 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1719]),
			.N(gen[1720]),
			.NE(gen[1721]),

			.O(gen[1814]),
			.E(gen[1816]),

			.SO(gen[1909]),
			.S(gen[1910]),
			.SE(gen[1911]),

			.SELF(gen[1815]),
			.cell_state(gen[1815])
		); 

/******************* CELL 1816 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1816 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1720]),
			.N(gen[1721]),
			.NE(gen[1722]),

			.O(gen[1815]),
			.E(gen[1817]),

			.SO(gen[1910]),
			.S(gen[1911]),
			.SE(gen[1912]),

			.SELF(gen[1816]),
			.cell_state(gen[1816])
		); 

/******************* CELL 1817 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1817 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1721]),
			.N(gen[1722]),
			.NE(gen[1723]),

			.O(gen[1816]),
			.E(gen[1818]),

			.SO(gen[1911]),
			.S(gen[1912]),
			.SE(gen[1913]),

			.SELF(gen[1817]),
			.cell_state(gen[1817])
		); 

/******************* CELL 1818 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1818 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1722]),
			.N(gen[1723]),
			.NE(gen[1724]),

			.O(gen[1817]),
			.E(gen[1819]),

			.SO(gen[1912]),
			.S(gen[1913]),
			.SE(gen[1914]),

			.SELF(gen[1818]),
			.cell_state(gen[1818])
		); 

/******************* CELL 1819 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1819 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1723]),
			.N(gen[1724]),
			.NE(gen[1725]),

			.O(gen[1818]),
			.E(gen[1820]),

			.SO(gen[1913]),
			.S(gen[1914]),
			.SE(gen[1915]),

			.SELF(gen[1819]),
			.cell_state(gen[1819])
		); 

/******************* CELL 1820 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1820 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1724]),
			.N(gen[1725]),
			.NE(gen[1726]),

			.O(gen[1819]),
			.E(gen[1821]),

			.SO(gen[1914]),
			.S(gen[1915]),
			.SE(gen[1916]),

			.SELF(gen[1820]),
			.cell_state(gen[1820])
		); 

/******************* CELL 1821 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1821 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1725]),
			.N(gen[1726]),
			.NE(gen[1727]),

			.O(gen[1820]),
			.E(gen[1822]),

			.SO(gen[1915]),
			.S(gen[1916]),
			.SE(gen[1917]),

			.SELF(gen[1821]),
			.cell_state(gen[1821])
		); 

/******************* CELL 1822 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1822 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1726]),
			.N(gen[1727]),
			.NE(gen[1728]),

			.O(gen[1821]),
			.E(gen[1823]),

			.SO(gen[1916]),
			.S(gen[1917]),
			.SE(gen[1918]),

			.SELF(gen[1822]),
			.cell_state(gen[1822])
		); 

/******************* CELL 1823 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1823 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1727]),
			.N(gen[1728]),
			.NE(gen[1729]),

			.O(gen[1822]),
			.E(gen[1824]),

			.SO(gen[1917]),
			.S(gen[1918]),
			.SE(gen[1919]),

			.SELF(gen[1823]),
			.cell_state(gen[1823])
		); 

/******************* CELL 1824 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1824 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1728]),
			.N(gen[1729]),
			.NE(gen[1730]),

			.O(gen[1823]),
			.E(gen[1825]),

			.SO(gen[1918]),
			.S(gen[1919]),
			.SE(gen[1920]),

			.SELF(gen[1824]),
			.cell_state(gen[1824])
		); 

/******************* CELL 1825 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1825 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1729]),
			.N(gen[1730]),
			.NE(gen[1731]),

			.O(gen[1824]),
			.E(gen[1826]),

			.SO(gen[1919]),
			.S(gen[1920]),
			.SE(gen[1921]),

			.SELF(gen[1825]),
			.cell_state(gen[1825])
		); 

/******************* CELL 1826 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1826 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1730]),
			.N(gen[1731]),
			.NE(gen[1732]),

			.O(gen[1825]),
			.E(gen[1827]),

			.SO(gen[1920]),
			.S(gen[1921]),
			.SE(gen[1922]),

			.SELF(gen[1826]),
			.cell_state(gen[1826])
		); 

/******************* CELL 1827 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1827 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1731]),
			.N(gen[1732]),
			.NE(gen[1733]),

			.O(gen[1826]),
			.E(gen[1828]),

			.SO(gen[1921]),
			.S(gen[1922]),
			.SE(gen[1923]),

			.SELF(gen[1827]),
			.cell_state(gen[1827])
		); 

/******************* CELL 1828 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1828 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1732]),
			.N(gen[1733]),
			.NE(gen[1734]),

			.O(gen[1827]),
			.E(gen[1829]),

			.SO(gen[1922]),
			.S(gen[1923]),
			.SE(gen[1924]),

			.SELF(gen[1828]),
			.cell_state(gen[1828])
		); 

/******************* CELL 1829 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1829 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1733]),
			.N(gen[1734]),
			.NE(gen[1735]),

			.O(gen[1828]),
			.E(gen[1830]),

			.SO(gen[1923]),
			.S(gen[1924]),
			.SE(gen[1925]),

			.SELF(gen[1829]),
			.cell_state(gen[1829])
		); 

/******************* CELL 1830 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1830 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1734]),
			.N(gen[1735]),
			.NE(gen[1736]),

			.O(gen[1829]),
			.E(gen[1831]),

			.SO(gen[1924]),
			.S(gen[1925]),
			.SE(gen[1926]),

			.SELF(gen[1830]),
			.cell_state(gen[1830])
		); 

/******************* CELL 1831 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1831 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1735]),
			.N(gen[1736]),
			.NE(gen[1737]),

			.O(gen[1830]),
			.E(gen[1832]),

			.SO(gen[1925]),
			.S(gen[1926]),
			.SE(gen[1927]),

			.SELF(gen[1831]),
			.cell_state(gen[1831])
		); 

/******************* CELL 1832 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1832 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1736]),
			.N(gen[1737]),
			.NE(gen[1738]),

			.O(gen[1831]),
			.E(gen[1833]),

			.SO(gen[1926]),
			.S(gen[1927]),
			.SE(gen[1928]),

			.SELF(gen[1832]),
			.cell_state(gen[1832])
		); 

/******************* CELL 1833 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1833 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1737]),
			.N(gen[1738]),
			.NE(gen[1739]),

			.O(gen[1832]),
			.E(gen[1834]),

			.SO(gen[1927]),
			.S(gen[1928]),
			.SE(gen[1929]),

			.SELF(gen[1833]),
			.cell_state(gen[1833])
		); 

/******************* CELL 1834 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1834 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1738]),
			.N(gen[1739]),
			.NE(gen[1740]),

			.O(gen[1833]),
			.E(gen[1835]),

			.SO(gen[1928]),
			.S(gen[1929]),
			.SE(gen[1930]),

			.SELF(gen[1834]),
			.cell_state(gen[1834])
		); 

/******************* CELL 1835 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1835 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1739]),
			.N(gen[1740]),
			.NE(gen[1741]),

			.O(gen[1834]),
			.E(gen[1836]),

			.SO(gen[1929]),
			.S(gen[1930]),
			.SE(gen[1931]),

			.SELF(gen[1835]),
			.cell_state(gen[1835])
		); 

/******************* CELL 1836 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1836 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1740]),
			.N(gen[1741]),
			.NE(gen[1742]),

			.O(gen[1835]),
			.E(gen[1837]),

			.SO(gen[1930]),
			.S(gen[1931]),
			.SE(gen[1932]),

			.SELF(gen[1836]),
			.cell_state(gen[1836])
		); 

/******************* CELL 1837 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1837 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1741]),
			.N(gen[1742]),
			.NE(gen[1743]),

			.O(gen[1836]),
			.E(gen[1838]),

			.SO(gen[1931]),
			.S(gen[1932]),
			.SE(gen[1933]),

			.SELF(gen[1837]),
			.cell_state(gen[1837])
		); 

/******************* CELL 1838 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1838 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1742]),
			.N(gen[1743]),
			.NE(gen[1744]),

			.O(gen[1837]),
			.E(gen[1839]),

			.SO(gen[1932]),
			.S(gen[1933]),
			.SE(gen[1934]),

			.SELF(gen[1838]),
			.cell_state(gen[1838])
		); 

/******************* CELL 1839 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1839 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1743]),
			.N(gen[1744]),
			.NE(gen[1745]),

			.O(gen[1838]),
			.E(gen[1840]),

			.SO(gen[1933]),
			.S(gen[1934]),
			.SE(gen[1935]),

			.SELF(gen[1839]),
			.cell_state(gen[1839])
		); 

/******************* CELL 1840 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1840 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1744]),
			.N(gen[1745]),
			.NE(gen[1746]),

			.O(gen[1839]),
			.E(gen[1841]),

			.SO(gen[1934]),
			.S(gen[1935]),
			.SE(gen[1936]),

			.SELF(gen[1840]),
			.cell_state(gen[1840])
		); 

/******************* CELL 1841 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1841 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1745]),
			.N(gen[1746]),
			.NE(gen[1747]),

			.O(gen[1840]),
			.E(gen[1842]),

			.SO(gen[1935]),
			.S(gen[1936]),
			.SE(gen[1937]),

			.SELF(gen[1841]),
			.cell_state(gen[1841])
		); 

/******************* CELL 1842 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1842 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1746]),
			.N(gen[1747]),
			.NE(gen[1748]),

			.O(gen[1841]),
			.E(gen[1843]),

			.SO(gen[1936]),
			.S(gen[1937]),
			.SE(gen[1938]),

			.SELF(gen[1842]),
			.cell_state(gen[1842])
		); 

/******************* CELL 1843 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1843 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1747]),
			.N(gen[1748]),
			.NE(gen[1749]),

			.O(gen[1842]),
			.E(gen[1844]),

			.SO(gen[1937]),
			.S(gen[1938]),
			.SE(gen[1939]),

			.SELF(gen[1843]),
			.cell_state(gen[1843])
		); 

/******************* CELL 1844 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1844 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1748]),
			.N(gen[1749]),
			.NE(gen[1750]),

			.O(gen[1843]),
			.E(gen[1845]),

			.SO(gen[1938]),
			.S(gen[1939]),
			.SE(gen[1940]),

			.SELF(gen[1844]),
			.cell_state(gen[1844])
		); 

/******************* CELL 1845 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1845 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1749]),
			.N(gen[1750]),
			.NE(gen[1751]),

			.O(gen[1844]),
			.E(gen[1846]),

			.SO(gen[1939]),
			.S(gen[1940]),
			.SE(gen[1941]),

			.SELF(gen[1845]),
			.cell_state(gen[1845])
		); 

/******************* CELL 1846 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1846 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1750]),
			.N(gen[1751]),
			.NE(gen[1752]),

			.O(gen[1845]),
			.E(gen[1847]),

			.SO(gen[1940]),
			.S(gen[1941]),
			.SE(gen[1942]),

			.SELF(gen[1846]),
			.cell_state(gen[1846])
		); 

/******************* CELL 1847 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1847 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1751]),
			.N(gen[1752]),
			.NE(gen[1753]),

			.O(gen[1846]),
			.E(gen[1848]),

			.SO(gen[1941]),
			.S(gen[1942]),
			.SE(gen[1943]),

			.SELF(gen[1847]),
			.cell_state(gen[1847])
		); 

/******************* CELL 1848 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1848 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1752]),
			.N(gen[1753]),
			.NE(gen[1754]),

			.O(gen[1847]),
			.E(gen[1849]),

			.SO(gen[1942]),
			.S(gen[1943]),
			.SE(gen[1944]),

			.SELF(gen[1848]),
			.cell_state(gen[1848])
		); 

/******************* CELL 1849 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1849 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1753]),
			.N(gen[1754]),
			.NE(gen[1755]),

			.O(gen[1848]),
			.E(gen[1850]),

			.SO(gen[1943]),
			.S(gen[1944]),
			.SE(gen[1945]),

			.SELF(gen[1849]),
			.cell_state(gen[1849])
		); 

/******************* CELL 1850 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1850 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1754]),
			.N(gen[1755]),
			.NE(gen[1756]),

			.O(gen[1849]),
			.E(gen[1851]),

			.SO(gen[1944]),
			.S(gen[1945]),
			.SE(gen[1946]),

			.SELF(gen[1850]),
			.cell_state(gen[1850])
		); 

/******************* CELL 1851 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1851 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1755]),
			.N(gen[1756]),
			.NE(gen[1757]),

			.O(gen[1850]),
			.E(gen[1852]),

			.SO(gen[1945]),
			.S(gen[1946]),
			.SE(gen[1947]),

			.SELF(gen[1851]),
			.cell_state(gen[1851])
		); 

/******************* CELL 1852 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1852 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1756]),
			.N(gen[1757]),
			.NE(gen[1758]),

			.O(gen[1851]),
			.E(gen[1853]),

			.SO(gen[1946]),
			.S(gen[1947]),
			.SE(gen[1948]),

			.SELF(gen[1852]),
			.cell_state(gen[1852])
		); 

/******************* CELL 1853 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1853 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1757]),
			.N(gen[1758]),
			.NE(gen[1759]),

			.O(gen[1852]),
			.E(gen[1854]),

			.SO(gen[1947]),
			.S(gen[1948]),
			.SE(gen[1949]),

			.SELF(gen[1853]),
			.cell_state(gen[1853])
		); 

/******************* CELL 1854 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1854 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1758]),
			.N(gen[1759]),
			.NE(gen[1760]),

			.O(gen[1853]),
			.E(gen[1855]),

			.SO(gen[1948]),
			.S(gen[1949]),
			.SE(gen[1950]),

			.SELF(gen[1854]),
			.cell_state(gen[1854])
		); 

/******************* CELL 1855 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1855 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1759]),
			.N(gen[1760]),
			.NE(gen[1761]),

			.O(gen[1854]),
			.E(gen[1856]),

			.SO(gen[1949]),
			.S(gen[1950]),
			.SE(gen[1951]),

			.SELF(gen[1855]),
			.cell_state(gen[1855])
		); 

/******************* CELL 1856 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1856 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1760]),
			.N(gen[1761]),
			.NE(gen[1762]),

			.O(gen[1855]),
			.E(gen[1857]),

			.SO(gen[1950]),
			.S(gen[1951]),
			.SE(gen[1952]),

			.SELF(gen[1856]),
			.cell_state(gen[1856])
		); 

/******************* CELL 1857 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1857 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1761]),
			.N(gen[1762]),
			.NE(gen[1763]),

			.O(gen[1856]),
			.E(gen[1858]),

			.SO(gen[1951]),
			.S(gen[1952]),
			.SE(gen[1953]),

			.SELF(gen[1857]),
			.cell_state(gen[1857])
		); 

/******************* CELL 1858 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1858 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1762]),
			.N(gen[1763]),
			.NE(gen[1764]),

			.O(gen[1857]),
			.E(gen[1859]),

			.SO(gen[1952]),
			.S(gen[1953]),
			.SE(gen[1954]),

			.SELF(gen[1858]),
			.cell_state(gen[1858])
		); 

/******************* CELL 1859 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1859 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1763]),
			.N(gen[1764]),
			.NE(gen[1765]),

			.O(gen[1858]),
			.E(gen[1860]),

			.SO(gen[1953]),
			.S(gen[1954]),
			.SE(gen[1955]),

			.SELF(gen[1859]),
			.cell_state(gen[1859])
		); 

/******************* CELL 1860 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1860 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1764]),
			.N(gen[1765]),
			.NE(gen[1766]),

			.O(gen[1859]),
			.E(gen[1861]),

			.SO(gen[1954]),
			.S(gen[1955]),
			.SE(gen[1956]),

			.SELF(gen[1860]),
			.cell_state(gen[1860])
		); 

/******************* CELL 1861 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1861 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1765]),
			.N(gen[1766]),
			.NE(gen[1767]),

			.O(gen[1860]),
			.E(gen[1862]),

			.SO(gen[1955]),
			.S(gen[1956]),
			.SE(gen[1957]),

			.SELF(gen[1861]),
			.cell_state(gen[1861])
		); 

/******************* CELL 1862 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1862 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1766]),
			.N(gen[1767]),
			.NE(gen[1768]),

			.O(gen[1861]),
			.E(gen[1863]),

			.SO(gen[1956]),
			.S(gen[1957]),
			.SE(gen[1958]),

			.SELF(gen[1862]),
			.cell_state(gen[1862])
		); 

/******************* CELL 1863 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1863 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1767]),
			.N(gen[1768]),
			.NE(gen[1769]),

			.O(gen[1862]),
			.E(gen[1864]),

			.SO(gen[1957]),
			.S(gen[1958]),
			.SE(gen[1959]),

			.SELF(gen[1863]),
			.cell_state(gen[1863])
		); 

/******************* CELL 1864 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1864 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1768]),
			.N(gen[1769]),
			.NE(gen[1770]),

			.O(gen[1863]),
			.E(gen[1865]),

			.SO(gen[1958]),
			.S(gen[1959]),
			.SE(gen[1960]),

			.SELF(gen[1864]),
			.cell_state(gen[1864])
		); 

/******************* CELL 1865 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1865 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1769]),
			.N(gen[1770]),
			.NE(gen[1771]),

			.O(gen[1864]),
			.E(gen[1866]),

			.SO(gen[1959]),
			.S(gen[1960]),
			.SE(gen[1961]),

			.SELF(gen[1865]),
			.cell_state(gen[1865])
		); 

/******************* CELL 1866 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1866 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1770]),
			.N(gen[1771]),
			.NE(gen[1772]),

			.O(gen[1865]),
			.E(gen[1867]),

			.SO(gen[1960]),
			.S(gen[1961]),
			.SE(gen[1962]),

			.SELF(gen[1866]),
			.cell_state(gen[1866])
		); 

/******************* CELL 1867 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1867 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1771]),
			.N(gen[1772]),
			.NE(gen[1773]),

			.O(gen[1866]),
			.E(gen[1868]),

			.SO(gen[1961]),
			.S(gen[1962]),
			.SE(gen[1963]),

			.SELF(gen[1867]),
			.cell_state(gen[1867])
		); 

/******************* CELL 1868 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1868 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1772]),
			.N(gen[1773]),
			.NE(gen[1774]),

			.O(gen[1867]),
			.E(gen[1869]),

			.SO(gen[1962]),
			.S(gen[1963]),
			.SE(gen[1964]),

			.SELF(gen[1868]),
			.cell_state(gen[1868])
		); 

/******************* CELL 1869 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1869 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1773]),
			.N(gen[1774]),
			.NE(gen[1775]),

			.O(gen[1868]),
			.E(gen[1870]),

			.SO(gen[1963]),
			.S(gen[1964]),
			.SE(gen[1965]),

			.SELF(gen[1869]),
			.cell_state(gen[1869])
		); 

/******************* CELL 1870 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1870 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1774]),
			.N(gen[1775]),
			.NE(gen[1776]),

			.O(gen[1869]),
			.E(gen[1871]),

			.SO(gen[1964]),
			.S(gen[1965]),
			.SE(gen[1966]),

			.SELF(gen[1870]),
			.cell_state(gen[1870])
		); 

/******************* CELL 1871 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1871 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1775]),
			.N(gen[1776]),
			.NE(gen[1777]),

			.O(gen[1870]),
			.E(gen[1872]),

			.SO(gen[1965]),
			.S(gen[1966]),
			.SE(gen[1967]),

			.SELF(gen[1871]),
			.cell_state(gen[1871])
		); 

/******************* CELL 1872 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1872 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1776]),
			.N(gen[1777]),
			.NE(gen[1778]),

			.O(gen[1871]),
			.E(gen[1873]),

			.SO(gen[1966]),
			.S(gen[1967]),
			.SE(gen[1968]),

			.SELF(gen[1872]),
			.cell_state(gen[1872])
		); 

/******************* CELL 1873 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1873 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1777]),
			.N(gen[1778]),
			.NE(gen[1779]),

			.O(gen[1872]),
			.E(gen[1874]),

			.SO(gen[1967]),
			.S(gen[1968]),
			.SE(gen[1969]),

			.SELF(gen[1873]),
			.cell_state(gen[1873])
		); 

/******************* CELL 1874 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1874 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1778]),
			.N(gen[1779]),
			.NE(gen[1780]),

			.O(gen[1873]),
			.E(gen[1875]),

			.SO(gen[1968]),
			.S(gen[1969]),
			.SE(gen[1970]),

			.SELF(gen[1874]),
			.cell_state(gen[1874])
		); 

/******************* CELL 1875 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1875 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1779]),
			.N(gen[1780]),
			.NE(gen[1781]),

			.O(gen[1874]),
			.E(gen[1876]),

			.SO(gen[1969]),
			.S(gen[1970]),
			.SE(gen[1971]),

			.SELF(gen[1875]),
			.cell_state(gen[1875])
		); 

/******************* CELL 1876 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1876 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1780]),
			.N(gen[1781]),
			.NE(gen[1782]),

			.O(gen[1875]),
			.E(gen[1877]),

			.SO(gen[1970]),
			.S(gen[1971]),
			.SE(gen[1972]),

			.SELF(gen[1876]),
			.cell_state(gen[1876])
		); 

/******************* CELL 1877 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1877 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1781]),
			.N(gen[1782]),
			.NE(gen[1783]),

			.O(gen[1876]),
			.E(gen[1878]),

			.SO(gen[1971]),
			.S(gen[1972]),
			.SE(gen[1973]),

			.SELF(gen[1877]),
			.cell_state(gen[1877])
		); 

/******************* CELL 1878 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1878 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1782]),
			.N(gen[1783]),
			.NE(gen[1784]),

			.O(gen[1877]),
			.E(gen[1879]),

			.SO(gen[1972]),
			.S(gen[1973]),
			.SE(gen[1974]),

			.SELF(gen[1878]),
			.cell_state(gen[1878])
		); 

/******************* CELL 1879 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1879 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1783]),
			.N(gen[1784]),
			.NE(gen[1785]),

			.O(gen[1878]),
			.E(gen[1880]),

			.SO(gen[1973]),
			.S(gen[1974]),
			.SE(gen[1975]),

			.SELF(gen[1879]),
			.cell_state(gen[1879])
		); 

/******************* CELL 1880 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1880 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1784]),
			.N(gen[1785]),
			.NE(gen[1786]),

			.O(gen[1879]),
			.E(gen[1881]),

			.SO(gen[1974]),
			.S(gen[1975]),
			.SE(gen[1976]),

			.SELF(gen[1880]),
			.cell_state(gen[1880])
		); 

/******************* CELL 1881 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1881 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1785]),
			.N(gen[1786]),
			.NE(gen[1787]),

			.O(gen[1880]),
			.E(gen[1882]),

			.SO(gen[1975]),
			.S(gen[1976]),
			.SE(gen[1977]),

			.SELF(gen[1881]),
			.cell_state(gen[1881])
		); 

/******************* CELL 1882 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1882 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1786]),
			.N(gen[1787]),
			.NE(gen[1788]),

			.O(gen[1881]),
			.E(gen[1883]),

			.SO(gen[1976]),
			.S(gen[1977]),
			.SE(gen[1978]),

			.SELF(gen[1882]),
			.cell_state(gen[1882])
		); 

/******************* CELL 1883 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1883 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1787]),
			.N(gen[1788]),
			.NE(gen[1789]),

			.O(gen[1882]),
			.E(gen[1884]),

			.SO(gen[1977]),
			.S(gen[1978]),
			.SE(gen[1979]),

			.SELF(gen[1883]),
			.cell_state(gen[1883])
		); 

/******************* CELL 1884 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1884 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1788]),
			.N(gen[1789]),
			.NE(gen[1790]),

			.O(gen[1883]),
			.E(gen[1885]),

			.SO(gen[1978]),
			.S(gen[1979]),
			.SE(gen[1980]),

			.SELF(gen[1884]),
			.cell_state(gen[1884])
		); 

/******************* CELL 1885 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1885 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1789]),
			.N(gen[1790]),
			.NE(gen[1791]),

			.O(gen[1884]),
			.E(gen[1886]),

			.SO(gen[1979]),
			.S(gen[1980]),
			.SE(gen[1981]),

			.SELF(gen[1885]),
			.cell_state(gen[1885])
		); 

/******************* CELL 1886 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1886 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1790]),
			.N(gen[1791]),
			.NE(gen[1792]),

			.O(gen[1885]),
			.E(gen[1887]),

			.SO(gen[1980]),
			.S(gen[1981]),
			.SE(gen[1982]),

			.SELF(gen[1886]),
			.cell_state(gen[1886])
		); 

/******************* CELL 1887 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1887 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1791]),
			.N(gen[1792]),
			.NE(gen[1793]),

			.O(gen[1886]),
			.E(gen[1888]),

			.SO(gen[1981]),
			.S(gen[1982]),
			.SE(gen[1983]),

			.SELF(gen[1887]),
			.cell_state(gen[1887])
		); 

/******************* CELL 1888 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1888 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1792]),
			.N(gen[1793]),
			.NE(gen[1794]),

			.O(gen[1887]),
			.E(gen[1889]),

			.SO(gen[1982]),
			.S(gen[1983]),
			.SE(gen[1984]),

			.SELF(gen[1888]),
			.cell_state(gen[1888])
		); 

/******************* CELL 1889 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1889 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1793]),
			.N(gen[1794]),
			.NE(gen[1795]),

			.O(gen[1888]),
			.E(gen[1890]),

			.SO(gen[1983]),
			.S(gen[1984]),
			.SE(gen[1985]),

			.SELF(gen[1889]),
			.cell_state(gen[1889])
		); 

/******************* CELL 1890 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1890 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1794]),
			.N(gen[1795]),
			.NE(gen[1796]),

			.O(gen[1889]),
			.E(gen[1891]),

			.SO(gen[1984]),
			.S(gen[1985]),
			.SE(gen[1986]),

			.SELF(gen[1890]),
			.cell_state(gen[1890])
		); 

/******************* CELL 1891 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1891 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1795]),
			.N(gen[1796]),
			.NE(gen[1797]),

			.O(gen[1890]),
			.E(gen[1892]),

			.SO(gen[1985]),
			.S(gen[1986]),
			.SE(gen[1987]),

			.SELF(gen[1891]),
			.cell_state(gen[1891])
		); 

/******************* CELL 1892 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1892 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1796]),
			.N(gen[1797]),
			.NE(gen[1798]),

			.O(gen[1891]),
			.E(gen[1893]),

			.SO(gen[1986]),
			.S(gen[1987]),
			.SE(gen[1988]),

			.SELF(gen[1892]),
			.cell_state(gen[1892])
		); 

/******************* CELL 1893 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1893 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1797]),
			.N(gen[1798]),
			.NE(gen[1799]),

			.O(gen[1892]),
			.E(gen[1894]),

			.SO(gen[1987]),
			.S(gen[1988]),
			.SE(gen[1989]),

			.SELF(gen[1893]),
			.cell_state(gen[1893])
		); 

/******************* CELL 1894 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1894 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1798]),
			.N(gen[1799]),
			.NE(gen[1800]),

			.O(gen[1893]),
			.E(gen[1895]),

			.SO(gen[1988]),
			.S(gen[1989]),
			.SE(gen[1990]),

			.SELF(gen[1894]),
			.cell_state(gen[1894])
		); 

/******************* CELL 1895 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1895 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1799]),
			.N(gen[1800]),
			.NE(gen[1801]),

			.O(gen[1894]),
			.E(gen[1896]),

			.SO(gen[1989]),
			.S(gen[1990]),
			.SE(gen[1991]),

			.SELF(gen[1895]),
			.cell_state(gen[1895])
		); 

/******************* CELL 1896 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1896 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1800]),
			.N(gen[1801]),
			.NE(gen[1802]),

			.O(gen[1895]),
			.E(gen[1897]),

			.SO(gen[1990]),
			.S(gen[1991]),
			.SE(gen[1992]),

			.SELF(gen[1896]),
			.cell_state(gen[1896])
		); 

/******************* CELL 1897 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1897 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1801]),
			.N(gen[1802]),
			.NE(gen[1803]),

			.O(gen[1896]),
			.E(gen[1898]),

			.SO(gen[1991]),
			.S(gen[1992]),
			.SE(gen[1993]),

			.SELF(gen[1897]),
			.cell_state(gen[1897])
		); 

/******************* CELL 1898 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1898 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1802]),
			.N(gen[1803]),
			.NE(gen[1804]),

			.O(gen[1897]),
			.E(gen[1899]),

			.SO(gen[1992]),
			.S(gen[1993]),
			.SE(gen[1994]),

			.SELF(gen[1898]),
			.cell_state(gen[1898])
		); 

/******************* CELL 1899 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1899 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1803]),
			.N(gen[1804]),
			.NE(gen[1803]),

			.O(gen[1898]),
			.E(gen[1898]),

			.SO(gen[1993]),
			.S(gen[1994]),
			.SE(gen[1993]),

			.SELF(gen[1899]),
			.cell_state(gen[1899])
		); 

/******************* CELL 1900 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1900 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1806]),
			.N(gen[1805]),
			.NE(gen[1806]),

			.O(gen[1901]),
			.E(gen[1901]),

			.SO(gen[1996]),
			.S(gen[1995]),
			.SE(gen[1996]),

			.SELF(gen[1900]),
			.cell_state(gen[1900])
		); 

/******************* CELL 1901 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1901 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1805]),
			.N(gen[1806]),
			.NE(gen[1807]),

			.O(gen[1900]),
			.E(gen[1902]),

			.SO(gen[1995]),
			.S(gen[1996]),
			.SE(gen[1997]),

			.SELF(gen[1901]),
			.cell_state(gen[1901])
		); 

/******************* CELL 1902 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1902 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1806]),
			.N(gen[1807]),
			.NE(gen[1808]),

			.O(gen[1901]),
			.E(gen[1903]),

			.SO(gen[1996]),
			.S(gen[1997]),
			.SE(gen[1998]),

			.SELF(gen[1902]),
			.cell_state(gen[1902])
		); 

/******************* CELL 1903 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1903 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1807]),
			.N(gen[1808]),
			.NE(gen[1809]),

			.O(gen[1902]),
			.E(gen[1904]),

			.SO(gen[1997]),
			.S(gen[1998]),
			.SE(gen[1999]),

			.SELF(gen[1903]),
			.cell_state(gen[1903])
		); 

/******************* CELL 1904 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1904 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1808]),
			.N(gen[1809]),
			.NE(gen[1810]),

			.O(gen[1903]),
			.E(gen[1905]),

			.SO(gen[1998]),
			.S(gen[1999]),
			.SE(gen[2000]),

			.SELF(gen[1904]),
			.cell_state(gen[1904])
		); 

/******************* CELL 1905 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1905 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1809]),
			.N(gen[1810]),
			.NE(gen[1811]),

			.O(gen[1904]),
			.E(gen[1906]),

			.SO(gen[1999]),
			.S(gen[2000]),
			.SE(gen[2001]),

			.SELF(gen[1905]),
			.cell_state(gen[1905])
		); 

/******************* CELL 1906 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1906 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1810]),
			.N(gen[1811]),
			.NE(gen[1812]),

			.O(gen[1905]),
			.E(gen[1907]),

			.SO(gen[2000]),
			.S(gen[2001]),
			.SE(gen[2002]),

			.SELF(gen[1906]),
			.cell_state(gen[1906])
		); 

/******************* CELL 1907 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1907 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1811]),
			.N(gen[1812]),
			.NE(gen[1813]),

			.O(gen[1906]),
			.E(gen[1908]),

			.SO(gen[2001]),
			.S(gen[2002]),
			.SE(gen[2003]),

			.SELF(gen[1907]),
			.cell_state(gen[1907])
		); 

/******************* CELL 1908 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1908 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1812]),
			.N(gen[1813]),
			.NE(gen[1814]),

			.O(gen[1907]),
			.E(gen[1909]),

			.SO(gen[2002]),
			.S(gen[2003]),
			.SE(gen[2004]),

			.SELF(gen[1908]),
			.cell_state(gen[1908])
		); 

/******************* CELL 1909 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1909 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1813]),
			.N(gen[1814]),
			.NE(gen[1815]),

			.O(gen[1908]),
			.E(gen[1910]),

			.SO(gen[2003]),
			.S(gen[2004]),
			.SE(gen[2005]),

			.SELF(gen[1909]),
			.cell_state(gen[1909])
		); 

/******************* CELL 1910 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1910 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1814]),
			.N(gen[1815]),
			.NE(gen[1816]),

			.O(gen[1909]),
			.E(gen[1911]),

			.SO(gen[2004]),
			.S(gen[2005]),
			.SE(gen[2006]),

			.SELF(gen[1910]),
			.cell_state(gen[1910])
		); 

/******************* CELL 1911 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1911 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1815]),
			.N(gen[1816]),
			.NE(gen[1817]),

			.O(gen[1910]),
			.E(gen[1912]),

			.SO(gen[2005]),
			.S(gen[2006]),
			.SE(gen[2007]),

			.SELF(gen[1911]),
			.cell_state(gen[1911])
		); 

/******************* CELL 1912 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1912 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1816]),
			.N(gen[1817]),
			.NE(gen[1818]),

			.O(gen[1911]),
			.E(gen[1913]),

			.SO(gen[2006]),
			.S(gen[2007]),
			.SE(gen[2008]),

			.SELF(gen[1912]),
			.cell_state(gen[1912])
		); 

/******************* CELL 1913 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1913 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1817]),
			.N(gen[1818]),
			.NE(gen[1819]),

			.O(gen[1912]),
			.E(gen[1914]),

			.SO(gen[2007]),
			.S(gen[2008]),
			.SE(gen[2009]),

			.SELF(gen[1913]),
			.cell_state(gen[1913])
		); 

/******************* CELL 1914 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1914 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1818]),
			.N(gen[1819]),
			.NE(gen[1820]),

			.O(gen[1913]),
			.E(gen[1915]),

			.SO(gen[2008]),
			.S(gen[2009]),
			.SE(gen[2010]),

			.SELF(gen[1914]),
			.cell_state(gen[1914])
		); 

/******************* CELL 1915 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1915 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1819]),
			.N(gen[1820]),
			.NE(gen[1821]),

			.O(gen[1914]),
			.E(gen[1916]),

			.SO(gen[2009]),
			.S(gen[2010]),
			.SE(gen[2011]),

			.SELF(gen[1915]),
			.cell_state(gen[1915])
		); 

/******************* CELL 1916 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1916 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1820]),
			.N(gen[1821]),
			.NE(gen[1822]),

			.O(gen[1915]),
			.E(gen[1917]),

			.SO(gen[2010]),
			.S(gen[2011]),
			.SE(gen[2012]),

			.SELF(gen[1916]),
			.cell_state(gen[1916])
		); 

/******************* CELL 1917 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1917 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1821]),
			.N(gen[1822]),
			.NE(gen[1823]),

			.O(gen[1916]),
			.E(gen[1918]),

			.SO(gen[2011]),
			.S(gen[2012]),
			.SE(gen[2013]),

			.SELF(gen[1917]),
			.cell_state(gen[1917])
		); 

/******************* CELL 1918 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1918 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1822]),
			.N(gen[1823]),
			.NE(gen[1824]),

			.O(gen[1917]),
			.E(gen[1919]),

			.SO(gen[2012]),
			.S(gen[2013]),
			.SE(gen[2014]),

			.SELF(gen[1918]),
			.cell_state(gen[1918])
		); 

/******************* CELL 1919 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1919 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1823]),
			.N(gen[1824]),
			.NE(gen[1825]),

			.O(gen[1918]),
			.E(gen[1920]),

			.SO(gen[2013]),
			.S(gen[2014]),
			.SE(gen[2015]),

			.SELF(gen[1919]),
			.cell_state(gen[1919])
		); 

/******************* CELL 1920 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1920 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1824]),
			.N(gen[1825]),
			.NE(gen[1826]),

			.O(gen[1919]),
			.E(gen[1921]),

			.SO(gen[2014]),
			.S(gen[2015]),
			.SE(gen[2016]),

			.SELF(gen[1920]),
			.cell_state(gen[1920])
		); 

/******************* CELL 1921 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1921 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1825]),
			.N(gen[1826]),
			.NE(gen[1827]),

			.O(gen[1920]),
			.E(gen[1922]),

			.SO(gen[2015]),
			.S(gen[2016]),
			.SE(gen[2017]),

			.SELF(gen[1921]),
			.cell_state(gen[1921])
		); 

/******************* CELL 1922 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1922 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1826]),
			.N(gen[1827]),
			.NE(gen[1828]),

			.O(gen[1921]),
			.E(gen[1923]),

			.SO(gen[2016]),
			.S(gen[2017]),
			.SE(gen[2018]),

			.SELF(gen[1922]),
			.cell_state(gen[1922])
		); 

/******************* CELL 1923 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1923 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1827]),
			.N(gen[1828]),
			.NE(gen[1829]),

			.O(gen[1922]),
			.E(gen[1924]),

			.SO(gen[2017]),
			.S(gen[2018]),
			.SE(gen[2019]),

			.SELF(gen[1923]),
			.cell_state(gen[1923])
		); 

/******************* CELL 1924 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1924 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1828]),
			.N(gen[1829]),
			.NE(gen[1830]),

			.O(gen[1923]),
			.E(gen[1925]),

			.SO(gen[2018]),
			.S(gen[2019]),
			.SE(gen[2020]),

			.SELF(gen[1924]),
			.cell_state(gen[1924])
		); 

/******************* CELL 1925 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1925 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1829]),
			.N(gen[1830]),
			.NE(gen[1831]),

			.O(gen[1924]),
			.E(gen[1926]),

			.SO(gen[2019]),
			.S(gen[2020]),
			.SE(gen[2021]),

			.SELF(gen[1925]),
			.cell_state(gen[1925])
		); 

/******************* CELL 1926 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1926 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1830]),
			.N(gen[1831]),
			.NE(gen[1832]),

			.O(gen[1925]),
			.E(gen[1927]),

			.SO(gen[2020]),
			.S(gen[2021]),
			.SE(gen[2022]),

			.SELF(gen[1926]),
			.cell_state(gen[1926])
		); 

/******************* CELL 1927 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1927 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1831]),
			.N(gen[1832]),
			.NE(gen[1833]),

			.O(gen[1926]),
			.E(gen[1928]),

			.SO(gen[2021]),
			.S(gen[2022]),
			.SE(gen[2023]),

			.SELF(gen[1927]),
			.cell_state(gen[1927])
		); 

/******************* CELL 1928 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1928 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1832]),
			.N(gen[1833]),
			.NE(gen[1834]),

			.O(gen[1927]),
			.E(gen[1929]),

			.SO(gen[2022]),
			.S(gen[2023]),
			.SE(gen[2024]),

			.SELF(gen[1928]),
			.cell_state(gen[1928])
		); 

/******************* CELL 1929 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1929 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1833]),
			.N(gen[1834]),
			.NE(gen[1835]),

			.O(gen[1928]),
			.E(gen[1930]),

			.SO(gen[2023]),
			.S(gen[2024]),
			.SE(gen[2025]),

			.SELF(gen[1929]),
			.cell_state(gen[1929])
		); 

/******************* CELL 1930 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1930 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1834]),
			.N(gen[1835]),
			.NE(gen[1836]),

			.O(gen[1929]),
			.E(gen[1931]),

			.SO(gen[2024]),
			.S(gen[2025]),
			.SE(gen[2026]),

			.SELF(gen[1930]),
			.cell_state(gen[1930])
		); 

/******************* CELL 1931 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1931 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1835]),
			.N(gen[1836]),
			.NE(gen[1837]),

			.O(gen[1930]),
			.E(gen[1932]),

			.SO(gen[2025]),
			.S(gen[2026]),
			.SE(gen[2027]),

			.SELF(gen[1931]),
			.cell_state(gen[1931])
		); 

/******************* CELL 1932 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1932 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1836]),
			.N(gen[1837]),
			.NE(gen[1838]),

			.O(gen[1931]),
			.E(gen[1933]),

			.SO(gen[2026]),
			.S(gen[2027]),
			.SE(gen[2028]),

			.SELF(gen[1932]),
			.cell_state(gen[1932])
		); 

/******************* CELL 1933 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1933 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1837]),
			.N(gen[1838]),
			.NE(gen[1839]),

			.O(gen[1932]),
			.E(gen[1934]),

			.SO(gen[2027]),
			.S(gen[2028]),
			.SE(gen[2029]),

			.SELF(gen[1933]),
			.cell_state(gen[1933])
		); 

/******************* CELL 1934 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1934 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1838]),
			.N(gen[1839]),
			.NE(gen[1840]),

			.O(gen[1933]),
			.E(gen[1935]),

			.SO(gen[2028]),
			.S(gen[2029]),
			.SE(gen[2030]),

			.SELF(gen[1934]),
			.cell_state(gen[1934])
		); 

/******************* CELL 1935 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1935 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1839]),
			.N(gen[1840]),
			.NE(gen[1841]),

			.O(gen[1934]),
			.E(gen[1936]),

			.SO(gen[2029]),
			.S(gen[2030]),
			.SE(gen[2031]),

			.SELF(gen[1935]),
			.cell_state(gen[1935])
		); 

/******************* CELL 1936 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1936 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1840]),
			.N(gen[1841]),
			.NE(gen[1842]),

			.O(gen[1935]),
			.E(gen[1937]),

			.SO(gen[2030]),
			.S(gen[2031]),
			.SE(gen[2032]),

			.SELF(gen[1936]),
			.cell_state(gen[1936])
		); 

/******************* CELL 1937 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1937 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1841]),
			.N(gen[1842]),
			.NE(gen[1843]),

			.O(gen[1936]),
			.E(gen[1938]),

			.SO(gen[2031]),
			.S(gen[2032]),
			.SE(gen[2033]),

			.SELF(gen[1937]),
			.cell_state(gen[1937])
		); 

/******************* CELL 1938 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1938 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1842]),
			.N(gen[1843]),
			.NE(gen[1844]),

			.O(gen[1937]),
			.E(gen[1939]),

			.SO(gen[2032]),
			.S(gen[2033]),
			.SE(gen[2034]),

			.SELF(gen[1938]),
			.cell_state(gen[1938])
		); 

/******************* CELL 1939 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1939 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1843]),
			.N(gen[1844]),
			.NE(gen[1845]),

			.O(gen[1938]),
			.E(gen[1940]),

			.SO(gen[2033]),
			.S(gen[2034]),
			.SE(gen[2035]),

			.SELF(gen[1939]),
			.cell_state(gen[1939])
		); 

/******************* CELL 1940 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1940 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1844]),
			.N(gen[1845]),
			.NE(gen[1846]),

			.O(gen[1939]),
			.E(gen[1941]),

			.SO(gen[2034]),
			.S(gen[2035]),
			.SE(gen[2036]),

			.SELF(gen[1940]),
			.cell_state(gen[1940])
		); 

/******************* CELL 1941 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1941 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1845]),
			.N(gen[1846]),
			.NE(gen[1847]),

			.O(gen[1940]),
			.E(gen[1942]),

			.SO(gen[2035]),
			.S(gen[2036]),
			.SE(gen[2037]),

			.SELF(gen[1941]),
			.cell_state(gen[1941])
		); 

/******************* CELL 1942 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1942 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1846]),
			.N(gen[1847]),
			.NE(gen[1848]),

			.O(gen[1941]),
			.E(gen[1943]),

			.SO(gen[2036]),
			.S(gen[2037]),
			.SE(gen[2038]),

			.SELF(gen[1942]),
			.cell_state(gen[1942])
		); 

/******************* CELL 1943 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1943 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1847]),
			.N(gen[1848]),
			.NE(gen[1849]),

			.O(gen[1942]),
			.E(gen[1944]),

			.SO(gen[2037]),
			.S(gen[2038]),
			.SE(gen[2039]),

			.SELF(gen[1943]),
			.cell_state(gen[1943])
		); 

/******************* CELL 1944 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1944 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1848]),
			.N(gen[1849]),
			.NE(gen[1850]),

			.O(gen[1943]),
			.E(gen[1945]),

			.SO(gen[2038]),
			.S(gen[2039]),
			.SE(gen[2040]),

			.SELF(gen[1944]),
			.cell_state(gen[1944])
		); 

/******************* CELL 1945 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1945 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1849]),
			.N(gen[1850]),
			.NE(gen[1851]),

			.O(gen[1944]),
			.E(gen[1946]),

			.SO(gen[2039]),
			.S(gen[2040]),
			.SE(gen[2041]),

			.SELF(gen[1945]),
			.cell_state(gen[1945])
		); 

/******************* CELL 1946 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1946 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1850]),
			.N(gen[1851]),
			.NE(gen[1852]),

			.O(gen[1945]),
			.E(gen[1947]),

			.SO(gen[2040]),
			.S(gen[2041]),
			.SE(gen[2042]),

			.SELF(gen[1946]),
			.cell_state(gen[1946])
		); 

/******************* CELL 1947 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1947 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1851]),
			.N(gen[1852]),
			.NE(gen[1853]),

			.O(gen[1946]),
			.E(gen[1948]),

			.SO(gen[2041]),
			.S(gen[2042]),
			.SE(gen[2043]),

			.SELF(gen[1947]),
			.cell_state(gen[1947])
		); 

/******************* CELL 1948 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1948 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1852]),
			.N(gen[1853]),
			.NE(gen[1854]),

			.O(gen[1947]),
			.E(gen[1949]),

			.SO(gen[2042]),
			.S(gen[2043]),
			.SE(gen[2044]),

			.SELF(gen[1948]),
			.cell_state(gen[1948])
		); 

/******************* CELL 1949 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1949 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1853]),
			.N(gen[1854]),
			.NE(gen[1855]),

			.O(gen[1948]),
			.E(gen[1950]),

			.SO(gen[2043]),
			.S(gen[2044]),
			.SE(gen[2045]),

			.SELF(gen[1949]),
			.cell_state(gen[1949])
		); 

/******************* CELL 1950 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1950 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1854]),
			.N(gen[1855]),
			.NE(gen[1856]),

			.O(gen[1949]),
			.E(gen[1951]),

			.SO(gen[2044]),
			.S(gen[2045]),
			.SE(gen[2046]),

			.SELF(gen[1950]),
			.cell_state(gen[1950])
		); 

/******************* CELL 1951 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1951 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1855]),
			.N(gen[1856]),
			.NE(gen[1857]),

			.O(gen[1950]),
			.E(gen[1952]),

			.SO(gen[2045]),
			.S(gen[2046]),
			.SE(gen[2047]),

			.SELF(gen[1951]),
			.cell_state(gen[1951])
		); 

/******************* CELL 1952 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1952 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1856]),
			.N(gen[1857]),
			.NE(gen[1858]),

			.O(gen[1951]),
			.E(gen[1953]),

			.SO(gen[2046]),
			.S(gen[2047]),
			.SE(gen[2048]),

			.SELF(gen[1952]),
			.cell_state(gen[1952])
		); 

/******************* CELL 1953 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1953 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1857]),
			.N(gen[1858]),
			.NE(gen[1859]),

			.O(gen[1952]),
			.E(gen[1954]),

			.SO(gen[2047]),
			.S(gen[2048]),
			.SE(gen[2049]),

			.SELF(gen[1953]),
			.cell_state(gen[1953])
		); 

/******************* CELL 1954 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1954 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1858]),
			.N(gen[1859]),
			.NE(gen[1860]),

			.O(gen[1953]),
			.E(gen[1955]),

			.SO(gen[2048]),
			.S(gen[2049]),
			.SE(gen[2050]),

			.SELF(gen[1954]),
			.cell_state(gen[1954])
		); 

/******************* CELL 1955 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1955 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1859]),
			.N(gen[1860]),
			.NE(gen[1861]),

			.O(gen[1954]),
			.E(gen[1956]),

			.SO(gen[2049]),
			.S(gen[2050]),
			.SE(gen[2051]),

			.SELF(gen[1955]),
			.cell_state(gen[1955])
		); 

/******************* CELL 1956 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1956 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1860]),
			.N(gen[1861]),
			.NE(gen[1862]),

			.O(gen[1955]),
			.E(gen[1957]),

			.SO(gen[2050]),
			.S(gen[2051]),
			.SE(gen[2052]),

			.SELF(gen[1956]),
			.cell_state(gen[1956])
		); 

/******************* CELL 1957 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1957 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1861]),
			.N(gen[1862]),
			.NE(gen[1863]),

			.O(gen[1956]),
			.E(gen[1958]),

			.SO(gen[2051]),
			.S(gen[2052]),
			.SE(gen[2053]),

			.SELF(gen[1957]),
			.cell_state(gen[1957])
		); 

/******************* CELL 1958 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1958 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1862]),
			.N(gen[1863]),
			.NE(gen[1864]),

			.O(gen[1957]),
			.E(gen[1959]),

			.SO(gen[2052]),
			.S(gen[2053]),
			.SE(gen[2054]),

			.SELF(gen[1958]),
			.cell_state(gen[1958])
		); 

/******************* CELL 1959 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1959 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1863]),
			.N(gen[1864]),
			.NE(gen[1865]),

			.O(gen[1958]),
			.E(gen[1960]),

			.SO(gen[2053]),
			.S(gen[2054]),
			.SE(gen[2055]),

			.SELF(gen[1959]),
			.cell_state(gen[1959])
		); 

/******************* CELL 1960 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1960 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1864]),
			.N(gen[1865]),
			.NE(gen[1866]),

			.O(gen[1959]),
			.E(gen[1961]),

			.SO(gen[2054]),
			.S(gen[2055]),
			.SE(gen[2056]),

			.SELF(gen[1960]),
			.cell_state(gen[1960])
		); 

/******************* CELL 1961 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1961 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1865]),
			.N(gen[1866]),
			.NE(gen[1867]),

			.O(gen[1960]),
			.E(gen[1962]),

			.SO(gen[2055]),
			.S(gen[2056]),
			.SE(gen[2057]),

			.SELF(gen[1961]),
			.cell_state(gen[1961])
		); 

/******************* CELL 1962 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1962 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1866]),
			.N(gen[1867]),
			.NE(gen[1868]),

			.O(gen[1961]),
			.E(gen[1963]),

			.SO(gen[2056]),
			.S(gen[2057]),
			.SE(gen[2058]),

			.SELF(gen[1962]),
			.cell_state(gen[1962])
		); 

/******************* CELL 1963 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1963 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1867]),
			.N(gen[1868]),
			.NE(gen[1869]),

			.O(gen[1962]),
			.E(gen[1964]),

			.SO(gen[2057]),
			.S(gen[2058]),
			.SE(gen[2059]),

			.SELF(gen[1963]),
			.cell_state(gen[1963])
		); 

/******************* CELL 1964 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1964 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1868]),
			.N(gen[1869]),
			.NE(gen[1870]),

			.O(gen[1963]),
			.E(gen[1965]),

			.SO(gen[2058]),
			.S(gen[2059]),
			.SE(gen[2060]),

			.SELF(gen[1964]),
			.cell_state(gen[1964])
		); 

/******************* CELL 1965 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1965 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1869]),
			.N(gen[1870]),
			.NE(gen[1871]),

			.O(gen[1964]),
			.E(gen[1966]),

			.SO(gen[2059]),
			.S(gen[2060]),
			.SE(gen[2061]),

			.SELF(gen[1965]),
			.cell_state(gen[1965])
		); 

/******************* CELL 1966 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1966 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1870]),
			.N(gen[1871]),
			.NE(gen[1872]),

			.O(gen[1965]),
			.E(gen[1967]),

			.SO(gen[2060]),
			.S(gen[2061]),
			.SE(gen[2062]),

			.SELF(gen[1966]),
			.cell_state(gen[1966])
		); 

/******************* CELL 1967 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1967 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1871]),
			.N(gen[1872]),
			.NE(gen[1873]),

			.O(gen[1966]),
			.E(gen[1968]),

			.SO(gen[2061]),
			.S(gen[2062]),
			.SE(gen[2063]),

			.SELF(gen[1967]),
			.cell_state(gen[1967])
		); 

/******************* CELL 1968 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1968 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1872]),
			.N(gen[1873]),
			.NE(gen[1874]),

			.O(gen[1967]),
			.E(gen[1969]),

			.SO(gen[2062]),
			.S(gen[2063]),
			.SE(gen[2064]),

			.SELF(gen[1968]),
			.cell_state(gen[1968])
		); 

/******************* CELL 1969 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1969 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1873]),
			.N(gen[1874]),
			.NE(gen[1875]),

			.O(gen[1968]),
			.E(gen[1970]),

			.SO(gen[2063]),
			.S(gen[2064]),
			.SE(gen[2065]),

			.SELF(gen[1969]),
			.cell_state(gen[1969])
		); 

/******************* CELL 1970 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1970 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1874]),
			.N(gen[1875]),
			.NE(gen[1876]),

			.O(gen[1969]),
			.E(gen[1971]),

			.SO(gen[2064]),
			.S(gen[2065]),
			.SE(gen[2066]),

			.SELF(gen[1970]),
			.cell_state(gen[1970])
		); 

/******************* CELL 1971 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1971 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1875]),
			.N(gen[1876]),
			.NE(gen[1877]),

			.O(gen[1970]),
			.E(gen[1972]),

			.SO(gen[2065]),
			.S(gen[2066]),
			.SE(gen[2067]),

			.SELF(gen[1971]),
			.cell_state(gen[1971])
		); 

/******************* CELL 1972 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1972 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1876]),
			.N(gen[1877]),
			.NE(gen[1878]),

			.O(gen[1971]),
			.E(gen[1973]),

			.SO(gen[2066]),
			.S(gen[2067]),
			.SE(gen[2068]),

			.SELF(gen[1972]),
			.cell_state(gen[1972])
		); 

/******************* CELL 1973 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1973 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1877]),
			.N(gen[1878]),
			.NE(gen[1879]),

			.O(gen[1972]),
			.E(gen[1974]),

			.SO(gen[2067]),
			.S(gen[2068]),
			.SE(gen[2069]),

			.SELF(gen[1973]),
			.cell_state(gen[1973])
		); 

/******************* CELL 1974 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1974 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1878]),
			.N(gen[1879]),
			.NE(gen[1880]),

			.O(gen[1973]),
			.E(gen[1975]),

			.SO(gen[2068]),
			.S(gen[2069]),
			.SE(gen[2070]),

			.SELF(gen[1974]),
			.cell_state(gen[1974])
		); 

/******************* CELL 1975 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1975 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1879]),
			.N(gen[1880]),
			.NE(gen[1881]),

			.O(gen[1974]),
			.E(gen[1976]),

			.SO(gen[2069]),
			.S(gen[2070]),
			.SE(gen[2071]),

			.SELF(gen[1975]),
			.cell_state(gen[1975])
		); 

/******************* CELL 1976 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1976 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1880]),
			.N(gen[1881]),
			.NE(gen[1882]),

			.O(gen[1975]),
			.E(gen[1977]),

			.SO(gen[2070]),
			.S(gen[2071]),
			.SE(gen[2072]),

			.SELF(gen[1976]),
			.cell_state(gen[1976])
		); 

/******************* CELL 1977 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1977 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1881]),
			.N(gen[1882]),
			.NE(gen[1883]),

			.O(gen[1976]),
			.E(gen[1978]),

			.SO(gen[2071]),
			.S(gen[2072]),
			.SE(gen[2073]),

			.SELF(gen[1977]),
			.cell_state(gen[1977])
		); 

/******************* CELL 1978 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1978 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1882]),
			.N(gen[1883]),
			.NE(gen[1884]),

			.O(gen[1977]),
			.E(gen[1979]),

			.SO(gen[2072]),
			.S(gen[2073]),
			.SE(gen[2074]),

			.SELF(gen[1978]),
			.cell_state(gen[1978])
		); 

/******************* CELL 1979 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1979 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1883]),
			.N(gen[1884]),
			.NE(gen[1885]),

			.O(gen[1978]),
			.E(gen[1980]),

			.SO(gen[2073]),
			.S(gen[2074]),
			.SE(gen[2075]),

			.SELF(gen[1979]),
			.cell_state(gen[1979])
		); 

/******************* CELL 1980 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1980 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1884]),
			.N(gen[1885]),
			.NE(gen[1886]),

			.O(gen[1979]),
			.E(gen[1981]),

			.SO(gen[2074]),
			.S(gen[2075]),
			.SE(gen[2076]),

			.SELF(gen[1980]),
			.cell_state(gen[1980])
		); 

/******************* CELL 1981 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1981 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1885]),
			.N(gen[1886]),
			.NE(gen[1887]),

			.O(gen[1980]),
			.E(gen[1982]),

			.SO(gen[2075]),
			.S(gen[2076]),
			.SE(gen[2077]),

			.SELF(gen[1981]),
			.cell_state(gen[1981])
		); 

/******************* CELL 1982 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1982 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1886]),
			.N(gen[1887]),
			.NE(gen[1888]),

			.O(gen[1981]),
			.E(gen[1983]),

			.SO(gen[2076]),
			.S(gen[2077]),
			.SE(gen[2078]),

			.SELF(gen[1982]),
			.cell_state(gen[1982])
		); 

/******************* CELL 1983 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1983 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1887]),
			.N(gen[1888]),
			.NE(gen[1889]),

			.O(gen[1982]),
			.E(gen[1984]),

			.SO(gen[2077]),
			.S(gen[2078]),
			.SE(gen[2079]),

			.SELF(gen[1983]),
			.cell_state(gen[1983])
		); 

/******************* CELL 1984 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1984 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1888]),
			.N(gen[1889]),
			.NE(gen[1890]),

			.O(gen[1983]),
			.E(gen[1985]),

			.SO(gen[2078]),
			.S(gen[2079]),
			.SE(gen[2080]),

			.SELF(gen[1984]),
			.cell_state(gen[1984])
		); 

/******************* CELL 1985 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1985 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1889]),
			.N(gen[1890]),
			.NE(gen[1891]),

			.O(gen[1984]),
			.E(gen[1986]),

			.SO(gen[2079]),
			.S(gen[2080]),
			.SE(gen[2081]),

			.SELF(gen[1985]),
			.cell_state(gen[1985])
		); 

/******************* CELL 1986 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1986 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1890]),
			.N(gen[1891]),
			.NE(gen[1892]),

			.O(gen[1985]),
			.E(gen[1987]),

			.SO(gen[2080]),
			.S(gen[2081]),
			.SE(gen[2082]),

			.SELF(gen[1986]),
			.cell_state(gen[1986])
		); 

/******************* CELL 1987 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1987 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1891]),
			.N(gen[1892]),
			.NE(gen[1893]),

			.O(gen[1986]),
			.E(gen[1988]),

			.SO(gen[2081]),
			.S(gen[2082]),
			.SE(gen[2083]),

			.SELF(gen[1987]),
			.cell_state(gen[1987])
		); 

/******************* CELL 1988 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1988 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1892]),
			.N(gen[1893]),
			.NE(gen[1894]),

			.O(gen[1987]),
			.E(gen[1989]),

			.SO(gen[2082]),
			.S(gen[2083]),
			.SE(gen[2084]),

			.SELF(gen[1988]),
			.cell_state(gen[1988])
		); 

/******************* CELL 1989 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1989 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1893]),
			.N(gen[1894]),
			.NE(gen[1895]),

			.O(gen[1988]),
			.E(gen[1990]),

			.SO(gen[2083]),
			.S(gen[2084]),
			.SE(gen[2085]),

			.SELF(gen[1989]),
			.cell_state(gen[1989])
		); 

/******************* CELL 1990 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1990 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1894]),
			.N(gen[1895]),
			.NE(gen[1896]),

			.O(gen[1989]),
			.E(gen[1991]),

			.SO(gen[2084]),
			.S(gen[2085]),
			.SE(gen[2086]),

			.SELF(gen[1990]),
			.cell_state(gen[1990])
		); 

/******************* CELL 1991 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1991 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1895]),
			.N(gen[1896]),
			.NE(gen[1897]),

			.O(gen[1990]),
			.E(gen[1992]),

			.SO(gen[2085]),
			.S(gen[2086]),
			.SE(gen[2087]),

			.SELF(gen[1991]),
			.cell_state(gen[1991])
		); 

/******************* CELL 1992 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1992 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1896]),
			.N(gen[1897]),
			.NE(gen[1898]),

			.O(gen[1991]),
			.E(gen[1993]),

			.SO(gen[2086]),
			.S(gen[2087]),
			.SE(gen[2088]),

			.SELF(gen[1992]),
			.cell_state(gen[1992])
		); 

/******************* CELL 1993 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1993 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1897]),
			.N(gen[1898]),
			.NE(gen[1899]),

			.O(gen[1992]),
			.E(gen[1994]),

			.SO(gen[2087]),
			.S(gen[2088]),
			.SE(gen[2089]),

			.SELF(gen[1993]),
			.cell_state(gen[1993])
		); 

/******************* CELL 1994 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1994 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1898]),
			.N(gen[1899]),
			.NE(gen[1898]),

			.O(gen[1993]),
			.E(gen[1993]),

			.SO(gen[2088]),
			.S(gen[2089]),
			.SE(gen[2088]),

			.SELF(gen[1994]),
			.cell_state(gen[1994])
		); 

/******************* CELL 1995 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1995 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1901]),
			.N(gen[1900]),
			.NE(gen[1901]),

			.O(gen[1996]),
			.E(gen[1996]),

			.SO(gen[2091]),
			.S(gen[2090]),
			.SE(gen[2091]),

			.SELF(gen[1995]),
			.cell_state(gen[1995])
		); 

/******************* CELL 1996 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1996 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1900]),
			.N(gen[1901]),
			.NE(gen[1902]),

			.O(gen[1995]),
			.E(gen[1997]),

			.SO(gen[2090]),
			.S(gen[2091]),
			.SE(gen[2092]),

			.SELF(gen[1996]),
			.cell_state(gen[1996])
		); 

/******************* CELL 1997 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1997 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1901]),
			.N(gen[1902]),
			.NE(gen[1903]),

			.O(gen[1996]),
			.E(gen[1998]),

			.SO(gen[2091]),
			.S(gen[2092]),
			.SE(gen[2093]),

			.SELF(gen[1997]),
			.cell_state(gen[1997])
		); 

/******************* CELL 1998 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1998 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1902]),
			.N(gen[1903]),
			.NE(gen[1904]),

			.O(gen[1997]),
			.E(gen[1999]),

			.SO(gen[2092]),
			.S(gen[2093]),
			.SE(gen[2094]),

			.SELF(gen[1998]),
			.cell_state(gen[1998])
		); 

/******************* CELL 1999 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1999 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1903]),
			.N(gen[1904]),
			.NE(gen[1905]),

			.O(gen[1998]),
			.E(gen[2000]),

			.SO(gen[2093]),
			.S(gen[2094]),
			.SE(gen[2095]),

			.SELF(gen[1999]),
			.cell_state(gen[1999])
		); 

/******************* CELL 2000 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2000 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1904]),
			.N(gen[1905]),
			.NE(gen[1906]),

			.O(gen[1999]),
			.E(gen[2001]),

			.SO(gen[2094]),
			.S(gen[2095]),
			.SE(gen[2096]),

			.SELF(gen[2000]),
			.cell_state(gen[2000])
		); 

/******************* CELL 2001 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2001 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1905]),
			.N(gen[1906]),
			.NE(gen[1907]),

			.O(gen[2000]),
			.E(gen[2002]),

			.SO(gen[2095]),
			.S(gen[2096]),
			.SE(gen[2097]),

			.SELF(gen[2001]),
			.cell_state(gen[2001])
		); 

/******************* CELL 2002 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2002 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1906]),
			.N(gen[1907]),
			.NE(gen[1908]),

			.O(gen[2001]),
			.E(gen[2003]),

			.SO(gen[2096]),
			.S(gen[2097]),
			.SE(gen[2098]),

			.SELF(gen[2002]),
			.cell_state(gen[2002])
		); 

/******************* CELL 2003 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2003 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1907]),
			.N(gen[1908]),
			.NE(gen[1909]),

			.O(gen[2002]),
			.E(gen[2004]),

			.SO(gen[2097]),
			.S(gen[2098]),
			.SE(gen[2099]),

			.SELF(gen[2003]),
			.cell_state(gen[2003])
		); 

/******************* CELL 2004 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2004 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1908]),
			.N(gen[1909]),
			.NE(gen[1910]),

			.O(gen[2003]),
			.E(gen[2005]),

			.SO(gen[2098]),
			.S(gen[2099]),
			.SE(gen[2100]),

			.SELF(gen[2004]),
			.cell_state(gen[2004])
		); 

/******************* CELL 2005 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2005 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1909]),
			.N(gen[1910]),
			.NE(gen[1911]),

			.O(gen[2004]),
			.E(gen[2006]),

			.SO(gen[2099]),
			.S(gen[2100]),
			.SE(gen[2101]),

			.SELF(gen[2005]),
			.cell_state(gen[2005])
		); 

/******************* CELL 2006 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2006 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1910]),
			.N(gen[1911]),
			.NE(gen[1912]),

			.O(gen[2005]),
			.E(gen[2007]),

			.SO(gen[2100]),
			.S(gen[2101]),
			.SE(gen[2102]),

			.SELF(gen[2006]),
			.cell_state(gen[2006])
		); 

/******************* CELL 2007 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2007 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1911]),
			.N(gen[1912]),
			.NE(gen[1913]),

			.O(gen[2006]),
			.E(gen[2008]),

			.SO(gen[2101]),
			.S(gen[2102]),
			.SE(gen[2103]),

			.SELF(gen[2007]),
			.cell_state(gen[2007])
		); 

/******************* CELL 2008 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2008 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1912]),
			.N(gen[1913]),
			.NE(gen[1914]),

			.O(gen[2007]),
			.E(gen[2009]),

			.SO(gen[2102]),
			.S(gen[2103]),
			.SE(gen[2104]),

			.SELF(gen[2008]),
			.cell_state(gen[2008])
		); 

/******************* CELL 2009 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2009 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1913]),
			.N(gen[1914]),
			.NE(gen[1915]),

			.O(gen[2008]),
			.E(gen[2010]),

			.SO(gen[2103]),
			.S(gen[2104]),
			.SE(gen[2105]),

			.SELF(gen[2009]),
			.cell_state(gen[2009])
		); 

/******************* CELL 2010 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2010 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1914]),
			.N(gen[1915]),
			.NE(gen[1916]),

			.O(gen[2009]),
			.E(gen[2011]),

			.SO(gen[2104]),
			.S(gen[2105]),
			.SE(gen[2106]),

			.SELF(gen[2010]),
			.cell_state(gen[2010])
		); 

/******************* CELL 2011 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2011 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1915]),
			.N(gen[1916]),
			.NE(gen[1917]),

			.O(gen[2010]),
			.E(gen[2012]),

			.SO(gen[2105]),
			.S(gen[2106]),
			.SE(gen[2107]),

			.SELF(gen[2011]),
			.cell_state(gen[2011])
		); 

/******************* CELL 2012 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2012 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1916]),
			.N(gen[1917]),
			.NE(gen[1918]),

			.O(gen[2011]),
			.E(gen[2013]),

			.SO(gen[2106]),
			.S(gen[2107]),
			.SE(gen[2108]),

			.SELF(gen[2012]),
			.cell_state(gen[2012])
		); 

/******************* CELL 2013 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2013 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1917]),
			.N(gen[1918]),
			.NE(gen[1919]),

			.O(gen[2012]),
			.E(gen[2014]),

			.SO(gen[2107]),
			.S(gen[2108]),
			.SE(gen[2109]),

			.SELF(gen[2013]),
			.cell_state(gen[2013])
		); 

/******************* CELL 2014 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2014 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1918]),
			.N(gen[1919]),
			.NE(gen[1920]),

			.O(gen[2013]),
			.E(gen[2015]),

			.SO(gen[2108]),
			.S(gen[2109]),
			.SE(gen[2110]),

			.SELF(gen[2014]),
			.cell_state(gen[2014])
		); 

/******************* CELL 2015 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2015 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1919]),
			.N(gen[1920]),
			.NE(gen[1921]),

			.O(gen[2014]),
			.E(gen[2016]),

			.SO(gen[2109]),
			.S(gen[2110]),
			.SE(gen[2111]),

			.SELF(gen[2015]),
			.cell_state(gen[2015])
		); 

/******************* CELL 2016 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2016 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1920]),
			.N(gen[1921]),
			.NE(gen[1922]),

			.O(gen[2015]),
			.E(gen[2017]),

			.SO(gen[2110]),
			.S(gen[2111]),
			.SE(gen[2112]),

			.SELF(gen[2016]),
			.cell_state(gen[2016])
		); 

/******************* CELL 2017 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2017 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1921]),
			.N(gen[1922]),
			.NE(gen[1923]),

			.O(gen[2016]),
			.E(gen[2018]),

			.SO(gen[2111]),
			.S(gen[2112]),
			.SE(gen[2113]),

			.SELF(gen[2017]),
			.cell_state(gen[2017])
		); 

/******************* CELL 2018 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2018 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1922]),
			.N(gen[1923]),
			.NE(gen[1924]),

			.O(gen[2017]),
			.E(gen[2019]),

			.SO(gen[2112]),
			.S(gen[2113]),
			.SE(gen[2114]),

			.SELF(gen[2018]),
			.cell_state(gen[2018])
		); 

/******************* CELL 2019 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2019 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1923]),
			.N(gen[1924]),
			.NE(gen[1925]),

			.O(gen[2018]),
			.E(gen[2020]),

			.SO(gen[2113]),
			.S(gen[2114]),
			.SE(gen[2115]),

			.SELF(gen[2019]),
			.cell_state(gen[2019])
		); 

/******************* CELL 2020 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2020 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1924]),
			.N(gen[1925]),
			.NE(gen[1926]),

			.O(gen[2019]),
			.E(gen[2021]),

			.SO(gen[2114]),
			.S(gen[2115]),
			.SE(gen[2116]),

			.SELF(gen[2020]),
			.cell_state(gen[2020])
		); 

/******************* CELL 2021 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2021 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1925]),
			.N(gen[1926]),
			.NE(gen[1927]),

			.O(gen[2020]),
			.E(gen[2022]),

			.SO(gen[2115]),
			.S(gen[2116]),
			.SE(gen[2117]),

			.SELF(gen[2021]),
			.cell_state(gen[2021])
		); 

/******************* CELL 2022 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2022 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1926]),
			.N(gen[1927]),
			.NE(gen[1928]),

			.O(gen[2021]),
			.E(gen[2023]),

			.SO(gen[2116]),
			.S(gen[2117]),
			.SE(gen[2118]),

			.SELF(gen[2022]),
			.cell_state(gen[2022])
		); 

/******************* CELL 2023 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2023 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1927]),
			.N(gen[1928]),
			.NE(gen[1929]),

			.O(gen[2022]),
			.E(gen[2024]),

			.SO(gen[2117]),
			.S(gen[2118]),
			.SE(gen[2119]),

			.SELF(gen[2023]),
			.cell_state(gen[2023])
		); 

/******************* CELL 2024 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2024 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1928]),
			.N(gen[1929]),
			.NE(gen[1930]),

			.O(gen[2023]),
			.E(gen[2025]),

			.SO(gen[2118]),
			.S(gen[2119]),
			.SE(gen[2120]),

			.SELF(gen[2024]),
			.cell_state(gen[2024])
		); 

/******************* CELL 2025 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2025 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1929]),
			.N(gen[1930]),
			.NE(gen[1931]),

			.O(gen[2024]),
			.E(gen[2026]),

			.SO(gen[2119]),
			.S(gen[2120]),
			.SE(gen[2121]),

			.SELF(gen[2025]),
			.cell_state(gen[2025])
		); 

/******************* CELL 2026 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2026 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1930]),
			.N(gen[1931]),
			.NE(gen[1932]),

			.O(gen[2025]),
			.E(gen[2027]),

			.SO(gen[2120]),
			.S(gen[2121]),
			.SE(gen[2122]),

			.SELF(gen[2026]),
			.cell_state(gen[2026])
		); 

/******************* CELL 2027 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2027 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1931]),
			.N(gen[1932]),
			.NE(gen[1933]),

			.O(gen[2026]),
			.E(gen[2028]),

			.SO(gen[2121]),
			.S(gen[2122]),
			.SE(gen[2123]),

			.SELF(gen[2027]),
			.cell_state(gen[2027])
		); 

/******************* CELL 2028 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2028 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1932]),
			.N(gen[1933]),
			.NE(gen[1934]),

			.O(gen[2027]),
			.E(gen[2029]),

			.SO(gen[2122]),
			.S(gen[2123]),
			.SE(gen[2124]),

			.SELF(gen[2028]),
			.cell_state(gen[2028])
		); 

/******************* CELL 2029 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2029 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1933]),
			.N(gen[1934]),
			.NE(gen[1935]),

			.O(gen[2028]),
			.E(gen[2030]),

			.SO(gen[2123]),
			.S(gen[2124]),
			.SE(gen[2125]),

			.SELF(gen[2029]),
			.cell_state(gen[2029])
		); 

/******************* CELL 2030 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2030 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1934]),
			.N(gen[1935]),
			.NE(gen[1936]),

			.O(gen[2029]),
			.E(gen[2031]),

			.SO(gen[2124]),
			.S(gen[2125]),
			.SE(gen[2126]),

			.SELF(gen[2030]),
			.cell_state(gen[2030])
		); 

/******************* CELL 2031 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2031 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1935]),
			.N(gen[1936]),
			.NE(gen[1937]),

			.O(gen[2030]),
			.E(gen[2032]),

			.SO(gen[2125]),
			.S(gen[2126]),
			.SE(gen[2127]),

			.SELF(gen[2031]),
			.cell_state(gen[2031])
		); 

/******************* CELL 2032 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2032 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1936]),
			.N(gen[1937]),
			.NE(gen[1938]),

			.O(gen[2031]),
			.E(gen[2033]),

			.SO(gen[2126]),
			.S(gen[2127]),
			.SE(gen[2128]),

			.SELF(gen[2032]),
			.cell_state(gen[2032])
		); 

/******************* CELL 2033 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2033 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1937]),
			.N(gen[1938]),
			.NE(gen[1939]),

			.O(gen[2032]),
			.E(gen[2034]),

			.SO(gen[2127]),
			.S(gen[2128]),
			.SE(gen[2129]),

			.SELF(gen[2033]),
			.cell_state(gen[2033])
		); 

/******************* CELL 2034 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2034 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1938]),
			.N(gen[1939]),
			.NE(gen[1940]),

			.O(gen[2033]),
			.E(gen[2035]),

			.SO(gen[2128]),
			.S(gen[2129]),
			.SE(gen[2130]),

			.SELF(gen[2034]),
			.cell_state(gen[2034])
		); 

/******************* CELL 2035 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2035 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1939]),
			.N(gen[1940]),
			.NE(gen[1941]),

			.O(gen[2034]),
			.E(gen[2036]),

			.SO(gen[2129]),
			.S(gen[2130]),
			.SE(gen[2131]),

			.SELF(gen[2035]),
			.cell_state(gen[2035])
		); 

/******************* CELL 2036 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2036 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1940]),
			.N(gen[1941]),
			.NE(gen[1942]),

			.O(gen[2035]),
			.E(gen[2037]),

			.SO(gen[2130]),
			.S(gen[2131]),
			.SE(gen[2132]),

			.SELF(gen[2036]),
			.cell_state(gen[2036])
		); 

/******************* CELL 2037 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2037 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1941]),
			.N(gen[1942]),
			.NE(gen[1943]),

			.O(gen[2036]),
			.E(gen[2038]),

			.SO(gen[2131]),
			.S(gen[2132]),
			.SE(gen[2133]),

			.SELF(gen[2037]),
			.cell_state(gen[2037])
		); 

/******************* CELL 2038 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2038 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1942]),
			.N(gen[1943]),
			.NE(gen[1944]),

			.O(gen[2037]),
			.E(gen[2039]),

			.SO(gen[2132]),
			.S(gen[2133]),
			.SE(gen[2134]),

			.SELF(gen[2038]),
			.cell_state(gen[2038])
		); 

/******************* CELL 2039 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2039 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1943]),
			.N(gen[1944]),
			.NE(gen[1945]),

			.O(gen[2038]),
			.E(gen[2040]),

			.SO(gen[2133]),
			.S(gen[2134]),
			.SE(gen[2135]),

			.SELF(gen[2039]),
			.cell_state(gen[2039])
		); 

/******************* CELL 2040 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2040 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1944]),
			.N(gen[1945]),
			.NE(gen[1946]),

			.O(gen[2039]),
			.E(gen[2041]),

			.SO(gen[2134]),
			.S(gen[2135]),
			.SE(gen[2136]),

			.SELF(gen[2040]),
			.cell_state(gen[2040])
		); 

/******************* CELL 2041 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2041 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1945]),
			.N(gen[1946]),
			.NE(gen[1947]),

			.O(gen[2040]),
			.E(gen[2042]),

			.SO(gen[2135]),
			.S(gen[2136]),
			.SE(gen[2137]),

			.SELF(gen[2041]),
			.cell_state(gen[2041])
		); 

/******************* CELL 2042 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2042 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1946]),
			.N(gen[1947]),
			.NE(gen[1948]),

			.O(gen[2041]),
			.E(gen[2043]),

			.SO(gen[2136]),
			.S(gen[2137]),
			.SE(gen[2138]),

			.SELF(gen[2042]),
			.cell_state(gen[2042])
		); 

/******************* CELL 2043 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2043 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1947]),
			.N(gen[1948]),
			.NE(gen[1949]),

			.O(gen[2042]),
			.E(gen[2044]),

			.SO(gen[2137]),
			.S(gen[2138]),
			.SE(gen[2139]),

			.SELF(gen[2043]),
			.cell_state(gen[2043])
		); 

/******************* CELL 2044 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2044 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1948]),
			.N(gen[1949]),
			.NE(gen[1950]),

			.O(gen[2043]),
			.E(gen[2045]),

			.SO(gen[2138]),
			.S(gen[2139]),
			.SE(gen[2140]),

			.SELF(gen[2044]),
			.cell_state(gen[2044])
		); 

/******************* CELL 2045 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2045 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1949]),
			.N(gen[1950]),
			.NE(gen[1951]),

			.O(gen[2044]),
			.E(gen[2046]),

			.SO(gen[2139]),
			.S(gen[2140]),
			.SE(gen[2141]),

			.SELF(gen[2045]),
			.cell_state(gen[2045])
		); 

/******************* CELL 2046 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2046 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1950]),
			.N(gen[1951]),
			.NE(gen[1952]),

			.O(gen[2045]),
			.E(gen[2047]),

			.SO(gen[2140]),
			.S(gen[2141]),
			.SE(gen[2142]),

			.SELF(gen[2046]),
			.cell_state(gen[2046])
		); 

/******************* CELL 2047 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2047 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1951]),
			.N(gen[1952]),
			.NE(gen[1953]),

			.O(gen[2046]),
			.E(gen[2048]),

			.SO(gen[2141]),
			.S(gen[2142]),
			.SE(gen[2143]),

			.SELF(gen[2047]),
			.cell_state(gen[2047])
		); 

/******************* CELL 2048 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2048 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1952]),
			.N(gen[1953]),
			.NE(gen[1954]),

			.O(gen[2047]),
			.E(gen[2049]),

			.SO(gen[2142]),
			.S(gen[2143]),
			.SE(gen[2144]),

			.SELF(gen[2048]),
			.cell_state(gen[2048])
		); 

/******************* CELL 2049 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2049 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1953]),
			.N(gen[1954]),
			.NE(gen[1955]),

			.O(gen[2048]),
			.E(gen[2050]),

			.SO(gen[2143]),
			.S(gen[2144]),
			.SE(gen[2145]),

			.SELF(gen[2049]),
			.cell_state(gen[2049])
		); 

/******************* CELL 2050 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2050 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1954]),
			.N(gen[1955]),
			.NE(gen[1956]),

			.O(gen[2049]),
			.E(gen[2051]),

			.SO(gen[2144]),
			.S(gen[2145]),
			.SE(gen[2146]),

			.SELF(gen[2050]),
			.cell_state(gen[2050])
		); 

/******************* CELL 2051 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2051 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1955]),
			.N(gen[1956]),
			.NE(gen[1957]),

			.O(gen[2050]),
			.E(gen[2052]),

			.SO(gen[2145]),
			.S(gen[2146]),
			.SE(gen[2147]),

			.SELF(gen[2051]),
			.cell_state(gen[2051])
		); 

/******************* CELL 2052 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2052 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1956]),
			.N(gen[1957]),
			.NE(gen[1958]),

			.O(gen[2051]),
			.E(gen[2053]),

			.SO(gen[2146]),
			.S(gen[2147]),
			.SE(gen[2148]),

			.SELF(gen[2052]),
			.cell_state(gen[2052])
		); 

/******************* CELL 2053 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2053 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1957]),
			.N(gen[1958]),
			.NE(gen[1959]),

			.O(gen[2052]),
			.E(gen[2054]),

			.SO(gen[2147]),
			.S(gen[2148]),
			.SE(gen[2149]),

			.SELF(gen[2053]),
			.cell_state(gen[2053])
		); 

/******************* CELL 2054 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2054 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1958]),
			.N(gen[1959]),
			.NE(gen[1960]),

			.O(gen[2053]),
			.E(gen[2055]),

			.SO(gen[2148]),
			.S(gen[2149]),
			.SE(gen[2150]),

			.SELF(gen[2054]),
			.cell_state(gen[2054])
		); 

/******************* CELL 2055 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2055 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1959]),
			.N(gen[1960]),
			.NE(gen[1961]),

			.O(gen[2054]),
			.E(gen[2056]),

			.SO(gen[2149]),
			.S(gen[2150]),
			.SE(gen[2151]),

			.SELF(gen[2055]),
			.cell_state(gen[2055])
		); 

/******************* CELL 2056 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2056 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1960]),
			.N(gen[1961]),
			.NE(gen[1962]),

			.O(gen[2055]),
			.E(gen[2057]),

			.SO(gen[2150]),
			.S(gen[2151]),
			.SE(gen[2152]),

			.SELF(gen[2056]),
			.cell_state(gen[2056])
		); 

/******************* CELL 2057 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2057 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1961]),
			.N(gen[1962]),
			.NE(gen[1963]),

			.O(gen[2056]),
			.E(gen[2058]),

			.SO(gen[2151]),
			.S(gen[2152]),
			.SE(gen[2153]),

			.SELF(gen[2057]),
			.cell_state(gen[2057])
		); 

/******************* CELL 2058 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2058 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1962]),
			.N(gen[1963]),
			.NE(gen[1964]),

			.O(gen[2057]),
			.E(gen[2059]),

			.SO(gen[2152]),
			.S(gen[2153]),
			.SE(gen[2154]),

			.SELF(gen[2058]),
			.cell_state(gen[2058])
		); 

/******************* CELL 2059 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2059 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1963]),
			.N(gen[1964]),
			.NE(gen[1965]),

			.O(gen[2058]),
			.E(gen[2060]),

			.SO(gen[2153]),
			.S(gen[2154]),
			.SE(gen[2155]),

			.SELF(gen[2059]),
			.cell_state(gen[2059])
		); 

/******************* CELL 2060 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2060 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1964]),
			.N(gen[1965]),
			.NE(gen[1966]),

			.O(gen[2059]),
			.E(gen[2061]),

			.SO(gen[2154]),
			.S(gen[2155]),
			.SE(gen[2156]),

			.SELF(gen[2060]),
			.cell_state(gen[2060])
		); 

/******************* CELL 2061 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2061 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1965]),
			.N(gen[1966]),
			.NE(gen[1967]),

			.O(gen[2060]),
			.E(gen[2062]),

			.SO(gen[2155]),
			.S(gen[2156]),
			.SE(gen[2157]),

			.SELF(gen[2061]),
			.cell_state(gen[2061])
		); 

/******************* CELL 2062 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2062 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1966]),
			.N(gen[1967]),
			.NE(gen[1968]),

			.O(gen[2061]),
			.E(gen[2063]),

			.SO(gen[2156]),
			.S(gen[2157]),
			.SE(gen[2158]),

			.SELF(gen[2062]),
			.cell_state(gen[2062])
		); 

/******************* CELL 2063 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2063 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1967]),
			.N(gen[1968]),
			.NE(gen[1969]),

			.O(gen[2062]),
			.E(gen[2064]),

			.SO(gen[2157]),
			.S(gen[2158]),
			.SE(gen[2159]),

			.SELF(gen[2063]),
			.cell_state(gen[2063])
		); 

/******************* CELL 2064 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2064 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1968]),
			.N(gen[1969]),
			.NE(gen[1970]),

			.O(gen[2063]),
			.E(gen[2065]),

			.SO(gen[2158]),
			.S(gen[2159]),
			.SE(gen[2160]),

			.SELF(gen[2064]),
			.cell_state(gen[2064])
		); 

/******************* CELL 2065 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2065 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1969]),
			.N(gen[1970]),
			.NE(gen[1971]),

			.O(gen[2064]),
			.E(gen[2066]),

			.SO(gen[2159]),
			.S(gen[2160]),
			.SE(gen[2161]),

			.SELF(gen[2065]),
			.cell_state(gen[2065])
		); 

/******************* CELL 2066 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2066 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1970]),
			.N(gen[1971]),
			.NE(gen[1972]),

			.O(gen[2065]),
			.E(gen[2067]),

			.SO(gen[2160]),
			.S(gen[2161]),
			.SE(gen[2162]),

			.SELF(gen[2066]),
			.cell_state(gen[2066])
		); 

/******************* CELL 2067 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2067 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1971]),
			.N(gen[1972]),
			.NE(gen[1973]),

			.O(gen[2066]),
			.E(gen[2068]),

			.SO(gen[2161]),
			.S(gen[2162]),
			.SE(gen[2163]),

			.SELF(gen[2067]),
			.cell_state(gen[2067])
		); 

/******************* CELL 2068 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2068 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1972]),
			.N(gen[1973]),
			.NE(gen[1974]),

			.O(gen[2067]),
			.E(gen[2069]),

			.SO(gen[2162]),
			.S(gen[2163]),
			.SE(gen[2164]),

			.SELF(gen[2068]),
			.cell_state(gen[2068])
		); 

/******************* CELL 2069 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2069 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1973]),
			.N(gen[1974]),
			.NE(gen[1975]),

			.O(gen[2068]),
			.E(gen[2070]),

			.SO(gen[2163]),
			.S(gen[2164]),
			.SE(gen[2165]),

			.SELF(gen[2069]),
			.cell_state(gen[2069])
		); 

/******************* CELL 2070 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2070 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1974]),
			.N(gen[1975]),
			.NE(gen[1976]),

			.O(gen[2069]),
			.E(gen[2071]),

			.SO(gen[2164]),
			.S(gen[2165]),
			.SE(gen[2166]),

			.SELF(gen[2070]),
			.cell_state(gen[2070])
		); 

/******************* CELL 2071 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2071 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1975]),
			.N(gen[1976]),
			.NE(gen[1977]),

			.O(gen[2070]),
			.E(gen[2072]),

			.SO(gen[2165]),
			.S(gen[2166]),
			.SE(gen[2167]),

			.SELF(gen[2071]),
			.cell_state(gen[2071])
		); 

/******************* CELL 2072 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2072 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1976]),
			.N(gen[1977]),
			.NE(gen[1978]),

			.O(gen[2071]),
			.E(gen[2073]),

			.SO(gen[2166]),
			.S(gen[2167]),
			.SE(gen[2168]),

			.SELF(gen[2072]),
			.cell_state(gen[2072])
		); 

/******************* CELL 2073 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2073 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1977]),
			.N(gen[1978]),
			.NE(gen[1979]),

			.O(gen[2072]),
			.E(gen[2074]),

			.SO(gen[2167]),
			.S(gen[2168]),
			.SE(gen[2169]),

			.SELF(gen[2073]),
			.cell_state(gen[2073])
		); 

/******************* CELL 2074 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2074 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1978]),
			.N(gen[1979]),
			.NE(gen[1980]),

			.O(gen[2073]),
			.E(gen[2075]),

			.SO(gen[2168]),
			.S(gen[2169]),
			.SE(gen[2170]),

			.SELF(gen[2074]),
			.cell_state(gen[2074])
		); 

/******************* CELL 2075 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2075 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1979]),
			.N(gen[1980]),
			.NE(gen[1981]),

			.O(gen[2074]),
			.E(gen[2076]),

			.SO(gen[2169]),
			.S(gen[2170]),
			.SE(gen[2171]),

			.SELF(gen[2075]),
			.cell_state(gen[2075])
		); 

/******************* CELL 2076 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2076 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1980]),
			.N(gen[1981]),
			.NE(gen[1982]),

			.O(gen[2075]),
			.E(gen[2077]),

			.SO(gen[2170]),
			.S(gen[2171]),
			.SE(gen[2172]),

			.SELF(gen[2076]),
			.cell_state(gen[2076])
		); 

/******************* CELL 2077 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2077 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1981]),
			.N(gen[1982]),
			.NE(gen[1983]),

			.O(gen[2076]),
			.E(gen[2078]),

			.SO(gen[2171]),
			.S(gen[2172]),
			.SE(gen[2173]),

			.SELF(gen[2077]),
			.cell_state(gen[2077])
		); 

/******************* CELL 2078 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2078 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1982]),
			.N(gen[1983]),
			.NE(gen[1984]),

			.O(gen[2077]),
			.E(gen[2079]),

			.SO(gen[2172]),
			.S(gen[2173]),
			.SE(gen[2174]),

			.SELF(gen[2078]),
			.cell_state(gen[2078])
		); 

/******************* CELL 2079 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2079 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1983]),
			.N(gen[1984]),
			.NE(gen[1985]),

			.O(gen[2078]),
			.E(gen[2080]),

			.SO(gen[2173]),
			.S(gen[2174]),
			.SE(gen[2175]),

			.SELF(gen[2079]),
			.cell_state(gen[2079])
		); 

/******************* CELL 2080 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2080 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1984]),
			.N(gen[1985]),
			.NE(gen[1986]),

			.O(gen[2079]),
			.E(gen[2081]),

			.SO(gen[2174]),
			.S(gen[2175]),
			.SE(gen[2176]),

			.SELF(gen[2080]),
			.cell_state(gen[2080])
		); 

/******************* CELL 2081 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2081 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1985]),
			.N(gen[1986]),
			.NE(gen[1987]),

			.O(gen[2080]),
			.E(gen[2082]),

			.SO(gen[2175]),
			.S(gen[2176]),
			.SE(gen[2177]),

			.SELF(gen[2081]),
			.cell_state(gen[2081])
		); 

/******************* CELL 2082 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2082 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1986]),
			.N(gen[1987]),
			.NE(gen[1988]),

			.O(gen[2081]),
			.E(gen[2083]),

			.SO(gen[2176]),
			.S(gen[2177]),
			.SE(gen[2178]),

			.SELF(gen[2082]),
			.cell_state(gen[2082])
		); 

/******************* CELL 2083 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2083 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1987]),
			.N(gen[1988]),
			.NE(gen[1989]),

			.O(gen[2082]),
			.E(gen[2084]),

			.SO(gen[2177]),
			.S(gen[2178]),
			.SE(gen[2179]),

			.SELF(gen[2083]),
			.cell_state(gen[2083])
		); 

/******************* CELL 2084 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2084 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1988]),
			.N(gen[1989]),
			.NE(gen[1990]),

			.O(gen[2083]),
			.E(gen[2085]),

			.SO(gen[2178]),
			.S(gen[2179]),
			.SE(gen[2180]),

			.SELF(gen[2084]),
			.cell_state(gen[2084])
		); 

/******************* CELL 2085 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2085 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1989]),
			.N(gen[1990]),
			.NE(gen[1991]),

			.O(gen[2084]),
			.E(gen[2086]),

			.SO(gen[2179]),
			.S(gen[2180]),
			.SE(gen[2181]),

			.SELF(gen[2085]),
			.cell_state(gen[2085])
		); 

/******************* CELL 2086 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2086 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1990]),
			.N(gen[1991]),
			.NE(gen[1992]),

			.O(gen[2085]),
			.E(gen[2087]),

			.SO(gen[2180]),
			.S(gen[2181]),
			.SE(gen[2182]),

			.SELF(gen[2086]),
			.cell_state(gen[2086])
		); 

/******************* CELL 2087 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2087 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1991]),
			.N(gen[1992]),
			.NE(gen[1993]),

			.O(gen[2086]),
			.E(gen[2088]),

			.SO(gen[2181]),
			.S(gen[2182]),
			.SE(gen[2183]),

			.SELF(gen[2087]),
			.cell_state(gen[2087])
		); 

/******************* CELL 2088 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2088 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1992]),
			.N(gen[1993]),
			.NE(gen[1994]),

			.O(gen[2087]),
			.E(gen[2089]),

			.SO(gen[2182]),
			.S(gen[2183]),
			.SE(gen[2184]),

			.SELF(gen[2088]),
			.cell_state(gen[2088])
		); 

/******************* CELL 2089 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2089 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1993]),
			.N(gen[1994]),
			.NE(gen[1993]),

			.O(gen[2088]),
			.E(gen[2088]),

			.SO(gen[2183]),
			.S(gen[2184]),
			.SE(gen[2183]),

			.SELF(gen[2089]),
			.cell_state(gen[2089])
		); 

/******************* CELL 2090 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2090 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1996]),
			.N(gen[1995]),
			.NE(gen[1996]),

			.O(gen[2091]),
			.E(gen[2091]),

			.SO(gen[2186]),
			.S(gen[2185]),
			.SE(gen[2186]),

			.SELF(gen[2090]),
			.cell_state(gen[2090])
		); 

/******************* CELL 2091 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2091 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1995]),
			.N(gen[1996]),
			.NE(gen[1997]),

			.O(gen[2090]),
			.E(gen[2092]),

			.SO(gen[2185]),
			.S(gen[2186]),
			.SE(gen[2187]),

			.SELF(gen[2091]),
			.cell_state(gen[2091])
		); 

/******************* CELL 2092 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2092 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1996]),
			.N(gen[1997]),
			.NE(gen[1998]),

			.O(gen[2091]),
			.E(gen[2093]),

			.SO(gen[2186]),
			.S(gen[2187]),
			.SE(gen[2188]),

			.SELF(gen[2092]),
			.cell_state(gen[2092])
		); 

/******************* CELL 2093 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2093 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1997]),
			.N(gen[1998]),
			.NE(gen[1999]),

			.O(gen[2092]),
			.E(gen[2094]),

			.SO(gen[2187]),
			.S(gen[2188]),
			.SE(gen[2189]),

			.SELF(gen[2093]),
			.cell_state(gen[2093])
		); 

/******************* CELL 2094 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2094 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1998]),
			.N(gen[1999]),
			.NE(gen[2000]),

			.O(gen[2093]),
			.E(gen[2095]),

			.SO(gen[2188]),
			.S(gen[2189]),
			.SE(gen[2190]),

			.SELF(gen[2094]),
			.cell_state(gen[2094])
		); 

/******************* CELL 2095 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2095 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1999]),
			.N(gen[2000]),
			.NE(gen[2001]),

			.O(gen[2094]),
			.E(gen[2096]),

			.SO(gen[2189]),
			.S(gen[2190]),
			.SE(gen[2191]),

			.SELF(gen[2095]),
			.cell_state(gen[2095])
		); 

/******************* CELL 2096 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2096 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2000]),
			.N(gen[2001]),
			.NE(gen[2002]),

			.O(gen[2095]),
			.E(gen[2097]),

			.SO(gen[2190]),
			.S(gen[2191]),
			.SE(gen[2192]),

			.SELF(gen[2096]),
			.cell_state(gen[2096])
		); 

/******************* CELL 2097 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2097 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2001]),
			.N(gen[2002]),
			.NE(gen[2003]),

			.O(gen[2096]),
			.E(gen[2098]),

			.SO(gen[2191]),
			.S(gen[2192]),
			.SE(gen[2193]),

			.SELF(gen[2097]),
			.cell_state(gen[2097])
		); 

/******************* CELL 2098 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2098 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2002]),
			.N(gen[2003]),
			.NE(gen[2004]),

			.O(gen[2097]),
			.E(gen[2099]),

			.SO(gen[2192]),
			.S(gen[2193]),
			.SE(gen[2194]),

			.SELF(gen[2098]),
			.cell_state(gen[2098])
		); 

/******************* CELL 2099 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2099 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2003]),
			.N(gen[2004]),
			.NE(gen[2005]),

			.O(gen[2098]),
			.E(gen[2100]),

			.SO(gen[2193]),
			.S(gen[2194]),
			.SE(gen[2195]),

			.SELF(gen[2099]),
			.cell_state(gen[2099])
		); 

/******************* CELL 2100 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2100 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2004]),
			.N(gen[2005]),
			.NE(gen[2006]),

			.O(gen[2099]),
			.E(gen[2101]),

			.SO(gen[2194]),
			.S(gen[2195]),
			.SE(gen[2196]),

			.SELF(gen[2100]),
			.cell_state(gen[2100])
		); 

/******************* CELL 2101 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2101 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2005]),
			.N(gen[2006]),
			.NE(gen[2007]),

			.O(gen[2100]),
			.E(gen[2102]),

			.SO(gen[2195]),
			.S(gen[2196]),
			.SE(gen[2197]),

			.SELF(gen[2101]),
			.cell_state(gen[2101])
		); 

/******************* CELL 2102 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2102 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2006]),
			.N(gen[2007]),
			.NE(gen[2008]),

			.O(gen[2101]),
			.E(gen[2103]),

			.SO(gen[2196]),
			.S(gen[2197]),
			.SE(gen[2198]),

			.SELF(gen[2102]),
			.cell_state(gen[2102])
		); 

/******************* CELL 2103 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2103 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2007]),
			.N(gen[2008]),
			.NE(gen[2009]),

			.O(gen[2102]),
			.E(gen[2104]),

			.SO(gen[2197]),
			.S(gen[2198]),
			.SE(gen[2199]),

			.SELF(gen[2103]),
			.cell_state(gen[2103])
		); 

/******************* CELL 2104 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2104 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2008]),
			.N(gen[2009]),
			.NE(gen[2010]),

			.O(gen[2103]),
			.E(gen[2105]),

			.SO(gen[2198]),
			.S(gen[2199]),
			.SE(gen[2200]),

			.SELF(gen[2104]),
			.cell_state(gen[2104])
		); 

/******************* CELL 2105 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2105 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2009]),
			.N(gen[2010]),
			.NE(gen[2011]),

			.O(gen[2104]),
			.E(gen[2106]),

			.SO(gen[2199]),
			.S(gen[2200]),
			.SE(gen[2201]),

			.SELF(gen[2105]),
			.cell_state(gen[2105])
		); 

/******************* CELL 2106 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2106 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2010]),
			.N(gen[2011]),
			.NE(gen[2012]),

			.O(gen[2105]),
			.E(gen[2107]),

			.SO(gen[2200]),
			.S(gen[2201]),
			.SE(gen[2202]),

			.SELF(gen[2106]),
			.cell_state(gen[2106])
		); 

/******************* CELL 2107 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2107 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2011]),
			.N(gen[2012]),
			.NE(gen[2013]),

			.O(gen[2106]),
			.E(gen[2108]),

			.SO(gen[2201]),
			.S(gen[2202]),
			.SE(gen[2203]),

			.SELF(gen[2107]),
			.cell_state(gen[2107])
		); 

/******************* CELL 2108 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2108 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2012]),
			.N(gen[2013]),
			.NE(gen[2014]),

			.O(gen[2107]),
			.E(gen[2109]),

			.SO(gen[2202]),
			.S(gen[2203]),
			.SE(gen[2204]),

			.SELF(gen[2108]),
			.cell_state(gen[2108])
		); 

/******************* CELL 2109 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2109 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2013]),
			.N(gen[2014]),
			.NE(gen[2015]),

			.O(gen[2108]),
			.E(gen[2110]),

			.SO(gen[2203]),
			.S(gen[2204]),
			.SE(gen[2205]),

			.SELF(gen[2109]),
			.cell_state(gen[2109])
		); 

/******************* CELL 2110 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2110 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2014]),
			.N(gen[2015]),
			.NE(gen[2016]),

			.O(gen[2109]),
			.E(gen[2111]),

			.SO(gen[2204]),
			.S(gen[2205]),
			.SE(gen[2206]),

			.SELF(gen[2110]),
			.cell_state(gen[2110])
		); 

/******************* CELL 2111 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2111 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2015]),
			.N(gen[2016]),
			.NE(gen[2017]),

			.O(gen[2110]),
			.E(gen[2112]),

			.SO(gen[2205]),
			.S(gen[2206]),
			.SE(gen[2207]),

			.SELF(gen[2111]),
			.cell_state(gen[2111])
		); 

/******************* CELL 2112 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2112 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2016]),
			.N(gen[2017]),
			.NE(gen[2018]),

			.O(gen[2111]),
			.E(gen[2113]),

			.SO(gen[2206]),
			.S(gen[2207]),
			.SE(gen[2208]),

			.SELF(gen[2112]),
			.cell_state(gen[2112])
		); 

/******************* CELL 2113 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2113 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2017]),
			.N(gen[2018]),
			.NE(gen[2019]),

			.O(gen[2112]),
			.E(gen[2114]),

			.SO(gen[2207]),
			.S(gen[2208]),
			.SE(gen[2209]),

			.SELF(gen[2113]),
			.cell_state(gen[2113])
		); 

/******************* CELL 2114 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2114 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2018]),
			.N(gen[2019]),
			.NE(gen[2020]),

			.O(gen[2113]),
			.E(gen[2115]),

			.SO(gen[2208]),
			.S(gen[2209]),
			.SE(gen[2210]),

			.SELF(gen[2114]),
			.cell_state(gen[2114])
		); 

/******************* CELL 2115 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2115 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2019]),
			.N(gen[2020]),
			.NE(gen[2021]),

			.O(gen[2114]),
			.E(gen[2116]),

			.SO(gen[2209]),
			.S(gen[2210]),
			.SE(gen[2211]),

			.SELF(gen[2115]),
			.cell_state(gen[2115])
		); 

/******************* CELL 2116 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2116 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2020]),
			.N(gen[2021]),
			.NE(gen[2022]),

			.O(gen[2115]),
			.E(gen[2117]),

			.SO(gen[2210]),
			.S(gen[2211]),
			.SE(gen[2212]),

			.SELF(gen[2116]),
			.cell_state(gen[2116])
		); 

/******************* CELL 2117 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2117 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2021]),
			.N(gen[2022]),
			.NE(gen[2023]),

			.O(gen[2116]),
			.E(gen[2118]),

			.SO(gen[2211]),
			.S(gen[2212]),
			.SE(gen[2213]),

			.SELF(gen[2117]),
			.cell_state(gen[2117])
		); 

/******************* CELL 2118 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2118 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2022]),
			.N(gen[2023]),
			.NE(gen[2024]),

			.O(gen[2117]),
			.E(gen[2119]),

			.SO(gen[2212]),
			.S(gen[2213]),
			.SE(gen[2214]),

			.SELF(gen[2118]),
			.cell_state(gen[2118])
		); 

/******************* CELL 2119 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2119 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2023]),
			.N(gen[2024]),
			.NE(gen[2025]),

			.O(gen[2118]),
			.E(gen[2120]),

			.SO(gen[2213]),
			.S(gen[2214]),
			.SE(gen[2215]),

			.SELF(gen[2119]),
			.cell_state(gen[2119])
		); 

/******************* CELL 2120 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2120 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2024]),
			.N(gen[2025]),
			.NE(gen[2026]),

			.O(gen[2119]),
			.E(gen[2121]),

			.SO(gen[2214]),
			.S(gen[2215]),
			.SE(gen[2216]),

			.SELF(gen[2120]),
			.cell_state(gen[2120])
		); 

/******************* CELL 2121 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2121 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2025]),
			.N(gen[2026]),
			.NE(gen[2027]),

			.O(gen[2120]),
			.E(gen[2122]),

			.SO(gen[2215]),
			.S(gen[2216]),
			.SE(gen[2217]),

			.SELF(gen[2121]),
			.cell_state(gen[2121])
		); 

/******************* CELL 2122 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2122 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2026]),
			.N(gen[2027]),
			.NE(gen[2028]),

			.O(gen[2121]),
			.E(gen[2123]),

			.SO(gen[2216]),
			.S(gen[2217]),
			.SE(gen[2218]),

			.SELF(gen[2122]),
			.cell_state(gen[2122])
		); 

/******************* CELL 2123 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2123 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2027]),
			.N(gen[2028]),
			.NE(gen[2029]),

			.O(gen[2122]),
			.E(gen[2124]),

			.SO(gen[2217]),
			.S(gen[2218]),
			.SE(gen[2219]),

			.SELF(gen[2123]),
			.cell_state(gen[2123])
		); 

/******************* CELL 2124 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2124 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2028]),
			.N(gen[2029]),
			.NE(gen[2030]),

			.O(gen[2123]),
			.E(gen[2125]),

			.SO(gen[2218]),
			.S(gen[2219]),
			.SE(gen[2220]),

			.SELF(gen[2124]),
			.cell_state(gen[2124])
		); 

/******************* CELL 2125 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2125 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2029]),
			.N(gen[2030]),
			.NE(gen[2031]),

			.O(gen[2124]),
			.E(gen[2126]),

			.SO(gen[2219]),
			.S(gen[2220]),
			.SE(gen[2221]),

			.SELF(gen[2125]),
			.cell_state(gen[2125])
		); 

/******************* CELL 2126 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2126 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2030]),
			.N(gen[2031]),
			.NE(gen[2032]),

			.O(gen[2125]),
			.E(gen[2127]),

			.SO(gen[2220]),
			.S(gen[2221]),
			.SE(gen[2222]),

			.SELF(gen[2126]),
			.cell_state(gen[2126])
		); 

/******************* CELL 2127 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2127 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2031]),
			.N(gen[2032]),
			.NE(gen[2033]),

			.O(gen[2126]),
			.E(gen[2128]),

			.SO(gen[2221]),
			.S(gen[2222]),
			.SE(gen[2223]),

			.SELF(gen[2127]),
			.cell_state(gen[2127])
		); 

/******************* CELL 2128 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2128 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2032]),
			.N(gen[2033]),
			.NE(gen[2034]),

			.O(gen[2127]),
			.E(gen[2129]),

			.SO(gen[2222]),
			.S(gen[2223]),
			.SE(gen[2224]),

			.SELF(gen[2128]),
			.cell_state(gen[2128])
		); 

/******************* CELL 2129 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2129 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2033]),
			.N(gen[2034]),
			.NE(gen[2035]),

			.O(gen[2128]),
			.E(gen[2130]),

			.SO(gen[2223]),
			.S(gen[2224]),
			.SE(gen[2225]),

			.SELF(gen[2129]),
			.cell_state(gen[2129])
		); 

/******************* CELL 2130 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2130 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2034]),
			.N(gen[2035]),
			.NE(gen[2036]),

			.O(gen[2129]),
			.E(gen[2131]),

			.SO(gen[2224]),
			.S(gen[2225]),
			.SE(gen[2226]),

			.SELF(gen[2130]),
			.cell_state(gen[2130])
		); 

/******************* CELL 2131 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2131 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2035]),
			.N(gen[2036]),
			.NE(gen[2037]),

			.O(gen[2130]),
			.E(gen[2132]),

			.SO(gen[2225]),
			.S(gen[2226]),
			.SE(gen[2227]),

			.SELF(gen[2131]),
			.cell_state(gen[2131])
		); 

/******************* CELL 2132 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2132 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2036]),
			.N(gen[2037]),
			.NE(gen[2038]),

			.O(gen[2131]),
			.E(gen[2133]),

			.SO(gen[2226]),
			.S(gen[2227]),
			.SE(gen[2228]),

			.SELF(gen[2132]),
			.cell_state(gen[2132])
		); 

/******************* CELL 2133 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2133 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2037]),
			.N(gen[2038]),
			.NE(gen[2039]),

			.O(gen[2132]),
			.E(gen[2134]),

			.SO(gen[2227]),
			.S(gen[2228]),
			.SE(gen[2229]),

			.SELF(gen[2133]),
			.cell_state(gen[2133])
		); 

/******************* CELL 2134 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2134 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2038]),
			.N(gen[2039]),
			.NE(gen[2040]),

			.O(gen[2133]),
			.E(gen[2135]),

			.SO(gen[2228]),
			.S(gen[2229]),
			.SE(gen[2230]),

			.SELF(gen[2134]),
			.cell_state(gen[2134])
		); 

/******************* CELL 2135 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2135 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2039]),
			.N(gen[2040]),
			.NE(gen[2041]),

			.O(gen[2134]),
			.E(gen[2136]),

			.SO(gen[2229]),
			.S(gen[2230]),
			.SE(gen[2231]),

			.SELF(gen[2135]),
			.cell_state(gen[2135])
		); 

/******************* CELL 2136 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2136 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2040]),
			.N(gen[2041]),
			.NE(gen[2042]),

			.O(gen[2135]),
			.E(gen[2137]),

			.SO(gen[2230]),
			.S(gen[2231]),
			.SE(gen[2232]),

			.SELF(gen[2136]),
			.cell_state(gen[2136])
		); 

/******************* CELL 2137 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2137 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2041]),
			.N(gen[2042]),
			.NE(gen[2043]),

			.O(gen[2136]),
			.E(gen[2138]),

			.SO(gen[2231]),
			.S(gen[2232]),
			.SE(gen[2233]),

			.SELF(gen[2137]),
			.cell_state(gen[2137])
		); 

/******************* CELL 2138 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2138 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2042]),
			.N(gen[2043]),
			.NE(gen[2044]),

			.O(gen[2137]),
			.E(gen[2139]),

			.SO(gen[2232]),
			.S(gen[2233]),
			.SE(gen[2234]),

			.SELF(gen[2138]),
			.cell_state(gen[2138])
		); 

/******************* CELL 2139 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2139 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2043]),
			.N(gen[2044]),
			.NE(gen[2045]),

			.O(gen[2138]),
			.E(gen[2140]),

			.SO(gen[2233]),
			.S(gen[2234]),
			.SE(gen[2235]),

			.SELF(gen[2139]),
			.cell_state(gen[2139])
		); 

/******************* CELL 2140 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2140 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2044]),
			.N(gen[2045]),
			.NE(gen[2046]),

			.O(gen[2139]),
			.E(gen[2141]),

			.SO(gen[2234]),
			.S(gen[2235]),
			.SE(gen[2236]),

			.SELF(gen[2140]),
			.cell_state(gen[2140])
		); 

/******************* CELL 2141 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2141 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2045]),
			.N(gen[2046]),
			.NE(gen[2047]),

			.O(gen[2140]),
			.E(gen[2142]),

			.SO(gen[2235]),
			.S(gen[2236]),
			.SE(gen[2237]),

			.SELF(gen[2141]),
			.cell_state(gen[2141])
		); 

/******************* CELL 2142 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2142 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2046]),
			.N(gen[2047]),
			.NE(gen[2048]),

			.O(gen[2141]),
			.E(gen[2143]),

			.SO(gen[2236]),
			.S(gen[2237]),
			.SE(gen[2238]),

			.SELF(gen[2142]),
			.cell_state(gen[2142])
		); 

/******************* CELL 2143 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2143 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2047]),
			.N(gen[2048]),
			.NE(gen[2049]),

			.O(gen[2142]),
			.E(gen[2144]),

			.SO(gen[2237]),
			.S(gen[2238]),
			.SE(gen[2239]),

			.SELF(gen[2143]),
			.cell_state(gen[2143])
		); 

/******************* CELL 2144 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2144 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2048]),
			.N(gen[2049]),
			.NE(gen[2050]),

			.O(gen[2143]),
			.E(gen[2145]),

			.SO(gen[2238]),
			.S(gen[2239]),
			.SE(gen[2240]),

			.SELF(gen[2144]),
			.cell_state(gen[2144])
		); 

/******************* CELL 2145 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2145 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2049]),
			.N(gen[2050]),
			.NE(gen[2051]),

			.O(gen[2144]),
			.E(gen[2146]),

			.SO(gen[2239]),
			.S(gen[2240]),
			.SE(gen[2241]),

			.SELF(gen[2145]),
			.cell_state(gen[2145])
		); 

/******************* CELL 2146 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2146 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2050]),
			.N(gen[2051]),
			.NE(gen[2052]),

			.O(gen[2145]),
			.E(gen[2147]),

			.SO(gen[2240]),
			.S(gen[2241]),
			.SE(gen[2242]),

			.SELF(gen[2146]),
			.cell_state(gen[2146])
		); 

/******************* CELL 2147 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2147 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2051]),
			.N(gen[2052]),
			.NE(gen[2053]),

			.O(gen[2146]),
			.E(gen[2148]),

			.SO(gen[2241]),
			.S(gen[2242]),
			.SE(gen[2243]),

			.SELF(gen[2147]),
			.cell_state(gen[2147])
		); 

/******************* CELL 2148 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2148 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2052]),
			.N(gen[2053]),
			.NE(gen[2054]),

			.O(gen[2147]),
			.E(gen[2149]),

			.SO(gen[2242]),
			.S(gen[2243]),
			.SE(gen[2244]),

			.SELF(gen[2148]),
			.cell_state(gen[2148])
		); 

/******************* CELL 2149 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2149 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2053]),
			.N(gen[2054]),
			.NE(gen[2055]),

			.O(gen[2148]),
			.E(gen[2150]),

			.SO(gen[2243]),
			.S(gen[2244]),
			.SE(gen[2245]),

			.SELF(gen[2149]),
			.cell_state(gen[2149])
		); 

/******************* CELL 2150 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2150 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2054]),
			.N(gen[2055]),
			.NE(gen[2056]),

			.O(gen[2149]),
			.E(gen[2151]),

			.SO(gen[2244]),
			.S(gen[2245]),
			.SE(gen[2246]),

			.SELF(gen[2150]),
			.cell_state(gen[2150])
		); 

/******************* CELL 2151 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2151 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2055]),
			.N(gen[2056]),
			.NE(gen[2057]),

			.O(gen[2150]),
			.E(gen[2152]),

			.SO(gen[2245]),
			.S(gen[2246]),
			.SE(gen[2247]),

			.SELF(gen[2151]),
			.cell_state(gen[2151])
		); 

/******************* CELL 2152 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2152 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2056]),
			.N(gen[2057]),
			.NE(gen[2058]),

			.O(gen[2151]),
			.E(gen[2153]),

			.SO(gen[2246]),
			.S(gen[2247]),
			.SE(gen[2248]),

			.SELF(gen[2152]),
			.cell_state(gen[2152])
		); 

/******************* CELL 2153 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2153 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2057]),
			.N(gen[2058]),
			.NE(gen[2059]),

			.O(gen[2152]),
			.E(gen[2154]),

			.SO(gen[2247]),
			.S(gen[2248]),
			.SE(gen[2249]),

			.SELF(gen[2153]),
			.cell_state(gen[2153])
		); 

/******************* CELL 2154 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2154 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2058]),
			.N(gen[2059]),
			.NE(gen[2060]),

			.O(gen[2153]),
			.E(gen[2155]),

			.SO(gen[2248]),
			.S(gen[2249]),
			.SE(gen[2250]),

			.SELF(gen[2154]),
			.cell_state(gen[2154])
		); 

/******************* CELL 2155 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2155 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2059]),
			.N(gen[2060]),
			.NE(gen[2061]),

			.O(gen[2154]),
			.E(gen[2156]),

			.SO(gen[2249]),
			.S(gen[2250]),
			.SE(gen[2251]),

			.SELF(gen[2155]),
			.cell_state(gen[2155])
		); 

/******************* CELL 2156 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2156 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2060]),
			.N(gen[2061]),
			.NE(gen[2062]),

			.O(gen[2155]),
			.E(gen[2157]),

			.SO(gen[2250]),
			.S(gen[2251]),
			.SE(gen[2252]),

			.SELF(gen[2156]),
			.cell_state(gen[2156])
		); 

/******************* CELL 2157 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2157 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2061]),
			.N(gen[2062]),
			.NE(gen[2063]),

			.O(gen[2156]),
			.E(gen[2158]),

			.SO(gen[2251]),
			.S(gen[2252]),
			.SE(gen[2253]),

			.SELF(gen[2157]),
			.cell_state(gen[2157])
		); 

/******************* CELL 2158 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2158 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2062]),
			.N(gen[2063]),
			.NE(gen[2064]),

			.O(gen[2157]),
			.E(gen[2159]),

			.SO(gen[2252]),
			.S(gen[2253]),
			.SE(gen[2254]),

			.SELF(gen[2158]),
			.cell_state(gen[2158])
		); 

/******************* CELL 2159 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2159 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2063]),
			.N(gen[2064]),
			.NE(gen[2065]),

			.O(gen[2158]),
			.E(gen[2160]),

			.SO(gen[2253]),
			.S(gen[2254]),
			.SE(gen[2255]),

			.SELF(gen[2159]),
			.cell_state(gen[2159])
		); 

/******************* CELL 2160 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2160 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2064]),
			.N(gen[2065]),
			.NE(gen[2066]),

			.O(gen[2159]),
			.E(gen[2161]),

			.SO(gen[2254]),
			.S(gen[2255]),
			.SE(gen[2256]),

			.SELF(gen[2160]),
			.cell_state(gen[2160])
		); 

/******************* CELL 2161 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2161 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2065]),
			.N(gen[2066]),
			.NE(gen[2067]),

			.O(gen[2160]),
			.E(gen[2162]),

			.SO(gen[2255]),
			.S(gen[2256]),
			.SE(gen[2257]),

			.SELF(gen[2161]),
			.cell_state(gen[2161])
		); 

/******************* CELL 2162 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2162 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2066]),
			.N(gen[2067]),
			.NE(gen[2068]),

			.O(gen[2161]),
			.E(gen[2163]),

			.SO(gen[2256]),
			.S(gen[2257]),
			.SE(gen[2258]),

			.SELF(gen[2162]),
			.cell_state(gen[2162])
		); 

/******************* CELL 2163 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2163 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2067]),
			.N(gen[2068]),
			.NE(gen[2069]),

			.O(gen[2162]),
			.E(gen[2164]),

			.SO(gen[2257]),
			.S(gen[2258]),
			.SE(gen[2259]),

			.SELF(gen[2163]),
			.cell_state(gen[2163])
		); 

/******************* CELL 2164 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2164 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2068]),
			.N(gen[2069]),
			.NE(gen[2070]),

			.O(gen[2163]),
			.E(gen[2165]),

			.SO(gen[2258]),
			.S(gen[2259]),
			.SE(gen[2260]),

			.SELF(gen[2164]),
			.cell_state(gen[2164])
		); 

/******************* CELL 2165 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2165 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2069]),
			.N(gen[2070]),
			.NE(gen[2071]),

			.O(gen[2164]),
			.E(gen[2166]),

			.SO(gen[2259]),
			.S(gen[2260]),
			.SE(gen[2261]),

			.SELF(gen[2165]),
			.cell_state(gen[2165])
		); 

/******************* CELL 2166 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2166 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2070]),
			.N(gen[2071]),
			.NE(gen[2072]),

			.O(gen[2165]),
			.E(gen[2167]),

			.SO(gen[2260]),
			.S(gen[2261]),
			.SE(gen[2262]),

			.SELF(gen[2166]),
			.cell_state(gen[2166])
		); 

/******************* CELL 2167 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2167 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2071]),
			.N(gen[2072]),
			.NE(gen[2073]),

			.O(gen[2166]),
			.E(gen[2168]),

			.SO(gen[2261]),
			.S(gen[2262]),
			.SE(gen[2263]),

			.SELF(gen[2167]),
			.cell_state(gen[2167])
		); 

/******************* CELL 2168 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2168 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2072]),
			.N(gen[2073]),
			.NE(gen[2074]),

			.O(gen[2167]),
			.E(gen[2169]),

			.SO(gen[2262]),
			.S(gen[2263]),
			.SE(gen[2264]),

			.SELF(gen[2168]),
			.cell_state(gen[2168])
		); 

/******************* CELL 2169 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2169 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2073]),
			.N(gen[2074]),
			.NE(gen[2075]),

			.O(gen[2168]),
			.E(gen[2170]),

			.SO(gen[2263]),
			.S(gen[2264]),
			.SE(gen[2265]),

			.SELF(gen[2169]),
			.cell_state(gen[2169])
		); 

/******************* CELL 2170 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2170 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2074]),
			.N(gen[2075]),
			.NE(gen[2076]),

			.O(gen[2169]),
			.E(gen[2171]),

			.SO(gen[2264]),
			.S(gen[2265]),
			.SE(gen[2266]),

			.SELF(gen[2170]),
			.cell_state(gen[2170])
		); 

/******************* CELL 2171 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2171 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2075]),
			.N(gen[2076]),
			.NE(gen[2077]),

			.O(gen[2170]),
			.E(gen[2172]),

			.SO(gen[2265]),
			.S(gen[2266]),
			.SE(gen[2267]),

			.SELF(gen[2171]),
			.cell_state(gen[2171])
		); 

/******************* CELL 2172 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2172 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2076]),
			.N(gen[2077]),
			.NE(gen[2078]),

			.O(gen[2171]),
			.E(gen[2173]),

			.SO(gen[2266]),
			.S(gen[2267]),
			.SE(gen[2268]),

			.SELF(gen[2172]),
			.cell_state(gen[2172])
		); 

/******************* CELL 2173 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2173 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2077]),
			.N(gen[2078]),
			.NE(gen[2079]),

			.O(gen[2172]),
			.E(gen[2174]),

			.SO(gen[2267]),
			.S(gen[2268]),
			.SE(gen[2269]),

			.SELF(gen[2173]),
			.cell_state(gen[2173])
		); 

/******************* CELL 2174 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2174 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2078]),
			.N(gen[2079]),
			.NE(gen[2080]),

			.O(gen[2173]),
			.E(gen[2175]),

			.SO(gen[2268]),
			.S(gen[2269]),
			.SE(gen[2270]),

			.SELF(gen[2174]),
			.cell_state(gen[2174])
		); 

/******************* CELL 2175 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2175 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2079]),
			.N(gen[2080]),
			.NE(gen[2081]),

			.O(gen[2174]),
			.E(gen[2176]),

			.SO(gen[2269]),
			.S(gen[2270]),
			.SE(gen[2271]),

			.SELF(gen[2175]),
			.cell_state(gen[2175])
		); 

/******************* CELL 2176 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2176 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2080]),
			.N(gen[2081]),
			.NE(gen[2082]),

			.O(gen[2175]),
			.E(gen[2177]),

			.SO(gen[2270]),
			.S(gen[2271]),
			.SE(gen[2272]),

			.SELF(gen[2176]),
			.cell_state(gen[2176])
		); 

/******************* CELL 2177 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2177 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2081]),
			.N(gen[2082]),
			.NE(gen[2083]),

			.O(gen[2176]),
			.E(gen[2178]),

			.SO(gen[2271]),
			.S(gen[2272]),
			.SE(gen[2273]),

			.SELF(gen[2177]),
			.cell_state(gen[2177])
		); 

/******************* CELL 2178 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2178 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2082]),
			.N(gen[2083]),
			.NE(gen[2084]),

			.O(gen[2177]),
			.E(gen[2179]),

			.SO(gen[2272]),
			.S(gen[2273]),
			.SE(gen[2274]),

			.SELF(gen[2178]),
			.cell_state(gen[2178])
		); 

/******************* CELL 2179 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2179 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2083]),
			.N(gen[2084]),
			.NE(gen[2085]),

			.O(gen[2178]),
			.E(gen[2180]),

			.SO(gen[2273]),
			.S(gen[2274]),
			.SE(gen[2275]),

			.SELF(gen[2179]),
			.cell_state(gen[2179])
		); 

/******************* CELL 2180 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2180 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2084]),
			.N(gen[2085]),
			.NE(gen[2086]),

			.O(gen[2179]),
			.E(gen[2181]),

			.SO(gen[2274]),
			.S(gen[2275]),
			.SE(gen[2276]),

			.SELF(gen[2180]),
			.cell_state(gen[2180])
		); 

/******************* CELL 2181 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2181 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2085]),
			.N(gen[2086]),
			.NE(gen[2087]),

			.O(gen[2180]),
			.E(gen[2182]),

			.SO(gen[2275]),
			.S(gen[2276]),
			.SE(gen[2277]),

			.SELF(gen[2181]),
			.cell_state(gen[2181])
		); 

/******************* CELL 2182 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2182 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2086]),
			.N(gen[2087]),
			.NE(gen[2088]),

			.O(gen[2181]),
			.E(gen[2183]),

			.SO(gen[2276]),
			.S(gen[2277]),
			.SE(gen[2278]),

			.SELF(gen[2182]),
			.cell_state(gen[2182])
		); 

/******************* CELL 2183 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2183 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2087]),
			.N(gen[2088]),
			.NE(gen[2089]),

			.O(gen[2182]),
			.E(gen[2184]),

			.SO(gen[2277]),
			.S(gen[2278]),
			.SE(gen[2279]),

			.SELF(gen[2183]),
			.cell_state(gen[2183])
		); 

/******************* CELL 2184 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2184 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2088]),
			.N(gen[2089]),
			.NE(gen[2088]),

			.O(gen[2183]),
			.E(gen[2183]),

			.SO(gen[2278]),
			.S(gen[2279]),
			.SE(gen[2278]),

			.SELF(gen[2184]),
			.cell_state(gen[2184])
		); 

/******************* CELL 2185 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2185 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2091]),
			.N(gen[2090]),
			.NE(gen[2091]),

			.O(gen[2186]),
			.E(gen[2186]),

			.SO(gen[2281]),
			.S(gen[2280]),
			.SE(gen[2281]),

			.SELF(gen[2185]),
			.cell_state(gen[2185])
		); 

/******************* CELL 2186 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2186 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2090]),
			.N(gen[2091]),
			.NE(gen[2092]),

			.O(gen[2185]),
			.E(gen[2187]),

			.SO(gen[2280]),
			.S(gen[2281]),
			.SE(gen[2282]),

			.SELF(gen[2186]),
			.cell_state(gen[2186])
		); 

/******************* CELL 2187 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2187 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2091]),
			.N(gen[2092]),
			.NE(gen[2093]),

			.O(gen[2186]),
			.E(gen[2188]),

			.SO(gen[2281]),
			.S(gen[2282]),
			.SE(gen[2283]),

			.SELF(gen[2187]),
			.cell_state(gen[2187])
		); 

/******************* CELL 2188 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2188 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2092]),
			.N(gen[2093]),
			.NE(gen[2094]),

			.O(gen[2187]),
			.E(gen[2189]),

			.SO(gen[2282]),
			.S(gen[2283]),
			.SE(gen[2284]),

			.SELF(gen[2188]),
			.cell_state(gen[2188])
		); 

/******************* CELL 2189 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2189 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2093]),
			.N(gen[2094]),
			.NE(gen[2095]),

			.O(gen[2188]),
			.E(gen[2190]),

			.SO(gen[2283]),
			.S(gen[2284]),
			.SE(gen[2285]),

			.SELF(gen[2189]),
			.cell_state(gen[2189])
		); 

/******************* CELL 2190 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2190 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2094]),
			.N(gen[2095]),
			.NE(gen[2096]),

			.O(gen[2189]),
			.E(gen[2191]),

			.SO(gen[2284]),
			.S(gen[2285]),
			.SE(gen[2286]),

			.SELF(gen[2190]),
			.cell_state(gen[2190])
		); 

/******************* CELL 2191 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2191 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2095]),
			.N(gen[2096]),
			.NE(gen[2097]),

			.O(gen[2190]),
			.E(gen[2192]),

			.SO(gen[2285]),
			.S(gen[2286]),
			.SE(gen[2287]),

			.SELF(gen[2191]),
			.cell_state(gen[2191])
		); 

/******************* CELL 2192 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2192 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2096]),
			.N(gen[2097]),
			.NE(gen[2098]),

			.O(gen[2191]),
			.E(gen[2193]),

			.SO(gen[2286]),
			.S(gen[2287]),
			.SE(gen[2288]),

			.SELF(gen[2192]),
			.cell_state(gen[2192])
		); 

/******************* CELL 2193 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2193 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2097]),
			.N(gen[2098]),
			.NE(gen[2099]),

			.O(gen[2192]),
			.E(gen[2194]),

			.SO(gen[2287]),
			.S(gen[2288]),
			.SE(gen[2289]),

			.SELF(gen[2193]),
			.cell_state(gen[2193])
		); 

/******************* CELL 2194 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2194 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2098]),
			.N(gen[2099]),
			.NE(gen[2100]),

			.O(gen[2193]),
			.E(gen[2195]),

			.SO(gen[2288]),
			.S(gen[2289]),
			.SE(gen[2290]),

			.SELF(gen[2194]),
			.cell_state(gen[2194])
		); 

/******************* CELL 2195 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2195 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2099]),
			.N(gen[2100]),
			.NE(gen[2101]),

			.O(gen[2194]),
			.E(gen[2196]),

			.SO(gen[2289]),
			.S(gen[2290]),
			.SE(gen[2291]),

			.SELF(gen[2195]),
			.cell_state(gen[2195])
		); 

/******************* CELL 2196 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2196 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2100]),
			.N(gen[2101]),
			.NE(gen[2102]),

			.O(gen[2195]),
			.E(gen[2197]),

			.SO(gen[2290]),
			.S(gen[2291]),
			.SE(gen[2292]),

			.SELF(gen[2196]),
			.cell_state(gen[2196])
		); 

/******************* CELL 2197 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2197 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2101]),
			.N(gen[2102]),
			.NE(gen[2103]),

			.O(gen[2196]),
			.E(gen[2198]),

			.SO(gen[2291]),
			.S(gen[2292]),
			.SE(gen[2293]),

			.SELF(gen[2197]),
			.cell_state(gen[2197])
		); 

/******************* CELL 2198 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2198 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2102]),
			.N(gen[2103]),
			.NE(gen[2104]),

			.O(gen[2197]),
			.E(gen[2199]),

			.SO(gen[2292]),
			.S(gen[2293]),
			.SE(gen[2294]),

			.SELF(gen[2198]),
			.cell_state(gen[2198])
		); 

/******************* CELL 2199 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2199 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2103]),
			.N(gen[2104]),
			.NE(gen[2105]),

			.O(gen[2198]),
			.E(gen[2200]),

			.SO(gen[2293]),
			.S(gen[2294]),
			.SE(gen[2295]),

			.SELF(gen[2199]),
			.cell_state(gen[2199])
		); 

/******************* CELL 2200 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2200 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2104]),
			.N(gen[2105]),
			.NE(gen[2106]),

			.O(gen[2199]),
			.E(gen[2201]),

			.SO(gen[2294]),
			.S(gen[2295]),
			.SE(gen[2296]),

			.SELF(gen[2200]),
			.cell_state(gen[2200])
		); 

/******************* CELL 2201 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2201 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2105]),
			.N(gen[2106]),
			.NE(gen[2107]),

			.O(gen[2200]),
			.E(gen[2202]),

			.SO(gen[2295]),
			.S(gen[2296]),
			.SE(gen[2297]),

			.SELF(gen[2201]),
			.cell_state(gen[2201])
		); 

/******************* CELL 2202 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2202 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2106]),
			.N(gen[2107]),
			.NE(gen[2108]),

			.O(gen[2201]),
			.E(gen[2203]),

			.SO(gen[2296]),
			.S(gen[2297]),
			.SE(gen[2298]),

			.SELF(gen[2202]),
			.cell_state(gen[2202])
		); 

/******************* CELL 2203 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2203 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2107]),
			.N(gen[2108]),
			.NE(gen[2109]),

			.O(gen[2202]),
			.E(gen[2204]),

			.SO(gen[2297]),
			.S(gen[2298]),
			.SE(gen[2299]),

			.SELF(gen[2203]),
			.cell_state(gen[2203])
		); 

/******************* CELL 2204 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2204 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2108]),
			.N(gen[2109]),
			.NE(gen[2110]),

			.O(gen[2203]),
			.E(gen[2205]),

			.SO(gen[2298]),
			.S(gen[2299]),
			.SE(gen[2300]),

			.SELF(gen[2204]),
			.cell_state(gen[2204])
		); 

/******************* CELL 2205 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2205 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2109]),
			.N(gen[2110]),
			.NE(gen[2111]),

			.O(gen[2204]),
			.E(gen[2206]),

			.SO(gen[2299]),
			.S(gen[2300]),
			.SE(gen[2301]),

			.SELF(gen[2205]),
			.cell_state(gen[2205])
		); 

/******************* CELL 2206 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2206 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2110]),
			.N(gen[2111]),
			.NE(gen[2112]),

			.O(gen[2205]),
			.E(gen[2207]),

			.SO(gen[2300]),
			.S(gen[2301]),
			.SE(gen[2302]),

			.SELF(gen[2206]),
			.cell_state(gen[2206])
		); 

/******************* CELL 2207 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2207 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2111]),
			.N(gen[2112]),
			.NE(gen[2113]),

			.O(gen[2206]),
			.E(gen[2208]),

			.SO(gen[2301]),
			.S(gen[2302]),
			.SE(gen[2303]),

			.SELF(gen[2207]),
			.cell_state(gen[2207])
		); 

/******************* CELL 2208 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2208 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2112]),
			.N(gen[2113]),
			.NE(gen[2114]),

			.O(gen[2207]),
			.E(gen[2209]),

			.SO(gen[2302]),
			.S(gen[2303]),
			.SE(gen[2304]),

			.SELF(gen[2208]),
			.cell_state(gen[2208])
		); 

/******************* CELL 2209 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2209 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2113]),
			.N(gen[2114]),
			.NE(gen[2115]),

			.O(gen[2208]),
			.E(gen[2210]),

			.SO(gen[2303]),
			.S(gen[2304]),
			.SE(gen[2305]),

			.SELF(gen[2209]),
			.cell_state(gen[2209])
		); 

/******************* CELL 2210 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2210 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2114]),
			.N(gen[2115]),
			.NE(gen[2116]),

			.O(gen[2209]),
			.E(gen[2211]),

			.SO(gen[2304]),
			.S(gen[2305]),
			.SE(gen[2306]),

			.SELF(gen[2210]),
			.cell_state(gen[2210])
		); 

/******************* CELL 2211 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2211 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2115]),
			.N(gen[2116]),
			.NE(gen[2117]),

			.O(gen[2210]),
			.E(gen[2212]),

			.SO(gen[2305]),
			.S(gen[2306]),
			.SE(gen[2307]),

			.SELF(gen[2211]),
			.cell_state(gen[2211])
		); 

/******************* CELL 2212 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2212 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2116]),
			.N(gen[2117]),
			.NE(gen[2118]),

			.O(gen[2211]),
			.E(gen[2213]),

			.SO(gen[2306]),
			.S(gen[2307]),
			.SE(gen[2308]),

			.SELF(gen[2212]),
			.cell_state(gen[2212])
		); 

/******************* CELL 2213 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2213 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2117]),
			.N(gen[2118]),
			.NE(gen[2119]),

			.O(gen[2212]),
			.E(gen[2214]),

			.SO(gen[2307]),
			.S(gen[2308]),
			.SE(gen[2309]),

			.SELF(gen[2213]),
			.cell_state(gen[2213])
		); 

/******************* CELL 2214 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2214 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2118]),
			.N(gen[2119]),
			.NE(gen[2120]),

			.O(gen[2213]),
			.E(gen[2215]),

			.SO(gen[2308]),
			.S(gen[2309]),
			.SE(gen[2310]),

			.SELF(gen[2214]),
			.cell_state(gen[2214])
		); 

/******************* CELL 2215 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2215 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2119]),
			.N(gen[2120]),
			.NE(gen[2121]),

			.O(gen[2214]),
			.E(gen[2216]),

			.SO(gen[2309]),
			.S(gen[2310]),
			.SE(gen[2311]),

			.SELF(gen[2215]),
			.cell_state(gen[2215])
		); 

/******************* CELL 2216 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2216 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2120]),
			.N(gen[2121]),
			.NE(gen[2122]),

			.O(gen[2215]),
			.E(gen[2217]),

			.SO(gen[2310]),
			.S(gen[2311]),
			.SE(gen[2312]),

			.SELF(gen[2216]),
			.cell_state(gen[2216])
		); 

/******************* CELL 2217 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2217 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2121]),
			.N(gen[2122]),
			.NE(gen[2123]),

			.O(gen[2216]),
			.E(gen[2218]),

			.SO(gen[2311]),
			.S(gen[2312]),
			.SE(gen[2313]),

			.SELF(gen[2217]),
			.cell_state(gen[2217])
		); 

/******************* CELL 2218 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2218 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2122]),
			.N(gen[2123]),
			.NE(gen[2124]),

			.O(gen[2217]),
			.E(gen[2219]),

			.SO(gen[2312]),
			.S(gen[2313]),
			.SE(gen[2314]),

			.SELF(gen[2218]),
			.cell_state(gen[2218])
		); 

/******************* CELL 2219 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2219 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2123]),
			.N(gen[2124]),
			.NE(gen[2125]),

			.O(gen[2218]),
			.E(gen[2220]),

			.SO(gen[2313]),
			.S(gen[2314]),
			.SE(gen[2315]),

			.SELF(gen[2219]),
			.cell_state(gen[2219])
		); 

/******************* CELL 2220 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2220 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2124]),
			.N(gen[2125]),
			.NE(gen[2126]),

			.O(gen[2219]),
			.E(gen[2221]),

			.SO(gen[2314]),
			.S(gen[2315]),
			.SE(gen[2316]),

			.SELF(gen[2220]),
			.cell_state(gen[2220])
		); 

/******************* CELL 2221 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2221 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2125]),
			.N(gen[2126]),
			.NE(gen[2127]),

			.O(gen[2220]),
			.E(gen[2222]),

			.SO(gen[2315]),
			.S(gen[2316]),
			.SE(gen[2317]),

			.SELF(gen[2221]),
			.cell_state(gen[2221])
		); 

/******************* CELL 2222 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2222 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2126]),
			.N(gen[2127]),
			.NE(gen[2128]),

			.O(gen[2221]),
			.E(gen[2223]),

			.SO(gen[2316]),
			.S(gen[2317]),
			.SE(gen[2318]),

			.SELF(gen[2222]),
			.cell_state(gen[2222])
		); 

/******************* CELL 2223 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2223 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2127]),
			.N(gen[2128]),
			.NE(gen[2129]),

			.O(gen[2222]),
			.E(gen[2224]),

			.SO(gen[2317]),
			.S(gen[2318]),
			.SE(gen[2319]),

			.SELF(gen[2223]),
			.cell_state(gen[2223])
		); 

/******************* CELL 2224 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2224 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2128]),
			.N(gen[2129]),
			.NE(gen[2130]),

			.O(gen[2223]),
			.E(gen[2225]),

			.SO(gen[2318]),
			.S(gen[2319]),
			.SE(gen[2320]),

			.SELF(gen[2224]),
			.cell_state(gen[2224])
		); 

/******************* CELL 2225 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2225 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2129]),
			.N(gen[2130]),
			.NE(gen[2131]),

			.O(gen[2224]),
			.E(gen[2226]),

			.SO(gen[2319]),
			.S(gen[2320]),
			.SE(gen[2321]),

			.SELF(gen[2225]),
			.cell_state(gen[2225])
		); 

/******************* CELL 2226 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2226 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2130]),
			.N(gen[2131]),
			.NE(gen[2132]),

			.O(gen[2225]),
			.E(gen[2227]),

			.SO(gen[2320]),
			.S(gen[2321]),
			.SE(gen[2322]),

			.SELF(gen[2226]),
			.cell_state(gen[2226])
		); 

/******************* CELL 2227 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2227 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2131]),
			.N(gen[2132]),
			.NE(gen[2133]),

			.O(gen[2226]),
			.E(gen[2228]),

			.SO(gen[2321]),
			.S(gen[2322]),
			.SE(gen[2323]),

			.SELF(gen[2227]),
			.cell_state(gen[2227])
		); 

/******************* CELL 2228 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2228 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2132]),
			.N(gen[2133]),
			.NE(gen[2134]),

			.O(gen[2227]),
			.E(gen[2229]),

			.SO(gen[2322]),
			.S(gen[2323]),
			.SE(gen[2324]),

			.SELF(gen[2228]),
			.cell_state(gen[2228])
		); 

/******************* CELL 2229 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2229 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2133]),
			.N(gen[2134]),
			.NE(gen[2135]),

			.O(gen[2228]),
			.E(gen[2230]),

			.SO(gen[2323]),
			.S(gen[2324]),
			.SE(gen[2325]),

			.SELF(gen[2229]),
			.cell_state(gen[2229])
		); 

/******************* CELL 2230 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2230 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2134]),
			.N(gen[2135]),
			.NE(gen[2136]),

			.O(gen[2229]),
			.E(gen[2231]),

			.SO(gen[2324]),
			.S(gen[2325]),
			.SE(gen[2326]),

			.SELF(gen[2230]),
			.cell_state(gen[2230])
		); 

/******************* CELL 2231 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2231 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2135]),
			.N(gen[2136]),
			.NE(gen[2137]),

			.O(gen[2230]),
			.E(gen[2232]),

			.SO(gen[2325]),
			.S(gen[2326]),
			.SE(gen[2327]),

			.SELF(gen[2231]),
			.cell_state(gen[2231])
		); 

/******************* CELL 2232 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2232 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2136]),
			.N(gen[2137]),
			.NE(gen[2138]),

			.O(gen[2231]),
			.E(gen[2233]),

			.SO(gen[2326]),
			.S(gen[2327]),
			.SE(gen[2328]),

			.SELF(gen[2232]),
			.cell_state(gen[2232])
		); 

/******************* CELL 2233 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2233 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2137]),
			.N(gen[2138]),
			.NE(gen[2139]),

			.O(gen[2232]),
			.E(gen[2234]),

			.SO(gen[2327]),
			.S(gen[2328]),
			.SE(gen[2329]),

			.SELF(gen[2233]),
			.cell_state(gen[2233])
		); 

/******************* CELL 2234 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2234 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2138]),
			.N(gen[2139]),
			.NE(gen[2140]),

			.O(gen[2233]),
			.E(gen[2235]),

			.SO(gen[2328]),
			.S(gen[2329]),
			.SE(gen[2330]),

			.SELF(gen[2234]),
			.cell_state(gen[2234])
		); 

/******************* CELL 2235 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2235 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2139]),
			.N(gen[2140]),
			.NE(gen[2141]),

			.O(gen[2234]),
			.E(gen[2236]),

			.SO(gen[2329]),
			.S(gen[2330]),
			.SE(gen[2331]),

			.SELF(gen[2235]),
			.cell_state(gen[2235])
		); 

/******************* CELL 2236 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2236 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2140]),
			.N(gen[2141]),
			.NE(gen[2142]),

			.O(gen[2235]),
			.E(gen[2237]),

			.SO(gen[2330]),
			.S(gen[2331]),
			.SE(gen[2332]),

			.SELF(gen[2236]),
			.cell_state(gen[2236])
		); 

/******************* CELL 2237 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2237 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2141]),
			.N(gen[2142]),
			.NE(gen[2143]),

			.O(gen[2236]),
			.E(gen[2238]),

			.SO(gen[2331]),
			.S(gen[2332]),
			.SE(gen[2333]),

			.SELF(gen[2237]),
			.cell_state(gen[2237])
		); 

/******************* CELL 2238 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2238 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2142]),
			.N(gen[2143]),
			.NE(gen[2144]),

			.O(gen[2237]),
			.E(gen[2239]),

			.SO(gen[2332]),
			.S(gen[2333]),
			.SE(gen[2334]),

			.SELF(gen[2238]),
			.cell_state(gen[2238])
		); 

/******************* CELL 2239 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2239 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2143]),
			.N(gen[2144]),
			.NE(gen[2145]),

			.O(gen[2238]),
			.E(gen[2240]),

			.SO(gen[2333]),
			.S(gen[2334]),
			.SE(gen[2335]),

			.SELF(gen[2239]),
			.cell_state(gen[2239])
		); 

/******************* CELL 2240 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2240 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2144]),
			.N(gen[2145]),
			.NE(gen[2146]),

			.O(gen[2239]),
			.E(gen[2241]),

			.SO(gen[2334]),
			.S(gen[2335]),
			.SE(gen[2336]),

			.SELF(gen[2240]),
			.cell_state(gen[2240])
		); 

/******************* CELL 2241 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2241 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2145]),
			.N(gen[2146]),
			.NE(gen[2147]),

			.O(gen[2240]),
			.E(gen[2242]),

			.SO(gen[2335]),
			.S(gen[2336]),
			.SE(gen[2337]),

			.SELF(gen[2241]),
			.cell_state(gen[2241])
		); 

/******************* CELL 2242 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2242 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2146]),
			.N(gen[2147]),
			.NE(gen[2148]),

			.O(gen[2241]),
			.E(gen[2243]),

			.SO(gen[2336]),
			.S(gen[2337]),
			.SE(gen[2338]),

			.SELF(gen[2242]),
			.cell_state(gen[2242])
		); 

/******************* CELL 2243 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2243 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2147]),
			.N(gen[2148]),
			.NE(gen[2149]),

			.O(gen[2242]),
			.E(gen[2244]),

			.SO(gen[2337]),
			.S(gen[2338]),
			.SE(gen[2339]),

			.SELF(gen[2243]),
			.cell_state(gen[2243])
		); 

/******************* CELL 2244 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2244 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2148]),
			.N(gen[2149]),
			.NE(gen[2150]),

			.O(gen[2243]),
			.E(gen[2245]),

			.SO(gen[2338]),
			.S(gen[2339]),
			.SE(gen[2340]),

			.SELF(gen[2244]),
			.cell_state(gen[2244])
		); 

/******************* CELL 2245 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2245 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2149]),
			.N(gen[2150]),
			.NE(gen[2151]),

			.O(gen[2244]),
			.E(gen[2246]),

			.SO(gen[2339]),
			.S(gen[2340]),
			.SE(gen[2341]),

			.SELF(gen[2245]),
			.cell_state(gen[2245])
		); 

/******************* CELL 2246 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2246 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2150]),
			.N(gen[2151]),
			.NE(gen[2152]),

			.O(gen[2245]),
			.E(gen[2247]),

			.SO(gen[2340]),
			.S(gen[2341]),
			.SE(gen[2342]),

			.SELF(gen[2246]),
			.cell_state(gen[2246])
		); 

/******************* CELL 2247 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2247 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2151]),
			.N(gen[2152]),
			.NE(gen[2153]),

			.O(gen[2246]),
			.E(gen[2248]),

			.SO(gen[2341]),
			.S(gen[2342]),
			.SE(gen[2343]),

			.SELF(gen[2247]),
			.cell_state(gen[2247])
		); 

/******************* CELL 2248 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2248 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2152]),
			.N(gen[2153]),
			.NE(gen[2154]),

			.O(gen[2247]),
			.E(gen[2249]),

			.SO(gen[2342]),
			.S(gen[2343]),
			.SE(gen[2344]),

			.SELF(gen[2248]),
			.cell_state(gen[2248])
		); 

/******************* CELL 2249 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2249 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2153]),
			.N(gen[2154]),
			.NE(gen[2155]),

			.O(gen[2248]),
			.E(gen[2250]),

			.SO(gen[2343]),
			.S(gen[2344]),
			.SE(gen[2345]),

			.SELF(gen[2249]),
			.cell_state(gen[2249])
		); 

/******************* CELL 2250 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2250 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2154]),
			.N(gen[2155]),
			.NE(gen[2156]),

			.O(gen[2249]),
			.E(gen[2251]),

			.SO(gen[2344]),
			.S(gen[2345]),
			.SE(gen[2346]),

			.SELF(gen[2250]),
			.cell_state(gen[2250])
		); 

/******************* CELL 2251 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2251 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2155]),
			.N(gen[2156]),
			.NE(gen[2157]),

			.O(gen[2250]),
			.E(gen[2252]),

			.SO(gen[2345]),
			.S(gen[2346]),
			.SE(gen[2347]),

			.SELF(gen[2251]),
			.cell_state(gen[2251])
		); 

/******************* CELL 2252 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2252 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2156]),
			.N(gen[2157]),
			.NE(gen[2158]),

			.O(gen[2251]),
			.E(gen[2253]),

			.SO(gen[2346]),
			.S(gen[2347]),
			.SE(gen[2348]),

			.SELF(gen[2252]),
			.cell_state(gen[2252])
		); 

/******************* CELL 2253 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2253 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2157]),
			.N(gen[2158]),
			.NE(gen[2159]),

			.O(gen[2252]),
			.E(gen[2254]),

			.SO(gen[2347]),
			.S(gen[2348]),
			.SE(gen[2349]),

			.SELF(gen[2253]),
			.cell_state(gen[2253])
		); 

/******************* CELL 2254 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2254 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2158]),
			.N(gen[2159]),
			.NE(gen[2160]),

			.O(gen[2253]),
			.E(gen[2255]),

			.SO(gen[2348]),
			.S(gen[2349]),
			.SE(gen[2350]),

			.SELF(gen[2254]),
			.cell_state(gen[2254])
		); 

/******************* CELL 2255 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2255 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2159]),
			.N(gen[2160]),
			.NE(gen[2161]),

			.O(gen[2254]),
			.E(gen[2256]),

			.SO(gen[2349]),
			.S(gen[2350]),
			.SE(gen[2351]),

			.SELF(gen[2255]),
			.cell_state(gen[2255])
		); 

/******************* CELL 2256 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2256 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2160]),
			.N(gen[2161]),
			.NE(gen[2162]),

			.O(gen[2255]),
			.E(gen[2257]),

			.SO(gen[2350]),
			.S(gen[2351]),
			.SE(gen[2352]),

			.SELF(gen[2256]),
			.cell_state(gen[2256])
		); 

/******************* CELL 2257 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2257 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2161]),
			.N(gen[2162]),
			.NE(gen[2163]),

			.O(gen[2256]),
			.E(gen[2258]),

			.SO(gen[2351]),
			.S(gen[2352]),
			.SE(gen[2353]),

			.SELF(gen[2257]),
			.cell_state(gen[2257])
		); 

/******************* CELL 2258 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2258 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2162]),
			.N(gen[2163]),
			.NE(gen[2164]),

			.O(gen[2257]),
			.E(gen[2259]),

			.SO(gen[2352]),
			.S(gen[2353]),
			.SE(gen[2354]),

			.SELF(gen[2258]),
			.cell_state(gen[2258])
		); 

/******************* CELL 2259 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2259 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2163]),
			.N(gen[2164]),
			.NE(gen[2165]),

			.O(gen[2258]),
			.E(gen[2260]),

			.SO(gen[2353]),
			.S(gen[2354]),
			.SE(gen[2355]),

			.SELF(gen[2259]),
			.cell_state(gen[2259])
		); 

/******************* CELL 2260 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2260 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2164]),
			.N(gen[2165]),
			.NE(gen[2166]),

			.O(gen[2259]),
			.E(gen[2261]),

			.SO(gen[2354]),
			.S(gen[2355]),
			.SE(gen[2356]),

			.SELF(gen[2260]),
			.cell_state(gen[2260])
		); 

/******************* CELL 2261 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2261 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2165]),
			.N(gen[2166]),
			.NE(gen[2167]),

			.O(gen[2260]),
			.E(gen[2262]),

			.SO(gen[2355]),
			.S(gen[2356]),
			.SE(gen[2357]),

			.SELF(gen[2261]),
			.cell_state(gen[2261])
		); 

/******************* CELL 2262 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2262 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2166]),
			.N(gen[2167]),
			.NE(gen[2168]),

			.O(gen[2261]),
			.E(gen[2263]),

			.SO(gen[2356]),
			.S(gen[2357]),
			.SE(gen[2358]),

			.SELF(gen[2262]),
			.cell_state(gen[2262])
		); 

/******************* CELL 2263 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2263 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2167]),
			.N(gen[2168]),
			.NE(gen[2169]),

			.O(gen[2262]),
			.E(gen[2264]),

			.SO(gen[2357]),
			.S(gen[2358]),
			.SE(gen[2359]),

			.SELF(gen[2263]),
			.cell_state(gen[2263])
		); 

/******************* CELL 2264 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2264 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2168]),
			.N(gen[2169]),
			.NE(gen[2170]),

			.O(gen[2263]),
			.E(gen[2265]),

			.SO(gen[2358]),
			.S(gen[2359]),
			.SE(gen[2360]),

			.SELF(gen[2264]),
			.cell_state(gen[2264])
		); 

/******************* CELL 2265 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2265 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2169]),
			.N(gen[2170]),
			.NE(gen[2171]),

			.O(gen[2264]),
			.E(gen[2266]),

			.SO(gen[2359]),
			.S(gen[2360]),
			.SE(gen[2361]),

			.SELF(gen[2265]),
			.cell_state(gen[2265])
		); 

/******************* CELL 2266 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2266 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2170]),
			.N(gen[2171]),
			.NE(gen[2172]),

			.O(gen[2265]),
			.E(gen[2267]),

			.SO(gen[2360]),
			.S(gen[2361]),
			.SE(gen[2362]),

			.SELF(gen[2266]),
			.cell_state(gen[2266])
		); 

/******************* CELL 2267 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2267 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2171]),
			.N(gen[2172]),
			.NE(gen[2173]),

			.O(gen[2266]),
			.E(gen[2268]),

			.SO(gen[2361]),
			.S(gen[2362]),
			.SE(gen[2363]),

			.SELF(gen[2267]),
			.cell_state(gen[2267])
		); 

/******************* CELL 2268 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2268 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2172]),
			.N(gen[2173]),
			.NE(gen[2174]),

			.O(gen[2267]),
			.E(gen[2269]),

			.SO(gen[2362]),
			.S(gen[2363]),
			.SE(gen[2364]),

			.SELF(gen[2268]),
			.cell_state(gen[2268])
		); 

/******************* CELL 2269 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2269 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2173]),
			.N(gen[2174]),
			.NE(gen[2175]),

			.O(gen[2268]),
			.E(gen[2270]),

			.SO(gen[2363]),
			.S(gen[2364]),
			.SE(gen[2365]),

			.SELF(gen[2269]),
			.cell_state(gen[2269])
		); 

/******************* CELL 2270 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2270 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2174]),
			.N(gen[2175]),
			.NE(gen[2176]),

			.O(gen[2269]),
			.E(gen[2271]),

			.SO(gen[2364]),
			.S(gen[2365]),
			.SE(gen[2366]),

			.SELF(gen[2270]),
			.cell_state(gen[2270])
		); 

/******************* CELL 2271 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2271 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2175]),
			.N(gen[2176]),
			.NE(gen[2177]),

			.O(gen[2270]),
			.E(gen[2272]),

			.SO(gen[2365]),
			.S(gen[2366]),
			.SE(gen[2367]),

			.SELF(gen[2271]),
			.cell_state(gen[2271])
		); 

/******************* CELL 2272 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2272 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2176]),
			.N(gen[2177]),
			.NE(gen[2178]),

			.O(gen[2271]),
			.E(gen[2273]),

			.SO(gen[2366]),
			.S(gen[2367]),
			.SE(gen[2368]),

			.SELF(gen[2272]),
			.cell_state(gen[2272])
		); 

/******************* CELL 2273 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2273 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2177]),
			.N(gen[2178]),
			.NE(gen[2179]),

			.O(gen[2272]),
			.E(gen[2274]),

			.SO(gen[2367]),
			.S(gen[2368]),
			.SE(gen[2369]),

			.SELF(gen[2273]),
			.cell_state(gen[2273])
		); 

/******************* CELL 2274 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2274 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2178]),
			.N(gen[2179]),
			.NE(gen[2180]),

			.O(gen[2273]),
			.E(gen[2275]),

			.SO(gen[2368]),
			.S(gen[2369]),
			.SE(gen[2370]),

			.SELF(gen[2274]),
			.cell_state(gen[2274])
		); 

/******************* CELL 2275 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2275 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2179]),
			.N(gen[2180]),
			.NE(gen[2181]),

			.O(gen[2274]),
			.E(gen[2276]),

			.SO(gen[2369]),
			.S(gen[2370]),
			.SE(gen[2371]),

			.SELF(gen[2275]),
			.cell_state(gen[2275])
		); 

/******************* CELL 2276 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2276 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2180]),
			.N(gen[2181]),
			.NE(gen[2182]),

			.O(gen[2275]),
			.E(gen[2277]),

			.SO(gen[2370]),
			.S(gen[2371]),
			.SE(gen[2372]),

			.SELF(gen[2276]),
			.cell_state(gen[2276])
		); 

/******************* CELL 2277 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2277 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2181]),
			.N(gen[2182]),
			.NE(gen[2183]),

			.O(gen[2276]),
			.E(gen[2278]),

			.SO(gen[2371]),
			.S(gen[2372]),
			.SE(gen[2373]),

			.SELF(gen[2277]),
			.cell_state(gen[2277])
		); 

/******************* CELL 2278 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2278 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2182]),
			.N(gen[2183]),
			.NE(gen[2184]),

			.O(gen[2277]),
			.E(gen[2279]),

			.SO(gen[2372]),
			.S(gen[2373]),
			.SE(gen[2374]),

			.SELF(gen[2278]),
			.cell_state(gen[2278])
		); 

/******************* CELL 2279 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2279 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2183]),
			.N(gen[2184]),
			.NE(gen[2183]),

			.O(gen[2278]),
			.E(gen[2278]),

			.SO(gen[2373]),
			.S(gen[2374]),
			.SE(gen[2373]),

			.SELF(gen[2279]),
			.cell_state(gen[2279])
		); 

/******************* CELL 2280 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2280 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2186]),
			.N(gen[2185]),
			.NE(gen[2186]),

			.O(gen[2281]),
			.E(gen[2281]),

			.SO(gen[2376]),
			.S(gen[2375]),
			.SE(gen[2376]),

			.SELF(gen[2280]),
			.cell_state(gen[2280])
		); 

/******************* CELL 2281 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2281 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2185]),
			.N(gen[2186]),
			.NE(gen[2187]),

			.O(gen[2280]),
			.E(gen[2282]),

			.SO(gen[2375]),
			.S(gen[2376]),
			.SE(gen[2377]),

			.SELF(gen[2281]),
			.cell_state(gen[2281])
		); 

/******************* CELL 2282 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2282 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2186]),
			.N(gen[2187]),
			.NE(gen[2188]),

			.O(gen[2281]),
			.E(gen[2283]),

			.SO(gen[2376]),
			.S(gen[2377]),
			.SE(gen[2378]),

			.SELF(gen[2282]),
			.cell_state(gen[2282])
		); 

/******************* CELL 2283 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2283 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2187]),
			.N(gen[2188]),
			.NE(gen[2189]),

			.O(gen[2282]),
			.E(gen[2284]),

			.SO(gen[2377]),
			.S(gen[2378]),
			.SE(gen[2379]),

			.SELF(gen[2283]),
			.cell_state(gen[2283])
		); 

/******************* CELL 2284 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2284 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2188]),
			.N(gen[2189]),
			.NE(gen[2190]),

			.O(gen[2283]),
			.E(gen[2285]),

			.SO(gen[2378]),
			.S(gen[2379]),
			.SE(gen[2380]),

			.SELF(gen[2284]),
			.cell_state(gen[2284])
		); 

/******************* CELL 2285 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2285 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2189]),
			.N(gen[2190]),
			.NE(gen[2191]),

			.O(gen[2284]),
			.E(gen[2286]),

			.SO(gen[2379]),
			.S(gen[2380]),
			.SE(gen[2381]),

			.SELF(gen[2285]),
			.cell_state(gen[2285])
		); 

/******************* CELL 2286 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2286 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2190]),
			.N(gen[2191]),
			.NE(gen[2192]),

			.O(gen[2285]),
			.E(gen[2287]),

			.SO(gen[2380]),
			.S(gen[2381]),
			.SE(gen[2382]),

			.SELF(gen[2286]),
			.cell_state(gen[2286])
		); 

/******************* CELL 2287 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2287 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2191]),
			.N(gen[2192]),
			.NE(gen[2193]),

			.O(gen[2286]),
			.E(gen[2288]),

			.SO(gen[2381]),
			.S(gen[2382]),
			.SE(gen[2383]),

			.SELF(gen[2287]),
			.cell_state(gen[2287])
		); 

/******************* CELL 2288 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2288 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2192]),
			.N(gen[2193]),
			.NE(gen[2194]),

			.O(gen[2287]),
			.E(gen[2289]),

			.SO(gen[2382]),
			.S(gen[2383]),
			.SE(gen[2384]),

			.SELF(gen[2288]),
			.cell_state(gen[2288])
		); 

/******************* CELL 2289 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2289 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2193]),
			.N(gen[2194]),
			.NE(gen[2195]),

			.O(gen[2288]),
			.E(gen[2290]),

			.SO(gen[2383]),
			.S(gen[2384]),
			.SE(gen[2385]),

			.SELF(gen[2289]),
			.cell_state(gen[2289])
		); 

/******************* CELL 2290 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2290 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2194]),
			.N(gen[2195]),
			.NE(gen[2196]),

			.O(gen[2289]),
			.E(gen[2291]),

			.SO(gen[2384]),
			.S(gen[2385]),
			.SE(gen[2386]),

			.SELF(gen[2290]),
			.cell_state(gen[2290])
		); 

/******************* CELL 2291 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2291 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2195]),
			.N(gen[2196]),
			.NE(gen[2197]),

			.O(gen[2290]),
			.E(gen[2292]),

			.SO(gen[2385]),
			.S(gen[2386]),
			.SE(gen[2387]),

			.SELF(gen[2291]),
			.cell_state(gen[2291])
		); 

/******************* CELL 2292 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2292 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2196]),
			.N(gen[2197]),
			.NE(gen[2198]),

			.O(gen[2291]),
			.E(gen[2293]),

			.SO(gen[2386]),
			.S(gen[2387]),
			.SE(gen[2388]),

			.SELF(gen[2292]),
			.cell_state(gen[2292])
		); 

/******************* CELL 2293 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2293 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2197]),
			.N(gen[2198]),
			.NE(gen[2199]),

			.O(gen[2292]),
			.E(gen[2294]),

			.SO(gen[2387]),
			.S(gen[2388]),
			.SE(gen[2389]),

			.SELF(gen[2293]),
			.cell_state(gen[2293])
		); 

/******************* CELL 2294 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2294 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2198]),
			.N(gen[2199]),
			.NE(gen[2200]),

			.O(gen[2293]),
			.E(gen[2295]),

			.SO(gen[2388]),
			.S(gen[2389]),
			.SE(gen[2390]),

			.SELF(gen[2294]),
			.cell_state(gen[2294])
		); 

/******************* CELL 2295 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2295 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2199]),
			.N(gen[2200]),
			.NE(gen[2201]),

			.O(gen[2294]),
			.E(gen[2296]),

			.SO(gen[2389]),
			.S(gen[2390]),
			.SE(gen[2391]),

			.SELF(gen[2295]),
			.cell_state(gen[2295])
		); 

/******************* CELL 2296 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2296 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2200]),
			.N(gen[2201]),
			.NE(gen[2202]),

			.O(gen[2295]),
			.E(gen[2297]),

			.SO(gen[2390]),
			.S(gen[2391]),
			.SE(gen[2392]),

			.SELF(gen[2296]),
			.cell_state(gen[2296])
		); 

/******************* CELL 2297 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2297 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2201]),
			.N(gen[2202]),
			.NE(gen[2203]),

			.O(gen[2296]),
			.E(gen[2298]),

			.SO(gen[2391]),
			.S(gen[2392]),
			.SE(gen[2393]),

			.SELF(gen[2297]),
			.cell_state(gen[2297])
		); 

/******************* CELL 2298 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2298 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2202]),
			.N(gen[2203]),
			.NE(gen[2204]),

			.O(gen[2297]),
			.E(gen[2299]),

			.SO(gen[2392]),
			.S(gen[2393]),
			.SE(gen[2394]),

			.SELF(gen[2298]),
			.cell_state(gen[2298])
		); 

/******************* CELL 2299 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2299 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2203]),
			.N(gen[2204]),
			.NE(gen[2205]),

			.O(gen[2298]),
			.E(gen[2300]),

			.SO(gen[2393]),
			.S(gen[2394]),
			.SE(gen[2395]),

			.SELF(gen[2299]),
			.cell_state(gen[2299])
		); 

/******************* CELL 2300 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2300 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2204]),
			.N(gen[2205]),
			.NE(gen[2206]),

			.O(gen[2299]),
			.E(gen[2301]),

			.SO(gen[2394]),
			.S(gen[2395]),
			.SE(gen[2396]),

			.SELF(gen[2300]),
			.cell_state(gen[2300])
		); 

/******************* CELL 2301 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2301 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2205]),
			.N(gen[2206]),
			.NE(gen[2207]),

			.O(gen[2300]),
			.E(gen[2302]),

			.SO(gen[2395]),
			.S(gen[2396]),
			.SE(gen[2397]),

			.SELF(gen[2301]),
			.cell_state(gen[2301])
		); 

/******************* CELL 2302 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2302 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2206]),
			.N(gen[2207]),
			.NE(gen[2208]),

			.O(gen[2301]),
			.E(gen[2303]),

			.SO(gen[2396]),
			.S(gen[2397]),
			.SE(gen[2398]),

			.SELF(gen[2302]),
			.cell_state(gen[2302])
		); 

/******************* CELL 2303 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2303 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2207]),
			.N(gen[2208]),
			.NE(gen[2209]),

			.O(gen[2302]),
			.E(gen[2304]),

			.SO(gen[2397]),
			.S(gen[2398]),
			.SE(gen[2399]),

			.SELF(gen[2303]),
			.cell_state(gen[2303])
		); 

/******************* CELL 2304 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2304 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2208]),
			.N(gen[2209]),
			.NE(gen[2210]),

			.O(gen[2303]),
			.E(gen[2305]),

			.SO(gen[2398]),
			.S(gen[2399]),
			.SE(gen[2400]),

			.SELF(gen[2304]),
			.cell_state(gen[2304])
		); 

/******************* CELL 2305 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2305 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2209]),
			.N(gen[2210]),
			.NE(gen[2211]),

			.O(gen[2304]),
			.E(gen[2306]),

			.SO(gen[2399]),
			.S(gen[2400]),
			.SE(gen[2401]),

			.SELF(gen[2305]),
			.cell_state(gen[2305])
		); 

/******************* CELL 2306 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2306 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2210]),
			.N(gen[2211]),
			.NE(gen[2212]),

			.O(gen[2305]),
			.E(gen[2307]),

			.SO(gen[2400]),
			.S(gen[2401]),
			.SE(gen[2402]),

			.SELF(gen[2306]),
			.cell_state(gen[2306])
		); 

/******************* CELL 2307 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2307 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2211]),
			.N(gen[2212]),
			.NE(gen[2213]),

			.O(gen[2306]),
			.E(gen[2308]),

			.SO(gen[2401]),
			.S(gen[2402]),
			.SE(gen[2403]),

			.SELF(gen[2307]),
			.cell_state(gen[2307])
		); 

/******************* CELL 2308 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2308 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2212]),
			.N(gen[2213]),
			.NE(gen[2214]),

			.O(gen[2307]),
			.E(gen[2309]),

			.SO(gen[2402]),
			.S(gen[2403]),
			.SE(gen[2404]),

			.SELF(gen[2308]),
			.cell_state(gen[2308])
		); 

/******************* CELL 2309 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2309 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2213]),
			.N(gen[2214]),
			.NE(gen[2215]),

			.O(gen[2308]),
			.E(gen[2310]),

			.SO(gen[2403]),
			.S(gen[2404]),
			.SE(gen[2405]),

			.SELF(gen[2309]),
			.cell_state(gen[2309])
		); 

/******************* CELL 2310 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2310 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2214]),
			.N(gen[2215]),
			.NE(gen[2216]),

			.O(gen[2309]),
			.E(gen[2311]),

			.SO(gen[2404]),
			.S(gen[2405]),
			.SE(gen[2406]),

			.SELF(gen[2310]),
			.cell_state(gen[2310])
		); 

/******************* CELL 2311 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2311 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2215]),
			.N(gen[2216]),
			.NE(gen[2217]),

			.O(gen[2310]),
			.E(gen[2312]),

			.SO(gen[2405]),
			.S(gen[2406]),
			.SE(gen[2407]),

			.SELF(gen[2311]),
			.cell_state(gen[2311])
		); 

/******************* CELL 2312 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2312 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2216]),
			.N(gen[2217]),
			.NE(gen[2218]),

			.O(gen[2311]),
			.E(gen[2313]),

			.SO(gen[2406]),
			.S(gen[2407]),
			.SE(gen[2408]),

			.SELF(gen[2312]),
			.cell_state(gen[2312])
		); 

/******************* CELL 2313 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2313 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2217]),
			.N(gen[2218]),
			.NE(gen[2219]),

			.O(gen[2312]),
			.E(gen[2314]),

			.SO(gen[2407]),
			.S(gen[2408]),
			.SE(gen[2409]),

			.SELF(gen[2313]),
			.cell_state(gen[2313])
		); 

/******************* CELL 2314 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2314 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2218]),
			.N(gen[2219]),
			.NE(gen[2220]),

			.O(gen[2313]),
			.E(gen[2315]),

			.SO(gen[2408]),
			.S(gen[2409]),
			.SE(gen[2410]),

			.SELF(gen[2314]),
			.cell_state(gen[2314])
		); 

/******************* CELL 2315 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2315 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2219]),
			.N(gen[2220]),
			.NE(gen[2221]),

			.O(gen[2314]),
			.E(gen[2316]),

			.SO(gen[2409]),
			.S(gen[2410]),
			.SE(gen[2411]),

			.SELF(gen[2315]),
			.cell_state(gen[2315])
		); 

/******************* CELL 2316 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2316 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2220]),
			.N(gen[2221]),
			.NE(gen[2222]),

			.O(gen[2315]),
			.E(gen[2317]),

			.SO(gen[2410]),
			.S(gen[2411]),
			.SE(gen[2412]),

			.SELF(gen[2316]),
			.cell_state(gen[2316])
		); 

/******************* CELL 2317 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2317 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2221]),
			.N(gen[2222]),
			.NE(gen[2223]),

			.O(gen[2316]),
			.E(gen[2318]),

			.SO(gen[2411]),
			.S(gen[2412]),
			.SE(gen[2413]),

			.SELF(gen[2317]),
			.cell_state(gen[2317])
		); 

/******************* CELL 2318 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2318 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2222]),
			.N(gen[2223]),
			.NE(gen[2224]),

			.O(gen[2317]),
			.E(gen[2319]),

			.SO(gen[2412]),
			.S(gen[2413]),
			.SE(gen[2414]),

			.SELF(gen[2318]),
			.cell_state(gen[2318])
		); 

/******************* CELL 2319 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2319 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2223]),
			.N(gen[2224]),
			.NE(gen[2225]),

			.O(gen[2318]),
			.E(gen[2320]),

			.SO(gen[2413]),
			.S(gen[2414]),
			.SE(gen[2415]),

			.SELF(gen[2319]),
			.cell_state(gen[2319])
		); 

/******************* CELL 2320 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2320 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2224]),
			.N(gen[2225]),
			.NE(gen[2226]),

			.O(gen[2319]),
			.E(gen[2321]),

			.SO(gen[2414]),
			.S(gen[2415]),
			.SE(gen[2416]),

			.SELF(gen[2320]),
			.cell_state(gen[2320])
		); 

/******************* CELL 2321 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2321 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2225]),
			.N(gen[2226]),
			.NE(gen[2227]),

			.O(gen[2320]),
			.E(gen[2322]),

			.SO(gen[2415]),
			.S(gen[2416]),
			.SE(gen[2417]),

			.SELF(gen[2321]),
			.cell_state(gen[2321])
		); 

/******************* CELL 2322 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2322 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2226]),
			.N(gen[2227]),
			.NE(gen[2228]),

			.O(gen[2321]),
			.E(gen[2323]),

			.SO(gen[2416]),
			.S(gen[2417]),
			.SE(gen[2418]),

			.SELF(gen[2322]),
			.cell_state(gen[2322])
		); 

/******************* CELL 2323 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2323 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2227]),
			.N(gen[2228]),
			.NE(gen[2229]),

			.O(gen[2322]),
			.E(gen[2324]),

			.SO(gen[2417]),
			.S(gen[2418]),
			.SE(gen[2419]),

			.SELF(gen[2323]),
			.cell_state(gen[2323])
		); 

/******************* CELL 2324 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2324 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2228]),
			.N(gen[2229]),
			.NE(gen[2230]),

			.O(gen[2323]),
			.E(gen[2325]),

			.SO(gen[2418]),
			.S(gen[2419]),
			.SE(gen[2420]),

			.SELF(gen[2324]),
			.cell_state(gen[2324])
		); 

/******************* CELL 2325 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2325 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2229]),
			.N(gen[2230]),
			.NE(gen[2231]),

			.O(gen[2324]),
			.E(gen[2326]),

			.SO(gen[2419]),
			.S(gen[2420]),
			.SE(gen[2421]),

			.SELF(gen[2325]),
			.cell_state(gen[2325])
		); 

/******************* CELL 2326 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2326 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2230]),
			.N(gen[2231]),
			.NE(gen[2232]),

			.O(gen[2325]),
			.E(gen[2327]),

			.SO(gen[2420]),
			.S(gen[2421]),
			.SE(gen[2422]),

			.SELF(gen[2326]),
			.cell_state(gen[2326])
		); 

/******************* CELL 2327 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2327 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2231]),
			.N(gen[2232]),
			.NE(gen[2233]),

			.O(gen[2326]),
			.E(gen[2328]),

			.SO(gen[2421]),
			.S(gen[2422]),
			.SE(gen[2423]),

			.SELF(gen[2327]),
			.cell_state(gen[2327])
		); 

/******************* CELL 2328 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2328 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2232]),
			.N(gen[2233]),
			.NE(gen[2234]),

			.O(gen[2327]),
			.E(gen[2329]),

			.SO(gen[2422]),
			.S(gen[2423]),
			.SE(gen[2424]),

			.SELF(gen[2328]),
			.cell_state(gen[2328])
		); 

/******************* CELL 2329 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2329 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2233]),
			.N(gen[2234]),
			.NE(gen[2235]),

			.O(gen[2328]),
			.E(gen[2330]),

			.SO(gen[2423]),
			.S(gen[2424]),
			.SE(gen[2425]),

			.SELF(gen[2329]),
			.cell_state(gen[2329])
		); 

/******************* CELL 2330 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2330 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2234]),
			.N(gen[2235]),
			.NE(gen[2236]),

			.O(gen[2329]),
			.E(gen[2331]),

			.SO(gen[2424]),
			.S(gen[2425]),
			.SE(gen[2426]),

			.SELF(gen[2330]),
			.cell_state(gen[2330])
		); 

/******************* CELL 2331 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2331 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2235]),
			.N(gen[2236]),
			.NE(gen[2237]),

			.O(gen[2330]),
			.E(gen[2332]),

			.SO(gen[2425]),
			.S(gen[2426]),
			.SE(gen[2427]),

			.SELF(gen[2331]),
			.cell_state(gen[2331])
		); 

/******************* CELL 2332 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2332 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2236]),
			.N(gen[2237]),
			.NE(gen[2238]),

			.O(gen[2331]),
			.E(gen[2333]),

			.SO(gen[2426]),
			.S(gen[2427]),
			.SE(gen[2428]),

			.SELF(gen[2332]),
			.cell_state(gen[2332])
		); 

/******************* CELL 2333 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2333 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2237]),
			.N(gen[2238]),
			.NE(gen[2239]),

			.O(gen[2332]),
			.E(gen[2334]),

			.SO(gen[2427]),
			.S(gen[2428]),
			.SE(gen[2429]),

			.SELF(gen[2333]),
			.cell_state(gen[2333])
		); 

/******************* CELL 2334 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2334 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2238]),
			.N(gen[2239]),
			.NE(gen[2240]),

			.O(gen[2333]),
			.E(gen[2335]),

			.SO(gen[2428]),
			.S(gen[2429]),
			.SE(gen[2430]),

			.SELF(gen[2334]),
			.cell_state(gen[2334])
		); 

/******************* CELL 2335 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2335 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2239]),
			.N(gen[2240]),
			.NE(gen[2241]),

			.O(gen[2334]),
			.E(gen[2336]),

			.SO(gen[2429]),
			.S(gen[2430]),
			.SE(gen[2431]),

			.SELF(gen[2335]),
			.cell_state(gen[2335])
		); 

/******************* CELL 2336 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2336 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2240]),
			.N(gen[2241]),
			.NE(gen[2242]),

			.O(gen[2335]),
			.E(gen[2337]),

			.SO(gen[2430]),
			.S(gen[2431]),
			.SE(gen[2432]),

			.SELF(gen[2336]),
			.cell_state(gen[2336])
		); 

/******************* CELL 2337 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2337 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2241]),
			.N(gen[2242]),
			.NE(gen[2243]),

			.O(gen[2336]),
			.E(gen[2338]),

			.SO(gen[2431]),
			.S(gen[2432]),
			.SE(gen[2433]),

			.SELF(gen[2337]),
			.cell_state(gen[2337])
		); 

/******************* CELL 2338 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2338 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2242]),
			.N(gen[2243]),
			.NE(gen[2244]),

			.O(gen[2337]),
			.E(gen[2339]),

			.SO(gen[2432]),
			.S(gen[2433]),
			.SE(gen[2434]),

			.SELF(gen[2338]),
			.cell_state(gen[2338])
		); 

/******************* CELL 2339 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2339 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2243]),
			.N(gen[2244]),
			.NE(gen[2245]),

			.O(gen[2338]),
			.E(gen[2340]),

			.SO(gen[2433]),
			.S(gen[2434]),
			.SE(gen[2435]),

			.SELF(gen[2339]),
			.cell_state(gen[2339])
		); 

/******************* CELL 2340 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2340 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2244]),
			.N(gen[2245]),
			.NE(gen[2246]),

			.O(gen[2339]),
			.E(gen[2341]),

			.SO(gen[2434]),
			.S(gen[2435]),
			.SE(gen[2436]),

			.SELF(gen[2340]),
			.cell_state(gen[2340])
		); 

/******************* CELL 2341 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2341 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2245]),
			.N(gen[2246]),
			.NE(gen[2247]),

			.O(gen[2340]),
			.E(gen[2342]),

			.SO(gen[2435]),
			.S(gen[2436]),
			.SE(gen[2437]),

			.SELF(gen[2341]),
			.cell_state(gen[2341])
		); 

/******************* CELL 2342 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2342 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2246]),
			.N(gen[2247]),
			.NE(gen[2248]),

			.O(gen[2341]),
			.E(gen[2343]),

			.SO(gen[2436]),
			.S(gen[2437]),
			.SE(gen[2438]),

			.SELF(gen[2342]),
			.cell_state(gen[2342])
		); 

/******************* CELL 2343 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2343 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2247]),
			.N(gen[2248]),
			.NE(gen[2249]),

			.O(gen[2342]),
			.E(gen[2344]),

			.SO(gen[2437]),
			.S(gen[2438]),
			.SE(gen[2439]),

			.SELF(gen[2343]),
			.cell_state(gen[2343])
		); 

/******************* CELL 2344 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2344 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2248]),
			.N(gen[2249]),
			.NE(gen[2250]),

			.O(gen[2343]),
			.E(gen[2345]),

			.SO(gen[2438]),
			.S(gen[2439]),
			.SE(gen[2440]),

			.SELF(gen[2344]),
			.cell_state(gen[2344])
		); 

/******************* CELL 2345 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2345 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2249]),
			.N(gen[2250]),
			.NE(gen[2251]),

			.O(gen[2344]),
			.E(gen[2346]),

			.SO(gen[2439]),
			.S(gen[2440]),
			.SE(gen[2441]),

			.SELF(gen[2345]),
			.cell_state(gen[2345])
		); 

/******************* CELL 2346 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2346 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2250]),
			.N(gen[2251]),
			.NE(gen[2252]),

			.O(gen[2345]),
			.E(gen[2347]),

			.SO(gen[2440]),
			.S(gen[2441]),
			.SE(gen[2442]),

			.SELF(gen[2346]),
			.cell_state(gen[2346])
		); 

/******************* CELL 2347 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2347 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2251]),
			.N(gen[2252]),
			.NE(gen[2253]),

			.O(gen[2346]),
			.E(gen[2348]),

			.SO(gen[2441]),
			.S(gen[2442]),
			.SE(gen[2443]),

			.SELF(gen[2347]),
			.cell_state(gen[2347])
		); 

/******************* CELL 2348 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2348 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2252]),
			.N(gen[2253]),
			.NE(gen[2254]),

			.O(gen[2347]),
			.E(gen[2349]),

			.SO(gen[2442]),
			.S(gen[2443]),
			.SE(gen[2444]),

			.SELF(gen[2348]),
			.cell_state(gen[2348])
		); 

/******************* CELL 2349 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2349 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2253]),
			.N(gen[2254]),
			.NE(gen[2255]),

			.O(gen[2348]),
			.E(gen[2350]),

			.SO(gen[2443]),
			.S(gen[2444]),
			.SE(gen[2445]),

			.SELF(gen[2349]),
			.cell_state(gen[2349])
		); 

/******************* CELL 2350 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2350 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2254]),
			.N(gen[2255]),
			.NE(gen[2256]),

			.O(gen[2349]),
			.E(gen[2351]),

			.SO(gen[2444]),
			.S(gen[2445]),
			.SE(gen[2446]),

			.SELF(gen[2350]),
			.cell_state(gen[2350])
		); 

/******************* CELL 2351 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2351 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2255]),
			.N(gen[2256]),
			.NE(gen[2257]),

			.O(gen[2350]),
			.E(gen[2352]),

			.SO(gen[2445]),
			.S(gen[2446]),
			.SE(gen[2447]),

			.SELF(gen[2351]),
			.cell_state(gen[2351])
		); 

/******************* CELL 2352 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2352 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2256]),
			.N(gen[2257]),
			.NE(gen[2258]),

			.O(gen[2351]),
			.E(gen[2353]),

			.SO(gen[2446]),
			.S(gen[2447]),
			.SE(gen[2448]),

			.SELF(gen[2352]),
			.cell_state(gen[2352])
		); 

/******************* CELL 2353 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2353 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2257]),
			.N(gen[2258]),
			.NE(gen[2259]),

			.O(gen[2352]),
			.E(gen[2354]),

			.SO(gen[2447]),
			.S(gen[2448]),
			.SE(gen[2449]),

			.SELF(gen[2353]),
			.cell_state(gen[2353])
		); 

/******************* CELL 2354 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2354 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2258]),
			.N(gen[2259]),
			.NE(gen[2260]),

			.O(gen[2353]),
			.E(gen[2355]),

			.SO(gen[2448]),
			.S(gen[2449]),
			.SE(gen[2450]),

			.SELF(gen[2354]),
			.cell_state(gen[2354])
		); 

/******************* CELL 2355 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2355 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2259]),
			.N(gen[2260]),
			.NE(gen[2261]),

			.O(gen[2354]),
			.E(gen[2356]),

			.SO(gen[2449]),
			.S(gen[2450]),
			.SE(gen[2451]),

			.SELF(gen[2355]),
			.cell_state(gen[2355])
		); 

/******************* CELL 2356 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2356 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2260]),
			.N(gen[2261]),
			.NE(gen[2262]),

			.O(gen[2355]),
			.E(gen[2357]),

			.SO(gen[2450]),
			.S(gen[2451]),
			.SE(gen[2452]),

			.SELF(gen[2356]),
			.cell_state(gen[2356])
		); 

/******************* CELL 2357 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2357 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2261]),
			.N(gen[2262]),
			.NE(gen[2263]),

			.O(gen[2356]),
			.E(gen[2358]),

			.SO(gen[2451]),
			.S(gen[2452]),
			.SE(gen[2453]),

			.SELF(gen[2357]),
			.cell_state(gen[2357])
		); 

/******************* CELL 2358 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2358 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2262]),
			.N(gen[2263]),
			.NE(gen[2264]),

			.O(gen[2357]),
			.E(gen[2359]),

			.SO(gen[2452]),
			.S(gen[2453]),
			.SE(gen[2454]),

			.SELF(gen[2358]),
			.cell_state(gen[2358])
		); 

/******************* CELL 2359 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2359 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2263]),
			.N(gen[2264]),
			.NE(gen[2265]),

			.O(gen[2358]),
			.E(gen[2360]),

			.SO(gen[2453]),
			.S(gen[2454]),
			.SE(gen[2455]),

			.SELF(gen[2359]),
			.cell_state(gen[2359])
		); 

/******************* CELL 2360 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2360 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2264]),
			.N(gen[2265]),
			.NE(gen[2266]),

			.O(gen[2359]),
			.E(gen[2361]),

			.SO(gen[2454]),
			.S(gen[2455]),
			.SE(gen[2456]),

			.SELF(gen[2360]),
			.cell_state(gen[2360])
		); 

/******************* CELL 2361 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2361 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2265]),
			.N(gen[2266]),
			.NE(gen[2267]),

			.O(gen[2360]),
			.E(gen[2362]),

			.SO(gen[2455]),
			.S(gen[2456]),
			.SE(gen[2457]),

			.SELF(gen[2361]),
			.cell_state(gen[2361])
		); 

/******************* CELL 2362 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2362 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2266]),
			.N(gen[2267]),
			.NE(gen[2268]),

			.O(gen[2361]),
			.E(gen[2363]),

			.SO(gen[2456]),
			.S(gen[2457]),
			.SE(gen[2458]),

			.SELF(gen[2362]),
			.cell_state(gen[2362])
		); 

/******************* CELL 2363 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2363 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2267]),
			.N(gen[2268]),
			.NE(gen[2269]),

			.O(gen[2362]),
			.E(gen[2364]),

			.SO(gen[2457]),
			.S(gen[2458]),
			.SE(gen[2459]),

			.SELF(gen[2363]),
			.cell_state(gen[2363])
		); 

/******************* CELL 2364 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2364 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2268]),
			.N(gen[2269]),
			.NE(gen[2270]),

			.O(gen[2363]),
			.E(gen[2365]),

			.SO(gen[2458]),
			.S(gen[2459]),
			.SE(gen[2460]),

			.SELF(gen[2364]),
			.cell_state(gen[2364])
		); 

/******************* CELL 2365 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2365 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2269]),
			.N(gen[2270]),
			.NE(gen[2271]),

			.O(gen[2364]),
			.E(gen[2366]),

			.SO(gen[2459]),
			.S(gen[2460]),
			.SE(gen[2461]),

			.SELF(gen[2365]),
			.cell_state(gen[2365])
		); 

/******************* CELL 2366 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2366 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2270]),
			.N(gen[2271]),
			.NE(gen[2272]),

			.O(gen[2365]),
			.E(gen[2367]),

			.SO(gen[2460]),
			.S(gen[2461]),
			.SE(gen[2462]),

			.SELF(gen[2366]),
			.cell_state(gen[2366])
		); 

/******************* CELL 2367 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2367 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2271]),
			.N(gen[2272]),
			.NE(gen[2273]),

			.O(gen[2366]),
			.E(gen[2368]),

			.SO(gen[2461]),
			.S(gen[2462]),
			.SE(gen[2463]),

			.SELF(gen[2367]),
			.cell_state(gen[2367])
		); 

/******************* CELL 2368 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2368 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2272]),
			.N(gen[2273]),
			.NE(gen[2274]),

			.O(gen[2367]),
			.E(gen[2369]),

			.SO(gen[2462]),
			.S(gen[2463]),
			.SE(gen[2464]),

			.SELF(gen[2368]),
			.cell_state(gen[2368])
		); 

/******************* CELL 2369 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2369 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2273]),
			.N(gen[2274]),
			.NE(gen[2275]),

			.O(gen[2368]),
			.E(gen[2370]),

			.SO(gen[2463]),
			.S(gen[2464]),
			.SE(gen[2465]),

			.SELF(gen[2369]),
			.cell_state(gen[2369])
		); 

/******************* CELL 2370 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2370 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2274]),
			.N(gen[2275]),
			.NE(gen[2276]),

			.O(gen[2369]),
			.E(gen[2371]),

			.SO(gen[2464]),
			.S(gen[2465]),
			.SE(gen[2466]),

			.SELF(gen[2370]),
			.cell_state(gen[2370])
		); 

/******************* CELL 2371 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2371 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2275]),
			.N(gen[2276]),
			.NE(gen[2277]),

			.O(gen[2370]),
			.E(gen[2372]),

			.SO(gen[2465]),
			.S(gen[2466]),
			.SE(gen[2467]),

			.SELF(gen[2371]),
			.cell_state(gen[2371])
		); 

/******************* CELL 2372 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2372 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2276]),
			.N(gen[2277]),
			.NE(gen[2278]),

			.O(gen[2371]),
			.E(gen[2373]),

			.SO(gen[2466]),
			.S(gen[2467]),
			.SE(gen[2468]),

			.SELF(gen[2372]),
			.cell_state(gen[2372])
		); 

/******************* CELL 2373 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2373 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2277]),
			.N(gen[2278]),
			.NE(gen[2279]),

			.O(gen[2372]),
			.E(gen[2374]),

			.SO(gen[2467]),
			.S(gen[2468]),
			.SE(gen[2469]),

			.SELF(gen[2373]),
			.cell_state(gen[2373])
		); 

/******************* CELL 2374 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2374 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2278]),
			.N(gen[2279]),
			.NE(gen[2278]),

			.O(gen[2373]),
			.E(gen[2373]),

			.SO(gen[2468]),
			.S(gen[2469]),
			.SE(gen[2468]),

			.SELF(gen[2374]),
			.cell_state(gen[2374])
		); 

/******************* CELL 2375 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2375 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2281]),
			.N(gen[2280]),
			.NE(gen[2281]),

			.O(gen[2376]),
			.E(gen[2376]),

			.SO(gen[2471]),
			.S(gen[2470]),
			.SE(gen[2471]),

			.SELF(gen[2375]),
			.cell_state(gen[2375])
		); 

/******************* CELL 2376 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2376 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2280]),
			.N(gen[2281]),
			.NE(gen[2282]),

			.O(gen[2375]),
			.E(gen[2377]),

			.SO(gen[2470]),
			.S(gen[2471]),
			.SE(gen[2472]),

			.SELF(gen[2376]),
			.cell_state(gen[2376])
		); 

/******************* CELL 2377 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2377 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2281]),
			.N(gen[2282]),
			.NE(gen[2283]),

			.O(gen[2376]),
			.E(gen[2378]),

			.SO(gen[2471]),
			.S(gen[2472]),
			.SE(gen[2473]),

			.SELF(gen[2377]),
			.cell_state(gen[2377])
		); 

/******************* CELL 2378 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2378 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2282]),
			.N(gen[2283]),
			.NE(gen[2284]),

			.O(gen[2377]),
			.E(gen[2379]),

			.SO(gen[2472]),
			.S(gen[2473]),
			.SE(gen[2474]),

			.SELF(gen[2378]),
			.cell_state(gen[2378])
		); 

/******************* CELL 2379 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2379 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2283]),
			.N(gen[2284]),
			.NE(gen[2285]),

			.O(gen[2378]),
			.E(gen[2380]),

			.SO(gen[2473]),
			.S(gen[2474]),
			.SE(gen[2475]),

			.SELF(gen[2379]),
			.cell_state(gen[2379])
		); 

/******************* CELL 2380 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2380 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2284]),
			.N(gen[2285]),
			.NE(gen[2286]),

			.O(gen[2379]),
			.E(gen[2381]),

			.SO(gen[2474]),
			.S(gen[2475]),
			.SE(gen[2476]),

			.SELF(gen[2380]),
			.cell_state(gen[2380])
		); 

/******************* CELL 2381 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2381 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2285]),
			.N(gen[2286]),
			.NE(gen[2287]),

			.O(gen[2380]),
			.E(gen[2382]),

			.SO(gen[2475]),
			.S(gen[2476]),
			.SE(gen[2477]),

			.SELF(gen[2381]),
			.cell_state(gen[2381])
		); 

/******************* CELL 2382 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2382 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2286]),
			.N(gen[2287]),
			.NE(gen[2288]),

			.O(gen[2381]),
			.E(gen[2383]),

			.SO(gen[2476]),
			.S(gen[2477]),
			.SE(gen[2478]),

			.SELF(gen[2382]),
			.cell_state(gen[2382])
		); 

/******************* CELL 2383 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2383 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2287]),
			.N(gen[2288]),
			.NE(gen[2289]),

			.O(gen[2382]),
			.E(gen[2384]),

			.SO(gen[2477]),
			.S(gen[2478]),
			.SE(gen[2479]),

			.SELF(gen[2383]),
			.cell_state(gen[2383])
		); 

/******************* CELL 2384 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2384 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2288]),
			.N(gen[2289]),
			.NE(gen[2290]),

			.O(gen[2383]),
			.E(gen[2385]),

			.SO(gen[2478]),
			.S(gen[2479]),
			.SE(gen[2480]),

			.SELF(gen[2384]),
			.cell_state(gen[2384])
		); 

/******************* CELL 2385 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2385 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2289]),
			.N(gen[2290]),
			.NE(gen[2291]),

			.O(gen[2384]),
			.E(gen[2386]),

			.SO(gen[2479]),
			.S(gen[2480]),
			.SE(gen[2481]),

			.SELF(gen[2385]),
			.cell_state(gen[2385])
		); 

/******************* CELL 2386 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2386 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2290]),
			.N(gen[2291]),
			.NE(gen[2292]),

			.O(gen[2385]),
			.E(gen[2387]),

			.SO(gen[2480]),
			.S(gen[2481]),
			.SE(gen[2482]),

			.SELF(gen[2386]),
			.cell_state(gen[2386])
		); 

/******************* CELL 2387 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2387 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2291]),
			.N(gen[2292]),
			.NE(gen[2293]),

			.O(gen[2386]),
			.E(gen[2388]),

			.SO(gen[2481]),
			.S(gen[2482]),
			.SE(gen[2483]),

			.SELF(gen[2387]),
			.cell_state(gen[2387])
		); 

/******************* CELL 2388 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2388 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2292]),
			.N(gen[2293]),
			.NE(gen[2294]),

			.O(gen[2387]),
			.E(gen[2389]),

			.SO(gen[2482]),
			.S(gen[2483]),
			.SE(gen[2484]),

			.SELF(gen[2388]),
			.cell_state(gen[2388])
		); 

/******************* CELL 2389 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2389 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2293]),
			.N(gen[2294]),
			.NE(gen[2295]),

			.O(gen[2388]),
			.E(gen[2390]),

			.SO(gen[2483]),
			.S(gen[2484]),
			.SE(gen[2485]),

			.SELF(gen[2389]),
			.cell_state(gen[2389])
		); 

/******************* CELL 2390 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2390 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2294]),
			.N(gen[2295]),
			.NE(gen[2296]),

			.O(gen[2389]),
			.E(gen[2391]),

			.SO(gen[2484]),
			.S(gen[2485]),
			.SE(gen[2486]),

			.SELF(gen[2390]),
			.cell_state(gen[2390])
		); 

/******************* CELL 2391 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2391 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2295]),
			.N(gen[2296]),
			.NE(gen[2297]),

			.O(gen[2390]),
			.E(gen[2392]),

			.SO(gen[2485]),
			.S(gen[2486]),
			.SE(gen[2487]),

			.SELF(gen[2391]),
			.cell_state(gen[2391])
		); 

/******************* CELL 2392 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2392 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2296]),
			.N(gen[2297]),
			.NE(gen[2298]),

			.O(gen[2391]),
			.E(gen[2393]),

			.SO(gen[2486]),
			.S(gen[2487]),
			.SE(gen[2488]),

			.SELF(gen[2392]),
			.cell_state(gen[2392])
		); 

/******************* CELL 2393 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2393 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2297]),
			.N(gen[2298]),
			.NE(gen[2299]),

			.O(gen[2392]),
			.E(gen[2394]),

			.SO(gen[2487]),
			.S(gen[2488]),
			.SE(gen[2489]),

			.SELF(gen[2393]),
			.cell_state(gen[2393])
		); 

/******************* CELL 2394 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2394 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2298]),
			.N(gen[2299]),
			.NE(gen[2300]),

			.O(gen[2393]),
			.E(gen[2395]),

			.SO(gen[2488]),
			.S(gen[2489]),
			.SE(gen[2490]),

			.SELF(gen[2394]),
			.cell_state(gen[2394])
		); 

/******************* CELL 2395 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2395 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2299]),
			.N(gen[2300]),
			.NE(gen[2301]),

			.O(gen[2394]),
			.E(gen[2396]),

			.SO(gen[2489]),
			.S(gen[2490]),
			.SE(gen[2491]),

			.SELF(gen[2395]),
			.cell_state(gen[2395])
		); 

/******************* CELL 2396 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2396 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2300]),
			.N(gen[2301]),
			.NE(gen[2302]),

			.O(gen[2395]),
			.E(gen[2397]),

			.SO(gen[2490]),
			.S(gen[2491]),
			.SE(gen[2492]),

			.SELF(gen[2396]),
			.cell_state(gen[2396])
		); 

/******************* CELL 2397 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2397 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2301]),
			.N(gen[2302]),
			.NE(gen[2303]),

			.O(gen[2396]),
			.E(gen[2398]),

			.SO(gen[2491]),
			.S(gen[2492]),
			.SE(gen[2493]),

			.SELF(gen[2397]),
			.cell_state(gen[2397])
		); 

/******************* CELL 2398 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2398 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2302]),
			.N(gen[2303]),
			.NE(gen[2304]),

			.O(gen[2397]),
			.E(gen[2399]),

			.SO(gen[2492]),
			.S(gen[2493]),
			.SE(gen[2494]),

			.SELF(gen[2398]),
			.cell_state(gen[2398])
		); 

/******************* CELL 2399 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2399 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2303]),
			.N(gen[2304]),
			.NE(gen[2305]),

			.O(gen[2398]),
			.E(gen[2400]),

			.SO(gen[2493]),
			.S(gen[2494]),
			.SE(gen[2495]),

			.SELF(gen[2399]),
			.cell_state(gen[2399])
		); 

/******************* CELL 2400 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2400 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2304]),
			.N(gen[2305]),
			.NE(gen[2306]),

			.O(gen[2399]),
			.E(gen[2401]),

			.SO(gen[2494]),
			.S(gen[2495]),
			.SE(gen[2496]),

			.SELF(gen[2400]),
			.cell_state(gen[2400])
		); 

/******************* CELL 2401 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2401 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2305]),
			.N(gen[2306]),
			.NE(gen[2307]),

			.O(gen[2400]),
			.E(gen[2402]),

			.SO(gen[2495]),
			.S(gen[2496]),
			.SE(gen[2497]),

			.SELF(gen[2401]),
			.cell_state(gen[2401])
		); 

/******************* CELL 2402 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2402 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2306]),
			.N(gen[2307]),
			.NE(gen[2308]),

			.O(gen[2401]),
			.E(gen[2403]),

			.SO(gen[2496]),
			.S(gen[2497]),
			.SE(gen[2498]),

			.SELF(gen[2402]),
			.cell_state(gen[2402])
		); 

/******************* CELL 2403 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2403 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2307]),
			.N(gen[2308]),
			.NE(gen[2309]),

			.O(gen[2402]),
			.E(gen[2404]),

			.SO(gen[2497]),
			.S(gen[2498]),
			.SE(gen[2499]),

			.SELF(gen[2403]),
			.cell_state(gen[2403])
		); 

/******************* CELL 2404 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2404 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2308]),
			.N(gen[2309]),
			.NE(gen[2310]),

			.O(gen[2403]),
			.E(gen[2405]),

			.SO(gen[2498]),
			.S(gen[2499]),
			.SE(gen[2500]),

			.SELF(gen[2404]),
			.cell_state(gen[2404])
		); 

/******************* CELL 2405 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2405 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2309]),
			.N(gen[2310]),
			.NE(gen[2311]),

			.O(gen[2404]),
			.E(gen[2406]),

			.SO(gen[2499]),
			.S(gen[2500]),
			.SE(gen[2501]),

			.SELF(gen[2405]),
			.cell_state(gen[2405])
		); 

/******************* CELL 2406 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2406 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2310]),
			.N(gen[2311]),
			.NE(gen[2312]),

			.O(gen[2405]),
			.E(gen[2407]),

			.SO(gen[2500]),
			.S(gen[2501]),
			.SE(gen[2502]),

			.SELF(gen[2406]),
			.cell_state(gen[2406])
		); 

/******************* CELL 2407 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2407 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2311]),
			.N(gen[2312]),
			.NE(gen[2313]),

			.O(gen[2406]),
			.E(gen[2408]),

			.SO(gen[2501]),
			.S(gen[2502]),
			.SE(gen[2503]),

			.SELF(gen[2407]),
			.cell_state(gen[2407])
		); 

/******************* CELL 2408 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2408 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2312]),
			.N(gen[2313]),
			.NE(gen[2314]),

			.O(gen[2407]),
			.E(gen[2409]),

			.SO(gen[2502]),
			.S(gen[2503]),
			.SE(gen[2504]),

			.SELF(gen[2408]),
			.cell_state(gen[2408])
		); 

/******************* CELL 2409 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2409 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2313]),
			.N(gen[2314]),
			.NE(gen[2315]),

			.O(gen[2408]),
			.E(gen[2410]),

			.SO(gen[2503]),
			.S(gen[2504]),
			.SE(gen[2505]),

			.SELF(gen[2409]),
			.cell_state(gen[2409])
		); 

/******************* CELL 2410 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2410 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2314]),
			.N(gen[2315]),
			.NE(gen[2316]),

			.O(gen[2409]),
			.E(gen[2411]),

			.SO(gen[2504]),
			.S(gen[2505]),
			.SE(gen[2506]),

			.SELF(gen[2410]),
			.cell_state(gen[2410])
		); 

/******************* CELL 2411 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2411 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2315]),
			.N(gen[2316]),
			.NE(gen[2317]),

			.O(gen[2410]),
			.E(gen[2412]),

			.SO(gen[2505]),
			.S(gen[2506]),
			.SE(gen[2507]),

			.SELF(gen[2411]),
			.cell_state(gen[2411])
		); 

/******************* CELL 2412 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2412 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2316]),
			.N(gen[2317]),
			.NE(gen[2318]),

			.O(gen[2411]),
			.E(gen[2413]),

			.SO(gen[2506]),
			.S(gen[2507]),
			.SE(gen[2508]),

			.SELF(gen[2412]),
			.cell_state(gen[2412])
		); 

/******************* CELL 2413 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2413 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2317]),
			.N(gen[2318]),
			.NE(gen[2319]),

			.O(gen[2412]),
			.E(gen[2414]),

			.SO(gen[2507]),
			.S(gen[2508]),
			.SE(gen[2509]),

			.SELF(gen[2413]),
			.cell_state(gen[2413])
		); 

/******************* CELL 2414 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2414 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2318]),
			.N(gen[2319]),
			.NE(gen[2320]),

			.O(gen[2413]),
			.E(gen[2415]),

			.SO(gen[2508]),
			.S(gen[2509]),
			.SE(gen[2510]),

			.SELF(gen[2414]),
			.cell_state(gen[2414])
		); 

/******************* CELL 2415 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2415 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2319]),
			.N(gen[2320]),
			.NE(gen[2321]),

			.O(gen[2414]),
			.E(gen[2416]),

			.SO(gen[2509]),
			.S(gen[2510]),
			.SE(gen[2511]),

			.SELF(gen[2415]),
			.cell_state(gen[2415])
		); 

/******************* CELL 2416 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2416 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2320]),
			.N(gen[2321]),
			.NE(gen[2322]),

			.O(gen[2415]),
			.E(gen[2417]),

			.SO(gen[2510]),
			.S(gen[2511]),
			.SE(gen[2512]),

			.SELF(gen[2416]),
			.cell_state(gen[2416])
		); 

/******************* CELL 2417 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2417 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2321]),
			.N(gen[2322]),
			.NE(gen[2323]),

			.O(gen[2416]),
			.E(gen[2418]),

			.SO(gen[2511]),
			.S(gen[2512]),
			.SE(gen[2513]),

			.SELF(gen[2417]),
			.cell_state(gen[2417])
		); 

/******************* CELL 2418 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2418 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2322]),
			.N(gen[2323]),
			.NE(gen[2324]),

			.O(gen[2417]),
			.E(gen[2419]),

			.SO(gen[2512]),
			.S(gen[2513]),
			.SE(gen[2514]),

			.SELF(gen[2418]),
			.cell_state(gen[2418])
		); 

/******************* CELL 2419 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2419 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2323]),
			.N(gen[2324]),
			.NE(gen[2325]),

			.O(gen[2418]),
			.E(gen[2420]),

			.SO(gen[2513]),
			.S(gen[2514]),
			.SE(gen[2515]),

			.SELF(gen[2419]),
			.cell_state(gen[2419])
		); 

/******************* CELL 2420 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2420 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2324]),
			.N(gen[2325]),
			.NE(gen[2326]),

			.O(gen[2419]),
			.E(gen[2421]),

			.SO(gen[2514]),
			.S(gen[2515]),
			.SE(gen[2516]),

			.SELF(gen[2420]),
			.cell_state(gen[2420])
		); 

/******************* CELL 2421 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2421 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2325]),
			.N(gen[2326]),
			.NE(gen[2327]),

			.O(gen[2420]),
			.E(gen[2422]),

			.SO(gen[2515]),
			.S(gen[2516]),
			.SE(gen[2517]),

			.SELF(gen[2421]),
			.cell_state(gen[2421])
		); 

/******************* CELL 2422 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2422 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2326]),
			.N(gen[2327]),
			.NE(gen[2328]),

			.O(gen[2421]),
			.E(gen[2423]),

			.SO(gen[2516]),
			.S(gen[2517]),
			.SE(gen[2518]),

			.SELF(gen[2422]),
			.cell_state(gen[2422])
		); 

/******************* CELL 2423 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2423 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2327]),
			.N(gen[2328]),
			.NE(gen[2329]),

			.O(gen[2422]),
			.E(gen[2424]),

			.SO(gen[2517]),
			.S(gen[2518]),
			.SE(gen[2519]),

			.SELF(gen[2423]),
			.cell_state(gen[2423])
		); 

/******************* CELL 2424 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2424 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2328]),
			.N(gen[2329]),
			.NE(gen[2330]),

			.O(gen[2423]),
			.E(gen[2425]),

			.SO(gen[2518]),
			.S(gen[2519]),
			.SE(gen[2520]),

			.SELF(gen[2424]),
			.cell_state(gen[2424])
		); 

/******************* CELL 2425 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2425 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2329]),
			.N(gen[2330]),
			.NE(gen[2331]),

			.O(gen[2424]),
			.E(gen[2426]),

			.SO(gen[2519]),
			.S(gen[2520]),
			.SE(gen[2521]),

			.SELF(gen[2425]),
			.cell_state(gen[2425])
		); 

/******************* CELL 2426 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2426 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2330]),
			.N(gen[2331]),
			.NE(gen[2332]),

			.O(gen[2425]),
			.E(gen[2427]),

			.SO(gen[2520]),
			.S(gen[2521]),
			.SE(gen[2522]),

			.SELF(gen[2426]),
			.cell_state(gen[2426])
		); 

/******************* CELL 2427 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2427 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2331]),
			.N(gen[2332]),
			.NE(gen[2333]),

			.O(gen[2426]),
			.E(gen[2428]),

			.SO(gen[2521]),
			.S(gen[2522]),
			.SE(gen[2523]),

			.SELF(gen[2427]),
			.cell_state(gen[2427])
		); 

/******************* CELL 2428 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2428 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2332]),
			.N(gen[2333]),
			.NE(gen[2334]),

			.O(gen[2427]),
			.E(gen[2429]),

			.SO(gen[2522]),
			.S(gen[2523]),
			.SE(gen[2524]),

			.SELF(gen[2428]),
			.cell_state(gen[2428])
		); 

/******************* CELL 2429 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2429 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2333]),
			.N(gen[2334]),
			.NE(gen[2335]),

			.O(gen[2428]),
			.E(gen[2430]),

			.SO(gen[2523]),
			.S(gen[2524]),
			.SE(gen[2525]),

			.SELF(gen[2429]),
			.cell_state(gen[2429])
		); 

/******************* CELL 2430 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2430 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2334]),
			.N(gen[2335]),
			.NE(gen[2336]),

			.O(gen[2429]),
			.E(gen[2431]),

			.SO(gen[2524]),
			.S(gen[2525]),
			.SE(gen[2526]),

			.SELF(gen[2430]),
			.cell_state(gen[2430])
		); 

/******************* CELL 2431 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2431 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2335]),
			.N(gen[2336]),
			.NE(gen[2337]),

			.O(gen[2430]),
			.E(gen[2432]),

			.SO(gen[2525]),
			.S(gen[2526]),
			.SE(gen[2527]),

			.SELF(gen[2431]),
			.cell_state(gen[2431])
		); 

/******************* CELL 2432 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2432 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2336]),
			.N(gen[2337]),
			.NE(gen[2338]),

			.O(gen[2431]),
			.E(gen[2433]),

			.SO(gen[2526]),
			.S(gen[2527]),
			.SE(gen[2528]),

			.SELF(gen[2432]),
			.cell_state(gen[2432])
		); 

/******************* CELL 2433 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2433 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2337]),
			.N(gen[2338]),
			.NE(gen[2339]),

			.O(gen[2432]),
			.E(gen[2434]),

			.SO(gen[2527]),
			.S(gen[2528]),
			.SE(gen[2529]),

			.SELF(gen[2433]),
			.cell_state(gen[2433])
		); 

/******************* CELL 2434 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2434 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2338]),
			.N(gen[2339]),
			.NE(gen[2340]),

			.O(gen[2433]),
			.E(gen[2435]),

			.SO(gen[2528]),
			.S(gen[2529]),
			.SE(gen[2530]),

			.SELF(gen[2434]),
			.cell_state(gen[2434])
		); 

/******************* CELL 2435 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2435 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2339]),
			.N(gen[2340]),
			.NE(gen[2341]),

			.O(gen[2434]),
			.E(gen[2436]),

			.SO(gen[2529]),
			.S(gen[2530]),
			.SE(gen[2531]),

			.SELF(gen[2435]),
			.cell_state(gen[2435])
		); 

/******************* CELL 2436 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2436 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2340]),
			.N(gen[2341]),
			.NE(gen[2342]),

			.O(gen[2435]),
			.E(gen[2437]),

			.SO(gen[2530]),
			.S(gen[2531]),
			.SE(gen[2532]),

			.SELF(gen[2436]),
			.cell_state(gen[2436])
		); 

/******************* CELL 2437 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2437 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2341]),
			.N(gen[2342]),
			.NE(gen[2343]),

			.O(gen[2436]),
			.E(gen[2438]),

			.SO(gen[2531]),
			.S(gen[2532]),
			.SE(gen[2533]),

			.SELF(gen[2437]),
			.cell_state(gen[2437])
		); 

/******************* CELL 2438 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2438 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2342]),
			.N(gen[2343]),
			.NE(gen[2344]),

			.O(gen[2437]),
			.E(gen[2439]),

			.SO(gen[2532]),
			.S(gen[2533]),
			.SE(gen[2534]),

			.SELF(gen[2438]),
			.cell_state(gen[2438])
		); 

/******************* CELL 2439 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2439 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2343]),
			.N(gen[2344]),
			.NE(gen[2345]),

			.O(gen[2438]),
			.E(gen[2440]),

			.SO(gen[2533]),
			.S(gen[2534]),
			.SE(gen[2535]),

			.SELF(gen[2439]),
			.cell_state(gen[2439])
		); 

/******************* CELL 2440 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2440 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2344]),
			.N(gen[2345]),
			.NE(gen[2346]),

			.O(gen[2439]),
			.E(gen[2441]),

			.SO(gen[2534]),
			.S(gen[2535]),
			.SE(gen[2536]),

			.SELF(gen[2440]),
			.cell_state(gen[2440])
		); 

/******************* CELL 2441 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2441 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2345]),
			.N(gen[2346]),
			.NE(gen[2347]),

			.O(gen[2440]),
			.E(gen[2442]),

			.SO(gen[2535]),
			.S(gen[2536]),
			.SE(gen[2537]),

			.SELF(gen[2441]),
			.cell_state(gen[2441])
		); 

/******************* CELL 2442 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2442 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2346]),
			.N(gen[2347]),
			.NE(gen[2348]),

			.O(gen[2441]),
			.E(gen[2443]),

			.SO(gen[2536]),
			.S(gen[2537]),
			.SE(gen[2538]),

			.SELF(gen[2442]),
			.cell_state(gen[2442])
		); 

/******************* CELL 2443 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2443 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2347]),
			.N(gen[2348]),
			.NE(gen[2349]),

			.O(gen[2442]),
			.E(gen[2444]),

			.SO(gen[2537]),
			.S(gen[2538]),
			.SE(gen[2539]),

			.SELF(gen[2443]),
			.cell_state(gen[2443])
		); 

/******************* CELL 2444 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2444 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2348]),
			.N(gen[2349]),
			.NE(gen[2350]),

			.O(gen[2443]),
			.E(gen[2445]),

			.SO(gen[2538]),
			.S(gen[2539]),
			.SE(gen[2540]),

			.SELF(gen[2444]),
			.cell_state(gen[2444])
		); 

/******************* CELL 2445 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2445 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2349]),
			.N(gen[2350]),
			.NE(gen[2351]),

			.O(gen[2444]),
			.E(gen[2446]),

			.SO(gen[2539]),
			.S(gen[2540]),
			.SE(gen[2541]),

			.SELF(gen[2445]),
			.cell_state(gen[2445])
		); 

/******************* CELL 2446 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2446 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2350]),
			.N(gen[2351]),
			.NE(gen[2352]),

			.O(gen[2445]),
			.E(gen[2447]),

			.SO(gen[2540]),
			.S(gen[2541]),
			.SE(gen[2542]),

			.SELF(gen[2446]),
			.cell_state(gen[2446])
		); 

/******************* CELL 2447 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2447 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2351]),
			.N(gen[2352]),
			.NE(gen[2353]),

			.O(gen[2446]),
			.E(gen[2448]),

			.SO(gen[2541]),
			.S(gen[2542]),
			.SE(gen[2543]),

			.SELF(gen[2447]),
			.cell_state(gen[2447])
		); 

/******************* CELL 2448 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2448 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2352]),
			.N(gen[2353]),
			.NE(gen[2354]),

			.O(gen[2447]),
			.E(gen[2449]),

			.SO(gen[2542]),
			.S(gen[2543]),
			.SE(gen[2544]),

			.SELF(gen[2448]),
			.cell_state(gen[2448])
		); 

/******************* CELL 2449 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2449 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2353]),
			.N(gen[2354]),
			.NE(gen[2355]),

			.O(gen[2448]),
			.E(gen[2450]),

			.SO(gen[2543]),
			.S(gen[2544]),
			.SE(gen[2545]),

			.SELF(gen[2449]),
			.cell_state(gen[2449])
		); 

/******************* CELL 2450 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2450 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2354]),
			.N(gen[2355]),
			.NE(gen[2356]),

			.O(gen[2449]),
			.E(gen[2451]),

			.SO(gen[2544]),
			.S(gen[2545]),
			.SE(gen[2546]),

			.SELF(gen[2450]),
			.cell_state(gen[2450])
		); 

/******************* CELL 2451 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2451 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2355]),
			.N(gen[2356]),
			.NE(gen[2357]),

			.O(gen[2450]),
			.E(gen[2452]),

			.SO(gen[2545]),
			.S(gen[2546]),
			.SE(gen[2547]),

			.SELF(gen[2451]),
			.cell_state(gen[2451])
		); 

/******************* CELL 2452 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2452 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2356]),
			.N(gen[2357]),
			.NE(gen[2358]),

			.O(gen[2451]),
			.E(gen[2453]),

			.SO(gen[2546]),
			.S(gen[2547]),
			.SE(gen[2548]),

			.SELF(gen[2452]),
			.cell_state(gen[2452])
		); 

/******************* CELL 2453 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2453 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2357]),
			.N(gen[2358]),
			.NE(gen[2359]),

			.O(gen[2452]),
			.E(gen[2454]),

			.SO(gen[2547]),
			.S(gen[2548]),
			.SE(gen[2549]),

			.SELF(gen[2453]),
			.cell_state(gen[2453])
		); 

/******************* CELL 2454 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2454 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2358]),
			.N(gen[2359]),
			.NE(gen[2360]),

			.O(gen[2453]),
			.E(gen[2455]),

			.SO(gen[2548]),
			.S(gen[2549]),
			.SE(gen[2550]),

			.SELF(gen[2454]),
			.cell_state(gen[2454])
		); 

/******************* CELL 2455 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2455 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2359]),
			.N(gen[2360]),
			.NE(gen[2361]),

			.O(gen[2454]),
			.E(gen[2456]),

			.SO(gen[2549]),
			.S(gen[2550]),
			.SE(gen[2551]),

			.SELF(gen[2455]),
			.cell_state(gen[2455])
		); 

/******************* CELL 2456 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2456 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2360]),
			.N(gen[2361]),
			.NE(gen[2362]),

			.O(gen[2455]),
			.E(gen[2457]),

			.SO(gen[2550]),
			.S(gen[2551]),
			.SE(gen[2552]),

			.SELF(gen[2456]),
			.cell_state(gen[2456])
		); 

/******************* CELL 2457 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2457 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2361]),
			.N(gen[2362]),
			.NE(gen[2363]),

			.O(gen[2456]),
			.E(gen[2458]),

			.SO(gen[2551]),
			.S(gen[2552]),
			.SE(gen[2553]),

			.SELF(gen[2457]),
			.cell_state(gen[2457])
		); 

/******************* CELL 2458 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2458 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2362]),
			.N(gen[2363]),
			.NE(gen[2364]),

			.O(gen[2457]),
			.E(gen[2459]),

			.SO(gen[2552]),
			.S(gen[2553]),
			.SE(gen[2554]),

			.SELF(gen[2458]),
			.cell_state(gen[2458])
		); 

/******************* CELL 2459 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2459 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2363]),
			.N(gen[2364]),
			.NE(gen[2365]),

			.O(gen[2458]),
			.E(gen[2460]),

			.SO(gen[2553]),
			.S(gen[2554]),
			.SE(gen[2555]),

			.SELF(gen[2459]),
			.cell_state(gen[2459])
		); 

/******************* CELL 2460 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2460 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2364]),
			.N(gen[2365]),
			.NE(gen[2366]),

			.O(gen[2459]),
			.E(gen[2461]),

			.SO(gen[2554]),
			.S(gen[2555]),
			.SE(gen[2556]),

			.SELF(gen[2460]),
			.cell_state(gen[2460])
		); 

/******************* CELL 2461 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2461 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2365]),
			.N(gen[2366]),
			.NE(gen[2367]),

			.O(gen[2460]),
			.E(gen[2462]),

			.SO(gen[2555]),
			.S(gen[2556]),
			.SE(gen[2557]),

			.SELF(gen[2461]),
			.cell_state(gen[2461])
		); 

/******************* CELL 2462 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2462 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2366]),
			.N(gen[2367]),
			.NE(gen[2368]),

			.O(gen[2461]),
			.E(gen[2463]),

			.SO(gen[2556]),
			.S(gen[2557]),
			.SE(gen[2558]),

			.SELF(gen[2462]),
			.cell_state(gen[2462])
		); 

/******************* CELL 2463 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2463 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2367]),
			.N(gen[2368]),
			.NE(gen[2369]),

			.O(gen[2462]),
			.E(gen[2464]),

			.SO(gen[2557]),
			.S(gen[2558]),
			.SE(gen[2559]),

			.SELF(gen[2463]),
			.cell_state(gen[2463])
		); 

/******************* CELL 2464 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2464 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2368]),
			.N(gen[2369]),
			.NE(gen[2370]),

			.O(gen[2463]),
			.E(gen[2465]),

			.SO(gen[2558]),
			.S(gen[2559]),
			.SE(gen[2560]),

			.SELF(gen[2464]),
			.cell_state(gen[2464])
		); 

/******************* CELL 2465 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2465 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2369]),
			.N(gen[2370]),
			.NE(gen[2371]),

			.O(gen[2464]),
			.E(gen[2466]),

			.SO(gen[2559]),
			.S(gen[2560]),
			.SE(gen[2561]),

			.SELF(gen[2465]),
			.cell_state(gen[2465])
		); 

/******************* CELL 2466 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2466 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2370]),
			.N(gen[2371]),
			.NE(gen[2372]),

			.O(gen[2465]),
			.E(gen[2467]),

			.SO(gen[2560]),
			.S(gen[2561]),
			.SE(gen[2562]),

			.SELF(gen[2466]),
			.cell_state(gen[2466])
		); 

/******************* CELL 2467 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2467 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2371]),
			.N(gen[2372]),
			.NE(gen[2373]),

			.O(gen[2466]),
			.E(gen[2468]),

			.SO(gen[2561]),
			.S(gen[2562]),
			.SE(gen[2563]),

			.SELF(gen[2467]),
			.cell_state(gen[2467])
		); 

/******************* CELL 2468 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2468 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2372]),
			.N(gen[2373]),
			.NE(gen[2374]),

			.O(gen[2467]),
			.E(gen[2469]),

			.SO(gen[2562]),
			.S(gen[2563]),
			.SE(gen[2564]),

			.SELF(gen[2468]),
			.cell_state(gen[2468])
		); 

/******************* CELL 2469 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2469 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2373]),
			.N(gen[2374]),
			.NE(gen[2373]),

			.O(gen[2468]),
			.E(gen[2468]),

			.SO(gen[2563]),
			.S(gen[2564]),
			.SE(gen[2563]),

			.SELF(gen[2469]),
			.cell_state(gen[2469])
		); 

/******************* CELL 2470 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2470 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2376]),
			.N(gen[2375]),
			.NE(gen[2376]),

			.O(gen[2471]),
			.E(gen[2471]),

			.SO(gen[2566]),
			.S(gen[2565]),
			.SE(gen[2566]),

			.SELF(gen[2470]),
			.cell_state(gen[2470])
		); 

/******************* CELL 2471 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2471 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2375]),
			.N(gen[2376]),
			.NE(gen[2377]),

			.O(gen[2470]),
			.E(gen[2472]),

			.SO(gen[2565]),
			.S(gen[2566]),
			.SE(gen[2567]),

			.SELF(gen[2471]),
			.cell_state(gen[2471])
		); 

/******************* CELL 2472 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2472 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2376]),
			.N(gen[2377]),
			.NE(gen[2378]),

			.O(gen[2471]),
			.E(gen[2473]),

			.SO(gen[2566]),
			.S(gen[2567]),
			.SE(gen[2568]),

			.SELF(gen[2472]),
			.cell_state(gen[2472])
		); 

/******************* CELL 2473 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2473 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2377]),
			.N(gen[2378]),
			.NE(gen[2379]),

			.O(gen[2472]),
			.E(gen[2474]),

			.SO(gen[2567]),
			.S(gen[2568]),
			.SE(gen[2569]),

			.SELF(gen[2473]),
			.cell_state(gen[2473])
		); 

/******************* CELL 2474 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2474 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2378]),
			.N(gen[2379]),
			.NE(gen[2380]),

			.O(gen[2473]),
			.E(gen[2475]),

			.SO(gen[2568]),
			.S(gen[2569]),
			.SE(gen[2570]),

			.SELF(gen[2474]),
			.cell_state(gen[2474])
		); 

/******************* CELL 2475 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2475 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2379]),
			.N(gen[2380]),
			.NE(gen[2381]),

			.O(gen[2474]),
			.E(gen[2476]),

			.SO(gen[2569]),
			.S(gen[2570]),
			.SE(gen[2571]),

			.SELF(gen[2475]),
			.cell_state(gen[2475])
		); 

/******************* CELL 2476 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2476 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2380]),
			.N(gen[2381]),
			.NE(gen[2382]),

			.O(gen[2475]),
			.E(gen[2477]),

			.SO(gen[2570]),
			.S(gen[2571]),
			.SE(gen[2572]),

			.SELF(gen[2476]),
			.cell_state(gen[2476])
		); 

/******************* CELL 2477 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2477 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2381]),
			.N(gen[2382]),
			.NE(gen[2383]),

			.O(gen[2476]),
			.E(gen[2478]),

			.SO(gen[2571]),
			.S(gen[2572]),
			.SE(gen[2573]),

			.SELF(gen[2477]),
			.cell_state(gen[2477])
		); 

/******************* CELL 2478 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2478 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2382]),
			.N(gen[2383]),
			.NE(gen[2384]),

			.O(gen[2477]),
			.E(gen[2479]),

			.SO(gen[2572]),
			.S(gen[2573]),
			.SE(gen[2574]),

			.SELF(gen[2478]),
			.cell_state(gen[2478])
		); 

/******************* CELL 2479 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2479 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2383]),
			.N(gen[2384]),
			.NE(gen[2385]),

			.O(gen[2478]),
			.E(gen[2480]),

			.SO(gen[2573]),
			.S(gen[2574]),
			.SE(gen[2575]),

			.SELF(gen[2479]),
			.cell_state(gen[2479])
		); 

/******************* CELL 2480 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2480 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2384]),
			.N(gen[2385]),
			.NE(gen[2386]),

			.O(gen[2479]),
			.E(gen[2481]),

			.SO(gen[2574]),
			.S(gen[2575]),
			.SE(gen[2576]),

			.SELF(gen[2480]),
			.cell_state(gen[2480])
		); 

/******************* CELL 2481 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2481 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2385]),
			.N(gen[2386]),
			.NE(gen[2387]),

			.O(gen[2480]),
			.E(gen[2482]),

			.SO(gen[2575]),
			.S(gen[2576]),
			.SE(gen[2577]),

			.SELF(gen[2481]),
			.cell_state(gen[2481])
		); 

/******************* CELL 2482 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2482 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2386]),
			.N(gen[2387]),
			.NE(gen[2388]),

			.O(gen[2481]),
			.E(gen[2483]),

			.SO(gen[2576]),
			.S(gen[2577]),
			.SE(gen[2578]),

			.SELF(gen[2482]),
			.cell_state(gen[2482])
		); 

/******************* CELL 2483 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2483 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2387]),
			.N(gen[2388]),
			.NE(gen[2389]),

			.O(gen[2482]),
			.E(gen[2484]),

			.SO(gen[2577]),
			.S(gen[2578]),
			.SE(gen[2579]),

			.SELF(gen[2483]),
			.cell_state(gen[2483])
		); 

/******************* CELL 2484 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2484 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2388]),
			.N(gen[2389]),
			.NE(gen[2390]),

			.O(gen[2483]),
			.E(gen[2485]),

			.SO(gen[2578]),
			.S(gen[2579]),
			.SE(gen[2580]),

			.SELF(gen[2484]),
			.cell_state(gen[2484])
		); 

/******************* CELL 2485 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2485 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2389]),
			.N(gen[2390]),
			.NE(gen[2391]),

			.O(gen[2484]),
			.E(gen[2486]),

			.SO(gen[2579]),
			.S(gen[2580]),
			.SE(gen[2581]),

			.SELF(gen[2485]),
			.cell_state(gen[2485])
		); 

/******************* CELL 2486 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2486 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2390]),
			.N(gen[2391]),
			.NE(gen[2392]),

			.O(gen[2485]),
			.E(gen[2487]),

			.SO(gen[2580]),
			.S(gen[2581]),
			.SE(gen[2582]),

			.SELF(gen[2486]),
			.cell_state(gen[2486])
		); 

/******************* CELL 2487 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2487 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2391]),
			.N(gen[2392]),
			.NE(gen[2393]),

			.O(gen[2486]),
			.E(gen[2488]),

			.SO(gen[2581]),
			.S(gen[2582]),
			.SE(gen[2583]),

			.SELF(gen[2487]),
			.cell_state(gen[2487])
		); 

/******************* CELL 2488 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2488 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2392]),
			.N(gen[2393]),
			.NE(gen[2394]),

			.O(gen[2487]),
			.E(gen[2489]),

			.SO(gen[2582]),
			.S(gen[2583]),
			.SE(gen[2584]),

			.SELF(gen[2488]),
			.cell_state(gen[2488])
		); 

/******************* CELL 2489 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2489 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2393]),
			.N(gen[2394]),
			.NE(gen[2395]),

			.O(gen[2488]),
			.E(gen[2490]),

			.SO(gen[2583]),
			.S(gen[2584]),
			.SE(gen[2585]),

			.SELF(gen[2489]),
			.cell_state(gen[2489])
		); 

/******************* CELL 2490 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2490 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2394]),
			.N(gen[2395]),
			.NE(gen[2396]),

			.O(gen[2489]),
			.E(gen[2491]),

			.SO(gen[2584]),
			.S(gen[2585]),
			.SE(gen[2586]),

			.SELF(gen[2490]),
			.cell_state(gen[2490])
		); 

/******************* CELL 2491 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2491 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2395]),
			.N(gen[2396]),
			.NE(gen[2397]),

			.O(gen[2490]),
			.E(gen[2492]),

			.SO(gen[2585]),
			.S(gen[2586]),
			.SE(gen[2587]),

			.SELF(gen[2491]),
			.cell_state(gen[2491])
		); 

/******************* CELL 2492 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2492 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2396]),
			.N(gen[2397]),
			.NE(gen[2398]),

			.O(gen[2491]),
			.E(gen[2493]),

			.SO(gen[2586]),
			.S(gen[2587]),
			.SE(gen[2588]),

			.SELF(gen[2492]),
			.cell_state(gen[2492])
		); 

/******************* CELL 2493 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2493 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2397]),
			.N(gen[2398]),
			.NE(gen[2399]),

			.O(gen[2492]),
			.E(gen[2494]),

			.SO(gen[2587]),
			.S(gen[2588]),
			.SE(gen[2589]),

			.SELF(gen[2493]),
			.cell_state(gen[2493])
		); 

/******************* CELL 2494 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2494 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2398]),
			.N(gen[2399]),
			.NE(gen[2400]),

			.O(gen[2493]),
			.E(gen[2495]),

			.SO(gen[2588]),
			.S(gen[2589]),
			.SE(gen[2590]),

			.SELF(gen[2494]),
			.cell_state(gen[2494])
		); 

/******************* CELL 2495 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2495 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2399]),
			.N(gen[2400]),
			.NE(gen[2401]),

			.O(gen[2494]),
			.E(gen[2496]),

			.SO(gen[2589]),
			.S(gen[2590]),
			.SE(gen[2591]),

			.SELF(gen[2495]),
			.cell_state(gen[2495])
		); 

/******************* CELL 2496 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2496 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2400]),
			.N(gen[2401]),
			.NE(gen[2402]),

			.O(gen[2495]),
			.E(gen[2497]),

			.SO(gen[2590]),
			.S(gen[2591]),
			.SE(gen[2592]),

			.SELF(gen[2496]),
			.cell_state(gen[2496])
		); 

/******************* CELL 2497 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2497 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2401]),
			.N(gen[2402]),
			.NE(gen[2403]),

			.O(gen[2496]),
			.E(gen[2498]),

			.SO(gen[2591]),
			.S(gen[2592]),
			.SE(gen[2593]),

			.SELF(gen[2497]),
			.cell_state(gen[2497])
		); 

/******************* CELL 2498 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2498 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2402]),
			.N(gen[2403]),
			.NE(gen[2404]),

			.O(gen[2497]),
			.E(gen[2499]),

			.SO(gen[2592]),
			.S(gen[2593]),
			.SE(gen[2594]),

			.SELF(gen[2498]),
			.cell_state(gen[2498])
		); 

/******************* CELL 2499 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2499 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2403]),
			.N(gen[2404]),
			.NE(gen[2405]),

			.O(gen[2498]),
			.E(gen[2500]),

			.SO(gen[2593]),
			.S(gen[2594]),
			.SE(gen[2595]),

			.SELF(gen[2499]),
			.cell_state(gen[2499])
		); 

/******************* CELL 2500 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2500 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2404]),
			.N(gen[2405]),
			.NE(gen[2406]),

			.O(gen[2499]),
			.E(gen[2501]),

			.SO(gen[2594]),
			.S(gen[2595]),
			.SE(gen[2596]),

			.SELF(gen[2500]),
			.cell_state(gen[2500])
		); 

/******************* CELL 2501 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2501 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2405]),
			.N(gen[2406]),
			.NE(gen[2407]),

			.O(gen[2500]),
			.E(gen[2502]),

			.SO(gen[2595]),
			.S(gen[2596]),
			.SE(gen[2597]),

			.SELF(gen[2501]),
			.cell_state(gen[2501])
		); 

/******************* CELL 2502 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2502 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2406]),
			.N(gen[2407]),
			.NE(gen[2408]),

			.O(gen[2501]),
			.E(gen[2503]),

			.SO(gen[2596]),
			.S(gen[2597]),
			.SE(gen[2598]),

			.SELF(gen[2502]),
			.cell_state(gen[2502])
		); 

/******************* CELL 2503 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2503 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2407]),
			.N(gen[2408]),
			.NE(gen[2409]),

			.O(gen[2502]),
			.E(gen[2504]),

			.SO(gen[2597]),
			.S(gen[2598]),
			.SE(gen[2599]),

			.SELF(gen[2503]),
			.cell_state(gen[2503])
		); 

/******************* CELL 2504 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2504 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2408]),
			.N(gen[2409]),
			.NE(gen[2410]),

			.O(gen[2503]),
			.E(gen[2505]),

			.SO(gen[2598]),
			.S(gen[2599]),
			.SE(gen[2600]),

			.SELF(gen[2504]),
			.cell_state(gen[2504])
		); 

/******************* CELL 2505 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2505 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2409]),
			.N(gen[2410]),
			.NE(gen[2411]),

			.O(gen[2504]),
			.E(gen[2506]),

			.SO(gen[2599]),
			.S(gen[2600]),
			.SE(gen[2601]),

			.SELF(gen[2505]),
			.cell_state(gen[2505])
		); 

/******************* CELL 2506 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2506 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2410]),
			.N(gen[2411]),
			.NE(gen[2412]),

			.O(gen[2505]),
			.E(gen[2507]),

			.SO(gen[2600]),
			.S(gen[2601]),
			.SE(gen[2602]),

			.SELF(gen[2506]),
			.cell_state(gen[2506])
		); 

/******************* CELL 2507 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2507 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2411]),
			.N(gen[2412]),
			.NE(gen[2413]),

			.O(gen[2506]),
			.E(gen[2508]),

			.SO(gen[2601]),
			.S(gen[2602]),
			.SE(gen[2603]),

			.SELF(gen[2507]),
			.cell_state(gen[2507])
		); 

/******************* CELL 2508 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2508 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2412]),
			.N(gen[2413]),
			.NE(gen[2414]),

			.O(gen[2507]),
			.E(gen[2509]),

			.SO(gen[2602]),
			.S(gen[2603]),
			.SE(gen[2604]),

			.SELF(gen[2508]),
			.cell_state(gen[2508])
		); 

/******************* CELL 2509 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2509 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2413]),
			.N(gen[2414]),
			.NE(gen[2415]),

			.O(gen[2508]),
			.E(gen[2510]),

			.SO(gen[2603]),
			.S(gen[2604]),
			.SE(gen[2605]),

			.SELF(gen[2509]),
			.cell_state(gen[2509])
		); 

/******************* CELL 2510 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2510 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2414]),
			.N(gen[2415]),
			.NE(gen[2416]),

			.O(gen[2509]),
			.E(gen[2511]),

			.SO(gen[2604]),
			.S(gen[2605]),
			.SE(gen[2606]),

			.SELF(gen[2510]),
			.cell_state(gen[2510])
		); 

/******************* CELL 2511 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2511 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2415]),
			.N(gen[2416]),
			.NE(gen[2417]),

			.O(gen[2510]),
			.E(gen[2512]),

			.SO(gen[2605]),
			.S(gen[2606]),
			.SE(gen[2607]),

			.SELF(gen[2511]),
			.cell_state(gen[2511])
		); 

/******************* CELL 2512 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2512 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2416]),
			.N(gen[2417]),
			.NE(gen[2418]),

			.O(gen[2511]),
			.E(gen[2513]),

			.SO(gen[2606]),
			.S(gen[2607]),
			.SE(gen[2608]),

			.SELF(gen[2512]),
			.cell_state(gen[2512])
		); 

/******************* CELL 2513 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2513 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2417]),
			.N(gen[2418]),
			.NE(gen[2419]),

			.O(gen[2512]),
			.E(gen[2514]),

			.SO(gen[2607]),
			.S(gen[2608]),
			.SE(gen[2609]),

			.SELF(gen[2513]),
			.cell_state(gen[2513])
		); 

/******************* CELL 2514 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2514 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2418]),
			.N(gen[2419]),
			.NE(gen[2420]),

			.O(gen[2513]),
			.E(gen[2515]),

			.SO(gen[2608]),
			.S(gen[2609]),
			.SE(gen[2610]),

			.SELF(gen[2514]),
			.cell_state(gen[2514])
		); 

/******************* CELL 2515 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2515 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2419]),
			.N(gen[2420]),
			.NE(gen[2421]),

			.O(gen[2514]),
			.E(gen[2516]),

			.SO(gen[2609]),
			.S(gen[2610]),
			.SE(gen[2611]),

			.SELF(gen[2515]),
			.cell_state(gen[2515])
		); 

/******************* CELL 2516 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2516 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2420]),
			.N(gen[2421]),
			.NE(gen[2422]),

			.O(gen[2515]),
			.E(gen[2517]),

			.SO(gen[2610]),
			.S(gen[2611]),
			.SE(gen[2612]),

			.SELF(gen[2516]),
			.cell_state(gen[2516])
		); 

/******************* CELL 2517 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2517 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2421]),
			.N(gen[2422]),
			.NE(gen[2423]),

			.O(gen[2516]),
			.E(gen[2518]),

			.SO(gen[2611]),
			.S(gen[2612]),
			.SE(gen[2613]),

			.SELF(gen[2517]),
			.cell_state(gen[2517])
		); 

/******************* CELL 2518 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2518 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2422]),
			.N(gen[2423]),
			.NE(gen[2424]),

			.O(gen[2517]),
			.E(gen[2519]),

			.SO(gen[2612]),
			.S(gen[2613]),
			.SE(gen[2614]),

			.SELF(gen[2518]),
			.cell_state(gen[2518])
		); 

/******************* CELL 2519 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2519 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2423]),
			.N(gen[2424]),
			.NE(gen[2425]),

			.O(gen[2518]),
			.E(gen[2520]),

			.SO(gen[2613]),
			.S(gen[2614]),
			.SE(gen[2615]),

			.SELF(gen[2519]),
			.cell_state(gen[2519])
		); 

/******************* CELL 2520 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2520 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2424]),
			.N(gen[2425]),
			.NE(gen[2426]),

			.O(gen[2519]),
			.E(gen[2521]),

			.SO(gen[2614]),
			.S(gen[2615]),
			.SE(gen[2616]),

			.SELF(gen[2520]),
			.cell_state(gen[2520])
		); 

/******************* CELL 2521 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2521 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2425]),
			.N(gen[2426]),
			.NE(gen[2427]),

			.O(gen[2520]),
			.E(gen[2522]),

			.SO(gen[2615]),
			.S(gen[2616]),
			.SE(gen[2617]),

			.SELF(gen[2521]),
			.cell_state(gen[2521])
		); 

/******************* CELL 2522 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2522 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2426]),
			.N(gen[2427]),
			.NE(gen[2428]),

			.O(gen[2521]),
			.E(gen[2523]),

			.SO(gen[2616]),
			.S(gen[2617]),
			.SE(gen[2618]),

			.SELF(gen[2522]),
			.cell_state(gen[2522])
		); 

/******************* CELL 2523 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2523 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2427]),
			.N(gen[2428]),
			.NE(gen[2429]),

			.O(gen[2522]),
			.E(gen[2524]),

			.SO(gen[2617]),
			.S(gen[2618]),
			.SE(gen[2619]),

			.SELF(gen[2523]),
			.cell_state(gen[2523])
		); 

/******************* CELL 2524 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2524 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2428]),
			.N(gen[2429]),
			.NE(gen[2430]),

			.O(gen[2523]),
			.E(gen[2525]),

			.SO(gen[2618]),
			.S(gen[2619]),
			.SE(gen[2620]),

			.SELF(gen[2524]),
			.cell_state(gen[2524])
		); 

/******************* CELL 2525 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2525 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2429]),
			.N(gen[2430]),
			.NE(gen[2431]),

			.O(gen[2524]),
			.E(gen[2526]),

			.SO(gen[2619]),
			.S(gen[2620]),
			.SE(gen[2621]),

			.SELF(gen[2525]),
			.cell_state(gen[2525])
		); 

/******************* CELL 2526 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2526 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2430]),
			.N(gen[2431]),
			.NE(gen[2432]),

			.O(gen[2525]),
			.E(gen[2527]),

			.SO(gen[2620]),
			.S(gen[2621]),
			.SE(gen[2622]),

			.SELF(gen[2526]),
			.cell_state(gen[2526])
		); 

/******************* CELL 2527 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2527 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2431]),
			.N(gen[2432]),
			.NE(gen[2433]),

			.O(gen[2526]),
			.E(gen[2528]),

			.SO(gen[2621]),
			.S(gen[2622]),
			.SE(gen[2623]),

			.SELF(gen[2527]),
			.cell_state(gen[2527])
		); 

/******************* CELL 2528 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2528 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2432]),
			.N(gen[2433]),
			.NE(gen[2434]),

			.O(gen[2527]),
			.E(gen[2529]),

			.SO(gen[2622]),
			.S(gen[2623]),
			.SE(gen[2624]),

			.SELF(gen[2528]),
			.cell_state(gen[2528])
		); 

/******************* CELL 2529 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2529 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2433]),
			.N(gen[2434]),
			.NE(gen[2435]),

			.O(gen[2528]),
			.E(gen[2530]),

			.SO(gen[2623]),
			.S(gen[2624]),
			.SE(gen[2625]),

			.SELF(gen[2529]),
			.cell_state(gen[2529])
		); 

/******************* CELL 2530 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2530 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2434]),
			.N(gen[2435]),
			.NE(gen[2436]),

			.O(gen[2529]),
			.E(gen[2531]),

			.SO(gen[2624]),
			.S(gen[2625]),
			.SE(gen[2626]),

			.SELF(gen[2530]),
			.cell_state(gen[2530])
		); 

/******************* CELL 2531 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2531 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2435]),
			.N(gen[2436]),
			.NE(gen[2437]),

			.O(gen[2530]),
			.E(gen[2532]),

			.SO(gen[2625]),
			.S(gen[2626]),
			.SE(gen[2627]),

			.SELF(gen[2531]),
			.cell_state(gen[2531])
		); 

/******************* CELL 2532 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2532 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2436]),
			.N(gen[2437]),
			.NE(gen[2438]),

			.O(gen[2531]),
			.E(gen[2533]),

			.SO(gen[2626]),
			.S(gen[2627]),
			.SE(gen[2628]),

			.SELF(gen[2532]),
			.cell_state(gen[2532])
		); 

/******************* CELL 2533 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2533 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2437]),
			.N(gen[2438]),
			.NE(gen[2439]),

			.O(gen[2532]),
			.E(gen[2534]),

			.SO(gen[2627]),
			.S(gen[2628]),
			.SE(gen[2629]),

			.SELF(gen[2533]),
			.cell_state(gen[2533])
		); 

/******************* CELL 2534 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2534 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2438]),
			.N(gen[2439]),
			.NE(gen[2440]),

			.O(gen[2533]),
			.E(gen[2535]),

			.SO(gen[2628]),
			.S(gen[2629]),
			.SE(gen[2630]),

			.SELF(gen[2534]),
			.cell_state(gen[2534])
		); 

/******************* CELL 2535 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2535 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2439]),
			.N(gen[2440]),
			.NE(gen[2441]),

			.O(gen[2534]),
			.E(gen[2536]),

			.SO(gen[2629]),
			.S(gen[2630]),
			.SE(gen[2631]),

			.SELF(gen[2535]),
			.cell_state(gen[2535])
		); 

/******************* CELL 2536 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2536 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2440]),
			.N(gen[2441]),
			.NE(gen[2442]),

			.O(gen[2535]),
			.E(gen[2537]),

			.SO(gen[2630]),
			.S(gen[2631]),
			.SE(gen[2632]),

			.SELF(gen[2536]),
			.cell_state(gen[2536])
		); 

/******************* CELL 2537 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2537 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2441]),
			.N(gen[2442]),
			.NE(gen[2443]),

			.O(gen[2536]),
			.E(gen[2538]),

			.SO(gen[2631]),
			.S(gen[2632]),
			.SE(gen[2633]),

			.SELF(gen[2537]),
			.cell_state(gen[2537])
		); 

/******************* CELL 2538 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2538 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2442]),
			.N(gen[2443]),
			.NE(gen[2444]),

			.O(gen[2537]),
			.E(gen[2539]),

			.SO(gen[2632]),
			.S(gen[2633]),
			.SE(gen[2634]),

			.SELF(gen[2538]),
			.cell_state(gen[2538])
		); 

/******************* CELL 2539 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2539 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2443]),
			.N(gen[2444]),
			.NE(gen[2445]),

			.O(gen[2538]),
			.E(gen[2540]),

			.SO(gen[2633]),
			.S(gen[2634]),
			.SE(gen[2635]),

			.SELF(gen[2539]),
			.cell_state(gen[2539])
		); 

/******************* CELL 2540 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2540 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2444]),
			.N(gen[2445]),
			.NE(gen[2446]),

			.O(gen[2539]),
			.E(gen[2541]),

			.SO(gen[2634]),
			.S(gen[2635]),
			.SE(gen[2636]),

			.SELF(gen[2540]),
			.cell_state(gen[2540])
		); 

/******************* CELL 2541 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2541 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2445]),
			.N(gen[2446]),
			.NE(gen[2447]),

			.O(gen[2540]),
			.E(gen[2542]),

			.SO(gen[2635]),
			.S(gen[2636]),
			.SE(gen[2637]),

			.SELF(gen[2541]),
			.cell_state(gen[2541])
		); 

/******************* CELL 2542 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2542 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2446]),
			.N(gen[2447]),
			.NE(gen[2448]),

			.O(gen[2541]),
			.E(gen[2543]),

			.SO(gen[2636]),
			.S(gen[2637]),
			.SE(gen[2638]),

			.SELF(gen[2542]),
			.cell_state(gen[2542])
		); 

/******************* CELL 2543 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2543 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2447]),
			.N(gen[2448]),
			.NE(gen[2449]),

			.O(gen[2542]),
			.E(gen[2544]),

			.SO(gen[2637]),
			.S(gen[2638]),
			.SE(gen[2639]),

			.SELF(gen[2543]),
			.cell_state(gen[2543])
		); 

/******************* CELL 2544 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2544 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2448]),
			.N(gen[2449]),
			.NE(gen[2450]),

			.O(gen[2543]),
			.E(gen[2545]),

			.SO(gen[2638]),
			.S(gen[2639]),
			.SE(gen[2640]),

			.SELF(gen[2544]),
			.cell_state(gen[2544])
		); 

/******************* CELL 2545 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2545 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2449]),
			.N(gen[2450]),
			.NE(gen[2451]),

			.O(gen[2544]),
			.E(gen[2546]),

			.SO(gen[2639]),
			.S(gen[2640]),
			.SE(gen[2641]),

			.SELF(gen[2545]),
			.cell_state(gen[2545])
		); 

/******************* CELL 2546 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2546 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2450]),
			.N(gen[2451]),
			.NE(gen[2452]),

			.O(gen[2545]),
			.E(gen[2547]),

			.SO(gen[2640]),
			.S(gen[2641]),
			.SE(gen[2642]),

			.SELF(gen[2546]),
			.cell_state(gen[2546])
		); 

/******************* CELL 2547 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2547 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2451]),
			.N(gen[2452]),
			.NE(gen[2453]),

			.O(gen[2546]),
			.E(gen[2548]),

			.SO(gen[2641]),
			.S(gen[2642]),
			.SE(gen[2643]),

			.SELF(gen[2547]),
			.cell_state(gen[2547])
		); 

/******************* CELL 2548 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2548 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2452]),
			.N(gen[2453]),
			.NE(gen[2454]),

			.O(gen[2547]),
			.E(gen[2549]),

			.SO(gen[2642]),
			.S(gen[2643]),
			.SE(gen[2644]),

			.SELF(gen[2548]),
			.cell_state(gen[2548])
		); 

/******************* CELL 2549 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2549 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2453]),
			.N(gen[2454]),
			.NE(gen[2455]),

			.O(gen[2548]),
			.E(gen[2550]),

			.SO(gen[2643]),
			.S(gen[2644]),
			.SE(gen[2645]),

			.SELF(gen[2549]),
			.cell_state(gen[2549])
		); 

/******************* CELL 2550 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2550 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2454]),
			.N(gen[2455]),
			.NE(gen[2456]),

			.O(gen[2549]),
			.E(gen[2551]),

			.SO(gen[2644]),
			.S(gen[2645]),
			.SE(gen[2646]),

			.SELF(gen[2550]),
			.cell_state(gen[2550])
		); 

/******************* CELL 2551 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2551 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2455]),
			.N(gen[2456]),
			.NE(gen[2457]),

			.O(gen[2550]),
			.E(gen[2552]),

			.SO(gen[2645]),
			.S(gen[2646]),
			.SE(gen[2647]),

			.SELF(gen[2551]),
			.cell_state(gen[2551])
		); 

/******************* CELL 2552 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2552 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2456]),
			.N(gen[2457]),
			.NE(gen[2458]),

			.O(gen[2551]),
			.E(gen[2553]),

			.SO(gen[2646]),
			.S(gen[2647]),
			.SE(gen[2648]),

			.SELF(gen[2552]),
			.cell_state(gen[2552])
		); 

/******************* CELL 2553 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2553 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2457]),
			.N(gen[2458]),
			.NE(gen[2459]),

			.O(gen[2552]),
			.E(gen[2554]),

			.SO(gen[2647]),
			.S(gen[2648]),
			.SE(gen[2649]),

			.SELF(gen[2553]),
			.cell_state(gen[2553])
		); 

/******************* CELL 2554 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2554 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2458]),
			.N(gen[2459]),
			.NE(gen[2460]),

			.O(gen[2553]),
			.E(gen[2555]),

			.SO(gen[2648]),
			.S(gen[2649]),
			.SE(gen[2650]),

			.SELF(gen[2554]),
			.cell_state(gen[2554])
		); 

/******************* CELL 2555 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2555 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2459]),
			.N(gen[2460]),
			.NE(gen[2461]),

			.O(gen[2554]),
			.E(gen[2556]),

			.SO(gen[2649]),
			.S(gen[2650]),
			.SE(gen[2651]),

			.SELF(gen[2555]),
			.cell_state(gen[2555])
		); 

/******************* CELL 2556 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2556 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2460]),
			.N(gen[2461]),
			.NE(gen[2462]),

			.O(gen[2555]),
			.E(gen[2557]),

			.SO(gen[2650]),
			.S(gen[2651]),
			.SE(gen[2652]),

			.SELF(gen[2556]),
			.cell_state(gen[2556])
		); 

/******************* CELL 2557 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2557 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2461]),
			.N(gen[2462]),
			.NE(gen[2463]),

			.O(gen[2556]),
			.E(gen[2558]),

			.SO(gen[2651]),
			.S(gen[2652]),
			.SE(gen[2653]),

			.SELF(gen[2557]),
			.cell_state(gen[2557])
		); 

/******************* CELL 2558 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2558 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2462]),
			.N(gen[2463]),
			.NE(gen[2464]),

			.O(gen[2557]),
			.E(gen[2559]),

			.SO(gen[2652]),
			.S(gen[2653]),
			.SE(gen[2654]),

			.SELF(gen[2558]),
			.cell_state(gen[2558])
		); 

/******************* CELL 2559 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2559 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2463]),
			.N(gen[2464]),
			.NE(gen[2465]),

			.O(gen[2558]),
			.E(gen[2560]),

			.SO(gen[2653]),
			.S(gen[2654]),
			.SE(gen[2655]),

			.SELF(gen[2559]),
			.cell_state(gen[2559])
		); 

/******************* CELL 2560 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2560 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2464]),
			.N(gen[2465]),
			.NE(gen[2466]),

			.O(gen[2559]),
			.E(gen[2561]),

			.SO(gen[2654]),
			.S(gen[2655]),
			.SE(gen[2656]),

			.SELF(gen[2560]),
			.cell_state(gen[2560])
		); 

/******************* CELL 2561 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2561 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2465]),
			.N(gen[2466]),
			.NE(gen[2467]),

			.O(gen[2560]),
			.E(gen[2562]),

			.SO(gen[2655]),
			.S(gen[2656]),
			.SE(gen[2657]),

			.SELF(gen[2561]),
			.cell_state(gen[2561])
		); 

/******************* CELL 2562 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2562 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2466]),
			.N(gen[2467]),
			.NE(gen[2468]),

			.O(gen[2561]),
			.E(gen[2563]),

			.SO(gen[2656]),
			.S(gen[2657]),
			.SE(gen[2658]),

			.SELF(gen[2562]),
			.cell_state(gen[2562])
		); 

/******************* CELL 2563 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2563 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2467]),
			.N(gen[2468]),
			.NE(gen[2469]),

			.O(gen[2562]),
			.E(gen[2564]),

			.SO(gen[2657]),
			.S(gen[2658]),
			.SE(gen[2659]),

			.SELF(gen[2563]),
			.cell_state(gen[2563])
		); 

/******************* CELL 2564 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2564 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2468]),
			.N(gen[2469]),
			.NE(gen[2468]),

			.O(gen[2563]),
			.E(gen[2563]),

			.SO(gen[2658]),
			.S(gen[2659]),
			.SE(gen[2658]),

			.SELF(gen[2564]),
			.cell_state(gen[2564])
		); 

/******************* CELL 2565 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2565 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2471]),
			.N(gen[2470]),
			.NE(gen[2471]),

			.O(gen[2566]),
			.E(gen[2566]),

			.SO(gen[2661]),
			.S(gen[2660]),
			.SE(gen[2661]),

			.SELF(gen[2565]),
			.cell_state(gen[2565])
		); 

/******************* CELL 2566 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2566 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2470]),
			.N(gen[2471]),
			.NE(gen[2472]),

			.O(gen[2565]),
			.E(gen[2567]),

			.SO(gen[2660]),
			.S(gen[2661]),
			.SE(gen[2662]),

			.SELF(gen[2566]),
			.cell_state(gen[2566])
		); 

/******************* CELL 2567 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2567 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2471]),
			.N(gen[2472]),
			.NE(gen[2473]),

			.O(gen[2566]),
			.E(gen[2568]),

			.SO(gen[2661]),
			.S(gen[2662]),
			.SE(gen[2663]),

			.SELF(gen[2567]),
			.cell_state(gen[2567])
		); 

/******************* CELL 2568 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2568 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2472]),
			.N(gen[2473]),
			.NE(gen[2474]),

			.O(gen[2567]),
			.E(gen[2569]),

			.SO(gen[2662]),
			.S(gen[2663]),
			.SE(gen[2664]),

			.SELF(gen[2568]),
			.cell_state(gen[2568])
		); 

/******************* CELL 2569 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2569 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2473]),
			.N(gen[2474]),
			.NE(gen[2475]),

			.O(gen[2568]),
			.E(gen[2570]),

			.SO(gen[2663]),
			.S(gen[2664]),
			.SE(gen[2665]),

			.SELF(gen[2569]),
			.cell_state(gen[2569])
		); 

/******************* CELL 2570 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2570 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2474]),
			.N(gen[2475]),
			.NE(gen[2476]),

			.O(gen[2569]),
			.E(gen[2571]),

			.SO(gen[2664]),
			.S(gen[2665]),
			.SE(gen[2666]),

			.SELF(gen[2570]),
			.cell_state(gen[2570])
		); 

/******************* CELL 2571 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2571 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2475]),
			.N(gen[2476]),
			.NE(gen[2477]),

			.O(gen[2570]),
			.E(gen[2572]),

			.SO(gen[2665]),
			.S(gen[2666]),
			.SE(gen[2667]),

			.SELF(gen[2571]),
			.cell_state(gen[2571])
		); 

/******************* CELL 2572 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2572 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2476]),
			.N(gen[2477]),
			.NE(gen[2478]),

			.O(gen[2571]),
			.E(gen[2573]),

			.SO(gen[2666]),
			.S(gen[2667]),
			.SE(gen[2668]),

			.SELF(gen[2572]),
			.cell_state(gen[2572])
		); 

/******************* CELL 2573 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2573 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2477]),
			.N(gen[2478]),
			.NE(gen[2479]),

			.O(gen[2572]),
			.E(gen[2574]),

			.SO(gen[2667]),
			.S(gen[2668]),
			.SE(gen[2669]),

			.SELF(gen[2573]),
			.cell_state(gen[2573])
		); 

/******************* CELL 2574 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2574 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2478]),
			.N(gen[2479]),
			.NE(gen[2480]),

			.O(gen[2573]),
			.E(gen[2575]),

			.SO(gen[2668]),
			.S(gen[2669]),
			.SE(gen[2670]),

			.SELF(gen[2574]),
			.cell_state(gen[2574])
		); 

/******************* CELL 2575 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2575 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2479]),
			.N(gen[2480]),
			.NE(gen[2481]),

			.O(gen[2574]),
			.E(gen[2576]),

			.SO(gen[2669]),
			.S(gen[2670]),
			.SE(gen[2671]),

			.SELF(gen[2575]),
			.cell_state(gen[2575])
		); 

/******************* CELL 2576 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2576 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2480]),
			.N(gen[2481]),
			.NE(gen[2482]),

			.O(gen[2575]),
			.E(gen[2577]),

			.SO(gen[2670]),
			.S(gen[2671]),
			.SE(gen[2672]),

			.SELF(gen[2576]),
			.cell_state(gen[2576])
		); 

/******************* CELL 2577 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2577 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2481]),
			.N(gen[2482]),
			.NE(gen[2483]),

			.O(gen[2576]),
			.E(gen[2578]),

			.SO(gen[2671]),
			.S(gen[2672]),
			.SE(gen[2673]),

			.SELF(gen[2577]),
			.cell_state(gen[2577])
		); 

/******************* CELL 2578 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2578 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2482]),
			.N(gen[2483]),
			.NE(gen[2484]),

			.O(gen[2577]),
			.E(gen[2579]),

			.SO(gen[2672]),
			.S(gen[2673]),
			.SE(gen[2674]),

			.SELF(gen[2578]),
			.cell_state(gen[2578])
		); 

/******************* CELL 2579 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2579 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2483]),
			.N(gen[2484]),
			.NE(gen[2485]),

			.O(gen[2578]),
			.E(gen[2580]),

			.SO(gen[2673]),
			.S(gen[2674]),
			.SE(gen[2675]),

			.SELF(gen[2579]),
			.cell_state(gen[2579])
		); 

/******************* CELL 2580 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2580 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2484]),
			.N(gen[2485]),
			.NE(gen[2486]),

			.O(gen[2579]),
			.E(gen[2581]),

			.SO(gen[2674]),
			.S(gen[2675]),
			.SE(gen[2676]),

			.SELF(gen[2580]),
			.cell_state(gen[2580])
		); 

/******************* CELL 2581 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2581 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2485]),
			.N(gen[2486]),
			.NE(gen[2487]),

			.O(gen[2580]),
			.E(gen[2582]),

			.SO(gen[2675]),
			.S(gen[2676]),
			.SE(gen[2677]),

			.SELF(gen[2581]),
			.cell_state(gen[2581])
		); 

/******************* CELL 2582 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2582 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2486]),
			.N(gen[2487]),
			.NE(gen[2488]),

			.O(gen[2581]),
			.E(gen[2583]),

			.SO(gen[2676]),
			.S(gen[2677]),
			.SE(gen[2678]),

			.SELF(gen[2582]),
			.cell_state(gen[2582])
		); 

/******************* CELL 2583 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2583 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2487]),
			.N(gen[2488]),
			.NE(gen[2489]),

			.O(gen[2582]),
			.E(gen[2584]),

			.SO(gen[2677]),
			.S(gen[2678]),
			.SE(gen[2679]),

			.SELF(gen[2583]),
			.cell_state(gen[2583])
		); 

/******************* CELL 2584 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2584 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2488]),
			.N(gen[2489]),
			.NE(gen[2490]),

			.O(gen[2583]),
			.E(gen[2585]),

			.SO(gen[2678]),
			.S(gen[2679]),
			.SE(gen[2680]),

			.SELF(gen[2584]),
			.cell_state(gen[2584])
		); 

/******************* CELL 2585 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2585 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2489]),
			.N(gen[2490]),
			.NE(gen[2491]),

			.O(gen[2584]),
			.E(gen[2586]),

			.SO(gen[2679]),
			.S(gen[2680]),
			.SE(gen[2681]),

			.SELF(gen[2585]),
			.cell_state(gen[2585])
		); 

/******************* CELL 2586 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2586 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2490]),
			.N(gen[2491]),
			.NE(gen[2492]),

			.O(gen[2585]),
			.E(gen[2587]),

			.SO(gen[2680]),
			.S(gen[2681]),
			.SE(gen[2682]),

			.SELF(gen[2586]),
			.cell_state(gen[2586])
		); 

/******************* CELL 2587 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2587 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2491]),
			.N(gen[2492]),
			.NE(gen[2493]),

			.O(gen[2586]),
			.E(gen[2588]),

			.SO(gen[2681]),
			.S(gen[2682]),
			.SE(gen[2683]),

			.SELF(gen[2587]),
			.cell_state(gen[2587])
		); 

/******************* CELL 2588 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2588 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2492]),
			.N(gen[2493]),
			.NE(gen[2494]),

			.O(gen[2587]),
			.E(gen[2589]),

			.SO(gen[2682]),
			.S(gen[2683]),
			.SE(gen[2684]),

			.SELF(gen[2588]),
			.cell_state(gen[2588])
		); 

/******************* CELL 2589 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2589 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2493]),
			.N(gen[2494]),
			.NE(gen[2495]),

			.O(gen[2588]),
			.E(gen[2590]),

			.SO(gen[2683]),
			.S(gen[2684]),
			.SE(gen[2685]),

			.SELF(gen[2589]),
			.cell_state(gen[2589])
		); 

/******************* CELL 2590 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2590 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2494]),
			.N(gen[2495]),
			.NE(gen[2496]),

			.O(gen[2589]),
			.E(gen[2591]),

			.SO(gen[2684]),
			.S(gen[2685]),
			.SE(gen[2686]),

			.SELF(gen[2590]),
			.cell_state(gen[2590])
		); 

/******************* CELL 2591 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2591 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2495]),
			.N(gen[2496]),
			.NE(gen[2497]),

			.O(gen[2590]),
			.E(gen[2592]),

			.SO(gen[2685]),
			.S(gen[2686]),
			.SE(gen[2687]),

			.SELF(gen[2591]),
			.cell_state(gen[2591])
		); 

/******************* CELL 2592 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2592 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2496]),
			.N(gen[2497]),
			.NE(gen[2498]),

			.O(gen[2591]),
			.E(gen[2593]),

			.SO(gen[2686]),
			.S(gen[2687]),
			.SE(gen[2688]),

			.SELF(gen[2592]),
			.cell_state(gen[2592])
		); 

/******************* CELL 2593 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2593 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2497]),
			.N(gen[2498]),
			.NE(gen[2499]),

			.O(gen[2592]),
			.E(gen[2594]),

			.SO(gen[2687]),
			.S(gen[2688]),
			.SE(gen[2689]),

			.SELF(gen[2593]),
			.cell_state(gen[2593])
		); 

/******************* CELL 2594 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2594 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2498]),
			.N(gen[2499]),
			.NE(gen[2500]),

			.O(gen[2593]),
			.E(gen[2595]),

			.SO(gen[2688]),
			.S(gen[2689]),
			.SE(gen[2690]),

			.SELF(gen[2594]),
			.cell_state(gen[2594])
		); 

/******************* CELL 2595 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2595 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2499]),
			.N(gen[2500]),
			.NE(gen[2501]),

			.O(gen[2594]),
			.E(gen[2596]),

			.SO(gen[2689]),
			.S(gen[2690]),
			.SE(gen[2691]),

			.SELF(gen[2595]),
			.cell_state(gen[2595])
		); 

/******************* CELL 2596 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2596 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2500]),
			.N(gen[2501]),
			.NE(gen[2502]),

			.O(gen[2595]),
			.E(gen[2597]),

			.SO(gen[2690]),
			.S(gen[2691]),
			.SE(gen[2692]),

			.SELF(gen[2596]),
			.cell_state(gen[2596])
		); 

/******************* CELL 2597 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2597 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2501]),
			.N(gen[2502]),
			.NE(gen[2503]),

			.O(gen[2596]),
			.E(gen[2598]),

			.SO(gen[2691]),
			.S(gen[2692]),
			.SE(gen[2693]),

			.SELF(gen[2597]),
			.cell_state(gen[2597])
		); 

/******************* CELL 2598 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2598 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2502]),
			.N(gen[2503]),
			.NE(gen[2504]),

			.O(gen[2597]),
			.E(gen[2599]),

			.SO(gen[2692]),
			.S(gen[2693]),
			.SE(gen[2694]),

			.SELF(gen[2598]),
			.cell_state(gen[2598])
		); 

/******************* CELL 2599 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2599 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2503]),
			.N(gen[2504]),
			.NE(gen[2505]),

			.O(gen[2598]),
			.E(gen[2600]),

			.SO(gen[2693]),
			.S(gen[2694]),
			.SE(gen[2695]),

			.SELF(gen[2599]),
			.cell_state(gen[2599])
		); 

/******************* CELL 2600 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2600 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2504]),
			.N(gen[2505]),
			.NE(gen[2506]),

			.O(gen[2599]),
			.E(gen[2601]),

			.SO(gen[2694]),
			.S(gen[2695]),
			.SE(gen[2696]),

			.SELF(gen[2600]),
			.cell_state(gen[2600])
		); 

/******************* CELL 2601 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2601 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2505]),
			.N(gen[2506]),
			.NE(gen[2507]),

			.O(gen[2600]),
			.E(gen[2602]),

			.SO(gen[2695]),
			.S(gen[2696]),
			.SE(gen[2697]),

			.SELF(gen[2601]),
			.cell_state(gen[2601])
		); 

/******************* CELL 2602 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2602 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2506]),
			.N(gen[2507]),
			.NE(gen[2508]),

			.O(gen[2601]),
			.E(gen[2603]),

			.SO(gen[2696]),
			.S(gen[2697]),
			.SE(gen[2698]),

			.SELF(gen[2602]),
			.cell_state(gen[2602])
		); 

/******************* CELL 2603 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2603 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2507]),
			.N(gen[2508]),
			.NE(gen[2509]),

			.O(gen[2602]),
			.E(gen[2604]),

			.SO(gen[2697]),
			.S(gen[2698]),
			.SE(gen[2699]),

			.SELF(gen[2603]),
			.cell_state(gen[2603])
		); 

/******************* CELL 2604 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2604 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2508]),
			.N(gen[2509]),
			.NE(gen[2510]),

			.O(gen[2603]),
			.E(gen[2605]),

			.SO(gen[2698]),
			.S(gen[2699]),
			.SE(gen[2700]),

			.SELF(gen[2604]),
			.cell_state(gen[2604])
		); 

/******************* CELL 2605 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2605 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2509]),
			.N(gen[2510]),
			.NE(gen[2511]),

			.O(gen[2604]),
			.E(gen[2606]),

			.SO(gen[2699]),
			.S(gen[2700]),
			.SE(gen[2701]),

			.SELF(gen[2605]),
			.cell_state(gen[2605])
		); 

/******************* CELL 2606 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2606 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2510]),
			.N(gen[2511]),
			.NE(gen[2512]),

			.O(gen[2605]),
			.E(gen[2607]),

			.SO(gen[2700]),
			.S(gen[2701]),
			.SE(gen[2702]),

			.SELF(gen[2606]),
			.cell_state(gen[2606])
		); 

/******************* CELL 2607 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2607 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2511]),
			.N(gen[2512]),
			.NE(gen[2513]),

			.O(gen[2606]),
			.E(gen[2608]),

			.SO(gen[2701]),
			.S(gen[2702]),
			.SE(gen[2703]),

			.SELF(gen[2607]),
			.cell_state(gen[2607])
		); 

/******************* CELL 2608 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2608 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2512]),
			.N(gen[2513]),
			.NE(gen[2514]),

			.O(gen[2607]),
			.E(gen[2609]),

			.SO(gen[2702]),
			.S(gen[2703]),
			.SE(gen[2704]),

			.SELF(gen[2608]),
			.cell_state(gen[2608])
		); 

/******************* CELL 2609 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2609 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2513]),
			.N(gen[2514]),
			.NE(gen[2515]),

			.O(gen[2608]),
			.E(gen[2610]),

			.SO(gen[2703]),
			.S(gen[2704]),
			.SE(gen[2705]),

			.SELF(gen[2609]),
			.cell_state(gen[2609])
		); 

/******************* CELL 2610 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2610 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2514]),
			.N(gen[2515]),
			.NE(gen[2516]),

			.O(gen[2609]),
			.E(gen[2611]),

			.SO(gen[2704]),
			.S(gen[2705]),
			.SE(gen[2706]),

			.SELF(gen[2610]),
			.cell_state(gen[2610])
		); 

/******************* CELL 2611 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2611 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2515]),
			.N(gen[2516]),
			.NE(gen[2517]),

			.O(gen[2610]),
			.E(gen[2612]),

			.SO(gen[2705]),
			.S(gen[2706]),
			.SE(gen[2707]),

			.SELF(gen[2611]),
			.cell_state(gen[2611])
		); 

/******************* CELL 2612 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2612 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2516]),
			.N(gen[2517]),
			.NE(gen[2518]),

			.O(gen[2611]),
			.E(gen[2613]),

			.SO(gen[2706]),
			.S(gen[2707]),
			.SE(gen[2708]),

			.SELF(gen[2612]),
			.cell_state(gen[2612])
		); 

/******************* CELL 2613 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2613 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2517]),
			.N(gen[2518]),
			.NE(gen[2519]),

			.O(gen[2612]),
			.E(gen[2614]),

			.SO(gen[2707]),
			.S(gen[2708]),
			.SE(gen[2709]),

			.SELF(gen[2613]),
			.cell_state(gen[2613])
		); 

/******************* CELL 2614 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2614 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2518]),
			.N(gen[2519]),
			.NE(gen[2520]),

			.O(gen[2613]),
			.E(gen[2615]),

			.SO(gen[2708]),
			.S(gen[2709]),
			.SE(gen[2710]),

			.SELF(gen[2614]),
			.cell_state(gen[2614])
		); 

/******************* CELL 2615 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2615 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2519]),
			.N(gen[2520]),
			.NE(gen[2521]),

			.O(gen[2614]),
			.E(gen[2616]),

			.SO(gen[2709]),
			.S(gen[2710]),
			.SE(gen[2711]),

			.SELF(gen[2615]),
			.cell_state(gen[2615])
		); 

/******************* CELL 2616 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2616 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2520]),
			.N(gen[2521]),
			.NE(gen[2522]),

			.O(gen[2615]),
			.E(gen[2617]),

			.SO(gen[2710]),
			.S(gen[2711]),
			.SE(gen[2712]),

			.SELF(gen[2616]),
			.cell_state(gen[2616])
		); 

/******************* CELL 2617 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2617 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2521]),
			.N(gen[2522]),
			.NE(gen[2523]),

			.O(gen[2616]),
			.E(gen[2618]),

			.SO(gen[2711]),
			.S(gen[2712]),
			.SE(gen[2713]),

			.SELF(gen[2617]),
			.cell_state(gen[2617])
		); 

/******************* CELL 2618 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2618 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2522]),
			.N(gen[2523]),
			.NE(gen[2524]),

			.O(gen[2617]),
			.E(gen[2619]),

			.SO(gen[2712]),
			.S(gen[2713]),
			.SE(gen[2714]),

			.SELF(gen[2618]),
			.cell_state(gen[2618])
		); 

/******************* CELL 2619 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2619 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2523]),
			.N(gen[2524]),
			.NE(gen[2525]),

			.O(gen[2618]),
			.E(gen[2620]),

			.SO(gen[2713]),
			.S(gen[2714]),
			.SE(gen[2715]),

			.SELF(gen[2619]),
			.cell_state(gen[2619])
		); 

/******************* CELL 2620 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2620 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2524]),
			.N(gen[2525]),
			.NE(gen[2526]),

			.O(gen[2619]),
			.E(gen[2621]),

			.SO(gen[2714]),
			.S(gen[2715]),
			.SE(gen[2716]),

			.SELF(gen[2620]),
			.cell_state(gen[2620])
		); 

/******************* CELL 2621 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2621 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2525]),
			.N(gen[2526]),
			.NE(gen[2527]),

			.O(gen[2620]),
			.E(gen[2622]),

			.SO(gen[2715]),
			.S(gen[2716]),
			.SE(gen[2717]),

			.SELF(gen[2621]),
			.cell_state(gen[2621])
		); 

/******************* CELL 2622 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2622 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2526]),
			.N(gen[2527]),
			.NE(gen[2528]),

			.O(gen[2621]),
			.E(gen[2623]),

			.SO(gen[2716]),
			.S(gen[2717]),
			.SE(gen[2718]),

			.SELF(gen[2622]),
			.cell_state(gen[2622])
		); 

/******************* CELL 2623 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2623 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2527]),
			.N(gen[2528]),
			.NE(gen[2529]),

			.O(gen[2622]),
			.E(gen[2624]),

			.SO(gen[2717]),
			.S(gen[2718]),
			.SE(gen[2719]),

			.SELF(gen[2623]),
			.cell_state(gen[2623])
		); 

/******************* CELL 2624 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2624 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2528]),
			.N(gen[2529]),
			.NE(gen[2530]),

			.O(gen[2623]),
			.E(gen[2625]),

			.SO(gen[2718]),
			.S(gen[2719]),
			.SE(gen[2720]),

			.SELF(gen[2624]),
			.cell_state(gen[2624])
		); 

/******************* CELL 2625 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2625 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2529]),
			.N(gen[2530]),
			.NE(gen[2531]),

			.O(gen[2624]),
			.E(gen[2626]),

			.SO(gen[2719]),
			.S(gen[2720]),
			.SE(gen[2721]),

			.SELF(gen[2625]),
			.cell_state(gen[2625])
		); 

/******************* CELL 2626 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2626 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2530]),
			.N(gen[2531]),
			.NE(gen[2532]),

			.O(gen[2625]),
			.E(gen[2627]),

			.SO(gen[2720]),
			.S(gen[2721]),
			.SE(gen[2722]),

			.SELF(gen[2626]),
			.cell_state(gen[2626])
		); 

/******************* CELL 2627 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2627 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2531]),
			.N(gen[2532]),
			.NE(gen[2533]),

			.O(gen[2626]),
			.E(gen[2628]),

			.SO(gen[2721]),
			.S(gen[2722]),
			.SE(gen[2723]),

			.SELF(gen[2627]),
			.cell_state(gen[2627])
		); 

/******************* CELL 2628 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2628 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2532]),
			.N(gen[2533]),
			.NE(gen[2534]),

			.O(gen[2627]),
			.E(gen[2629]),

			.SO(gen[2722]),
			.S(gen[2723]),
			.SE(gen[2724]),

			.SELF(gen[2628]),
			.cell_state(gen[2628])
		); 

/******************* CELL 2629 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2629 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2533]),
			.N(gen[2534]),
			.NE(gen[2535]),

			.O(gen[2628]),
			.E(gen[2630]),

			.SO(gen[2723]),
			.S(gen[2724]),
			.SE(gen[2725]),

			.SELF(gen[2629]),
			.cell_state(gen[2629])
		); 

/******************* CELL 2630 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2630 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2534]),
			.N(gen[2535]),
			.NE(gen[2536]),

			.O(gen[2629]),
			.E(gen[2631]),

			.SO(gen[2724]),
			.S(gen[2725]),
			.SE(gen[2726]),

			.SELF(gen[2630]),
			.cell_state(gen[2630])
		); 

/******************* CELL 2631 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2631 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2535]),
			.N(gen[2536]),
			.NE(gen[2537]),

			.O(gen[2630]),
			.E(gen[2632]),

			.SO(gen[2725]),
			.S(gen[2726]),
			.SE(gen[2727]),

			.SELF(gen[2631]),
			.cell_state(gen[2631])
		); 

/******************* CELL 2632 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2632 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2536]),
			.N(gen[2537]),
			.NE(gen[2538]),

			.O(gen[2631]),
			.E(gen[2633]),

			.SO(gen[2726]),
			.S(gen[2727]),
			.SE(gen[2728]),

			.SELF(gen[2632]),
			.cell_state(gen[2632])
		); 

/******************* CELL 2633 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2633 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2537]),
			.N(gen[2538]),
			.NE(gen[2539]),

			.O(gen[2632]),
			.E(gen[2634]),

			.SO(gen[2727]),
			.S(gen[2728]),
			.SE(gen[2729]),

			.SELF(gen[2633]),
			.cell_state(gen[2633])
		); 

/******************* CELL 2634 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2634 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2538]),
			.N(gen[2539]),
			.NE(gen[2540]),

			.O(gen[2633]),
			.E(gen[2635]),

			.SO(gen[2728]),
			.S(gen[2729]),
			.SE(gen[2730]),

			.SELF(gen[2634]),
			.cell_state(gen[2634])
		); 

/******************* CELL 2635 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2635 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2539]),
			.N(gen[2540]),
			.NE(gen[2541]),

			.O(gen[2634]),
			.E(gen[2636]),

			.SO(gen[2729]),
			.S(gen[2730]),
			.SE(gen[2731]),

			.SELF(gen[2635]),
			.cell_state(gen[2635])
		); 

/******************* CELL 2636 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2636 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2540]),
			.N(gen[2541]),
			.NE(gen[2542]),

			.O(gen[2635]),
			.E(gen[2637]),

			.SO(gen[2730]),
			.S(gen[2731]),
			.SE(gen[2732]),

			.SELF(gen[2636]),
			.cell_state(gen[2636])
		); 

/******************* CELL 2637 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2637 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2541]),
			.N(gen[2542]),
			.NE(gen[2543]),

			.O(gen[2636]),
			.E(gen[2638]),

			.SO(gen[2731]),
			.S(gen[2732]),
			.SE(gen[2733]),

			.SELF(gen[2637]),
			.cell_state(gen[2637])
		); 

/******************* CELL 2638 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2638 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2542]),
			.N(gen[2543]),
			.NE(gen[2544]),

			.O(gen[2637]),
			.E(gen[2639]),

			.SO(gen[2732]),
			.S(gen[2733]),
			.SE(gen[2734]),

			.SELF(gen[2638]),
			.cell_state(gen[2638])
		); 

/******************* CELL 2639 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2639 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2543]),
			.N(gen[2544]),
			.NE(gen[2545]),

			.O(gen[2638]),
			.E(gen[2640]),

			.SO(gen[2733]),
			.S(gen[2734]),
			.SE(gen[2735]),

			.SELF(gen[2639]),
			.cell_state(gen[2639])
		); 

/******************* CELL 2640 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2640 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2544]),
			.N(gen[2545]),
			.NE(gen[2546]),

			.O(gen[2639]),
			.E(gen[2641]),

			.SO(gen[2734]),
			.S(gen[2735]),
			.SE(gen[2736]),

			.SELF(gen[2640]),
			.cell_state(gen[2640])
		); 

/******************* CELL 2641 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2641 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2545]),
			.N(gen[2546]),
			.NE(gen[2547]),

			.O(gen[2640]),
			.E(gen[2642]),

			.SO(gen[2735]),
			.S(gen[2736]),
			.SE(gen[2737]),

			.SELF(gen[2641]),
			.cell_state(gen[2641])
		); 

/******************* CELL 2642 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2642 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2546]),
			.N(gen[2547]),
			.NE(gen[2548]),

			.O(gen[2641]),
			.E(gen[2643]),

			.SO(gen[2736]),
			.S(gen[2737]),
			.SE(gen[2738]),

			.SELF(gen[2642]),
			.cell_state(gen[2642])
		); 

/******************* CELL 2643 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2643 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2547]),
			.N(gen[2548]),
			.NE(gen[2549]),

			.O(gen[2642]),
			.E(gen[2644]),

			.SO(gen[2737]),
			.S(gen[2738]),
			.SE(gen[2739]),

			.SELF(gen[2643]),
			.cell_state(gen[2643])
		); 

/******************* CELL 2644 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2644 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2548]),
			.N(gen[2549]),
			.NE(gen[2550]),

			.O(gen[2643]),
			.E(gen[2645]),

			.SO(gen[2738]),
			.S(gen[2739]),
			.SE(gen[2740]),

			.SELF(gen[2644]),
			.cell_state(gen[2644])
		); 

/******************* CELL 2645 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2645 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2549]),
			.N(gen[2550]),
			.NE(gen[2551]),

			.O(gen[2644]),
			.E(gen[2646]),

			.SO(gen[2739]),
			.S(gen[2740]),
			.SE(gen[2741]),

			.SELF(gen[2645]),
			.cell_state(gen[2645])
		); 

/******************* CELL 2646 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2646 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2550]),
			.N(gen[2551]),
			.NE(gen[2552]),

			.O(gen[2645]),
			.E(gen[2647]),

			.SO(gen[2740]),
			.S(gen[2741]),
			.SE(gen[2742]),

			.SELF(gen[2646]),
			.cell_state(gen[2646])
		); 

/******************* CELL 2647 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2647 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2551]),
			.N(gen[2552]),
			.NE(gen[2553]),

			.O(gen[2646]),
			.E(gen[2648]),

			.SO(gen[2741]),
			.S(gen[2742]),
			.SE(gen[2743]),

			.SELF(gen[2647]),
			.cell_state(gen[2647])
		); 

/******************* CELL 2648 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2648 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2552]),
			.N(gen[2553]),
			.NE(gen[2554]),

			.O(gen[2647]),
			.E(gen[2649]),

			.SO(gen[2742]),
			.S(gen[2743]),
			.SE(gen[2744]),

			.SELF(gen[2648]),
			.cell_state(gen[2648])
		); 

/******************* CELL 2649 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2649 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2553]),
			.N(gen[2554]),
			.NE(gen[2555]),

			.O(gen[2648]),
			.E(gen[2650]),

			.SO(gen[2743]),
			.S(gen[2744]),
			.SE(gen[2745]),

			.SELF(gen[2649]),
			.cell_state(gen[2649])
		); 

/******************* CELL 2650 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2650 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2554]),
			.N(gen[2555]),
			.NE(gen[2556]),

			.O(gen[2649]),
			.E(gen[2651]),

			.SO(gen[2744]),
			.S(gen[2745]),
			.SE(gen[2746]),

			.SELF(gen[2650]),
			.cell_state(gen[2650])
		); 

/******************* CELL 2651 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2651 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2555]),
			.N(gen[2556]),
			.NE(gen[2557]),

			.O(gen[2650]),
			.E(gen[2652]),

			.SO(gen[2745]),
			.S(gen[2746]),
			.SE(gen[2747]),

			.SELF(gen[2651]),
			.cell_state(gen[2651])
		); 

/******************* CELL 2652 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2652 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2556]),
			.N(gen[2557]),
			.NE(gen[2558]),

			.O(gen[2651]),
			.E(gen[2653]),

			.SO(gen[2746]),
			.S(gen[2747]),
			.SE(gen[2748]),

			.SELF(gen[2652]),
			.cell_state(gen[2652])
		); 

/******************* CELL 2653 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2653 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2557]),
			.N(gen[2558]),
			.NE(gen[2559]),

			.O(gen[2652]),
			.E(gen[2654]),

			.SO(gen[2747]),
			.S(gen[2748]),
			.SE(gen[2749]),

			.SELF(gen[2653]),
			.cell_state(gen[2653])
		); 

/******************* CELL 2654 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2654 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2558]),
			.N(gen[2559]),
			.NE(gen[2560]),

			.O(gen[2653]),
			.E(gen[2655]),

			.SO(gen[2748]),
			.S(gen[2749]),
			.SE(gen[2750]),

			.SELF(gen[2654]),
			.cell_state(gen[2654])
		); 

/******************* CELL 2655 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2655 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2559]),
			.N(gen[2560]),
			.NE(gen[2561]),

			.O(gen[2654]),
			.E(gen[2656]),

			.SO(gen[2749]),
			.S(gen[2750]),
			.SE(gen[2751]),

			.SELF(gen[2655]),
			.cell_state(gen[2655])
		); 

/******************* CELL 2656 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2656 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2560]),
			.N(gen[2561]),
			.NE(gen[2562]),

			.O(gen[2655]),
			.E(gen[2657]),

			.SO(gen[2750]),
			.S(gen[2751]),
			.SE(gen[2752]),

			.SELF(gen[2656]),
			.cell_state(gen[2656])
		); 

/******************* CELL 2657 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2657 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2561]),
			.N(gen[2562]),
			.NE(gen[2563]),

			.O(gen[2656]),
			.E(gen[2658]),

			.SO(gen[2751]),
			.S(gen[2752]),
			.SE(gen[2753]),

			.SELF(gen[2657]),
			.cell_state(gen[2657])
		); 

/******************* CELL 2658 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2658 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2562]),
			.N(gen[2563]),
			.NE(gen[2564]),

			.O(gen[2657]),
			.E(gen[2659]),

			.SO(gen[2752]),
			.S(gen[2753]),
			.SE(gen[2754]),

			.SELF(gen[2658]),
			.cell_state(gen[2658])
		); 

/******************* CELL 2659 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2659 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2563]),
			.N(gen[2564]),
			.NE(gen[2563]),

			.O(gen[2658]),
			.E(gen[2658]),

			.SO(gen[2753]),
			.S(gen[2754]),
			.SE(gen[2753]),

			.SELF(gen[2659]),
			.cell_state(gen[2659])
		); 

/******************* CELL 2660 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2660 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2566]),
			.N(gen[2565]),
			.NE(gen[2566]),

			.O(gen[2661]),
			.E(gen[2661]),

			.SO(gen[2756]),
			.S(gen[2755]),
			.SE(gen[2756]),

			.SELF(gen[2660]),
			.cell_state(gen[2660])
		); 

/******************* CELL 2661 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2661 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2565]),
			.N(gen[2566]),
			.NE(gen[2567]),

			.O(gen[2660]),
			.E(gen[2662]),

			.SO(gen[2755]),
			.S(gen[2756]),
			.SE(gen[2757]),

			.SELF(gen[2661]),
			.cell_state(gen[2661])
		); 

/******************* CELL 2662 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2662 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2566]),
			.N(gen[2567]),
			.NE(gen[2568]),

			.O(gen[2661]),
			.E(gen[2663]),

			.SO(gen[2756]),
			.S(gen[2757]),
			.SE(gen[2758]),

			.SELF(gen[2662]),
			.cell_state(gen[2662])
		); 

/******************* CELL 2663 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2663 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2567]),
			.N(gen[2568]),
			.NE(gen[2569]),

			.O(gen[2662]),
			.E(gen[2664]),

			.SO(gen[2757]),
			.S(gen[2758]),
			.SE(gen[2759]),

			.SELF(gen[2663]),
			.cell_state(gen[2663])
		); 

/******************* CELL 2664 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2664 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2568]),
			.N(gen[2569]),
			.NE(gen[2570]),

			.O(gen[2663]),
			.E(gen[2665]),

			.SO(gen[2758]),
			.S(gen[2759]),
			.SE(gen[2760]),

			.SELF(gen[2664]),
			.cell_state(gen[2664])
		); 

/******************* CELL 2665 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2665 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2569]),
			.N(gen[2570]),
			.NE(gen[2571]),

			.O(gen[2664]),
			.E(gen[2666]),

			.SO(gen[2759]),
			.S(gen[2760]),
			.SE(gen[2761]),

			.SELF(gen[2665]),
			.cell_state(gen[2665])
		); 

/******************* CELL 2666 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2666 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2570]),
			.N(gen[2571]),
			.NE(gen[2572]),

			.O(gen[2665]),
			.E(gen[2667]),

			.SO(gen[2760]),
			.S(gen[2761]),
			.SE(gen[2762]),

			.SELF(gen[2666]),
			.cell_state(gen[2666])
		); 

/******************* CELL 2667 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2667 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2571]),
			.N(gen[2572]),
			.NE(gen[2573]),

			.O(gen[2666]),
			.E(gen[2668]),

			.SO(gen[2761]),
			.S(gen[2762]),
			.SE(gen[2763]),

			.SELF(gen[2667]),
			.cell_state(gen[2667])
		); 

/******************* CELL 2668 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2668 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2572]),
			.N(gen[2573]),
			.NE(gen[2574]),

			.O(gen[2667]),
			.E(gen[2669]),

			.SO(gen[2762]),
			.S(gen[2763]),
			.SE(gen[2764]),

			.SELF(gen[2668]),
			.cell_state(gen[2668])
		); 

/******************* CELL 2669 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2669 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2573]),
			.N(gen[2574]),
			.NE(gen[2575]),

			.O(gen[2668]),
			.E(gen[2670]),

			.SO(gen[2763]),
			.S(gen[2764]),
			.SE(gen[2765]),

			.SELF(gen[2669]),
			.cell_state(gen[2669])
		); 

/******************* CELL 2670 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2670 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2574]),
			.N(gen[2575]),
			.NE(gen[2576]),

			.O(gen[2669]),
			.E(gen[2671]),

			.SO(gen[2764]),
			.S(gen[2765]),
			.SE(gen[2766]),

			.SELF(gen[2670]),
			.cell_state(gen[2670])
		); 

/******************* CELL 2671 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2671 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2575]),
			.N(gen[2576]),
			.NE(gen[2577]),

			.O(gen[2670]),
			.E(gen[2672]),

			.SO(gen[2765]),
			.S(gen[2766]),
			.SE(gen[2767]),

			.SELF(gen[2671]),
			.cell_state(gen[2671])
		); 

/******************* CELL 2672 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2672 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2576]),
			.N(gen[2577]),
			.NE(gen[2578]),

			.O(gen[2671]),
			.E(gen[2673]),

			.SO(gen[2766]),
			.S(gen[2767]),
			.SE(gen[2768]),

			.SELF(gen[2672]),
			.cell_state(gen[2672])
		); 

/******************* CELL 2673 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2673 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2577]),
			.N(gen[2578]),
			.NE(gen[2579]),

			.O(gen[2672]),
			.E(gen[2674]),

			.SO(gen[2767]),
			.S(gen[2768]),
			.SE(gen[2769]),

			.SELF(gen[2673]),
			.cell_state(gen[2673])
		); 

/******************* CELL 2674 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2674 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2578]),
			.N(gen[2579]),
			.NE(gen[2580]),

			.O(gen[2673]),
			.E(gen[2675]),

			.SO(gen[2768]),
			.S(gen[2769]),
			.SE(gen[2770]),

			.SELF(gen[2674]),
			.cell_state(gen[2674])
		); 

/******************* CELL 2675 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2675 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2579]),
			.N(gen[2580]),
			.NE(gen[2581]),

			.O(gen[2674]),
			.E(gen[2676]),

			.SO(gen[2769]),
			.S(gen[2770]),
			.SE(gen[2771]),

			.SELF(gen[2675]),
			.cell_state(gen[2675])
		); 

/******************* CELL 2676 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2676 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2580]),
			.N(gen[2581]),
			.NE(gen[2582]),

			.O(gen[2675]),
			.E(gen[2677]),

			.SO(gen[2770]),
			.S(gen[2771]),
			.SE(gen[2772]),

			.SELF(gen[2676]),
			.cell_state(gen[2676])
		); 

/******************* CELL 2677 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2677 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2581]),
			.N(gen[2582]),
			.NE(gen[2583]),

			.O(gen[2676]),
			.E(gen[2678]),

			.SO(gen[2771]),
			.S(gen[2772]),
			.SE(gen[2773]),

			.SELF(gen[2677]),
			.cell_state(gen[2677])
		); 

/******************* CELL 2678 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2678 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2582]),
			.N(gen[2583]),
			.NE(gen[2584]),

			.O(gen[2677]),
			.E(gen[2679]),

			.SO(gen[2772]),
			.S(gen[2773]),
			.SE(gen[2774]),

			.SELF(gen[2678]),
			.cell_state(gen[2678])
		); 

/******************* CELL 2679 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2679 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2583]),
			.N(gen[2584]),
			.NE(gen[2585]),

			.O(gen[2678]),
			.E(gen[2680]),

			.SO(gen[2773]),
			.S(gen[2774]),
			.SE(gen[2775]),

			.SELF(gen[2679]),
			.cell_state(gen[2679])
		); 

/******************* CELL 2680 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2680 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2584]),
			.N(gen[2585]),
			.NE(gen[2586]),

			.O(gen[2679]),
			.E(gen[2681]),

			.SO(gen[2774]),
			.S(gen[2775]),
			.SE(gen[2776]),

			.SELF(gen[2680]),
			.cell_state(gen[2680])
		); 

/******************* CELL 2681 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2681 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2585]),
			.N(gen[2586]),
			.NE(gen[2587]),

			.O(gen[2680]),
			.E(gen[2682]),

			.SO(gen[2775]),
			.S(gen[2776]),
			.SE(gen[2777]),

			.SELF(gen[2681]),
			.cell_state(gen[2681])
		); 

/******************* CELL 2682 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2682 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2586]),
			.N(gen[2587]),
			.NE(gen[2588]),

			.O(gen[2681]),
			.E(gen[2683]),

			.SO(gen[2776]),
			.S(gen[2777]),
			.SE(gen[2778]),

			.SELF(gen[2682]),
			.cell_state(gen[2682])
		); 

/******************* CELL 2683 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2683 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2587]),
			.N(gen[2588]),
			.NE(gen[2589]),

			.O(gen[2682]),
			.E(gen[2684]),

			.SO(gen[2777]),
			.S(gen[2778]),
			.SE(gen[2779]),

			.SELF(gen[2683]),
			.cell_state(gen[2683])
		); 

/******************* CELL 2684 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2684 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2588]),
			.N(gen[2589]),
			.NE(gen[2590]),

			.O(gen[2683]),
			.E(gen[2685]),

			.SO(gen[2778]),
			.S(gen[2779]),
			.SE(gen[2780]),

			.SELF(gen[2684]),
			.cell_state(gen[2684])
		); 

/******************* CELL 2685 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2685 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2589]),
			.N(gen[2590]),
			.NE(gen[2591]),

			.O(gen[2684]),
			.E(gen[2686]),

			.SO(gen[2779]),
			.S(gen[2780]),
			.SE(gen[2781]),

			.SELF(gen[2685]),
			.cell_state(gen[2685])
		); 

/******************* CELL 2686 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2686 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2590]),
			.N(gen[2591]),
			.NE(gen[2592]),

			.O(gen[2685]),
			.E(gen[2687]),

			.SO(gen[2780]),
			.S(gen[2781]),
			.SE(gen[2782]),

			.SELF(gen[2686]),
			.cell_state(gen[2686])
		); 

/******************* CELL 2687 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2687 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2591]),
			.N(gen[2592]),
			.NE(gen[2593]),

			.O(gen[2686]),
			.E(gen[2688]),

			.SO(gen[2781]),
			.S(gen[2782]),
			.SE(gen[2783]),

			.SELF(gen[2687]),
			.cell_state(gen[2687])
		); 

/******************* CELL 2688 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2688 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2592]),
			.N(gen[2593]),
			.NE(gen[2594]),

			.O(gen[2687]),
			.E(gen[2689]),

			.SO(gen[2782]),
			.S(gen[2783]),
			.SE(gen[2784]),

			.SELF(gen[2688]),
			.cell_state(gen[2688])
		); 

/******************* CELL 2689 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2689 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2593]),
			.N(gen[2594]),
			.NE(gen[2595]),

			.O(gen[2688]),
			.E(gen[2690]),

			.SO(gen[2783]),
			.S(gen[2784]),
			.SE(gen[2785]),

			.SELF(gen[2689]),
			.cell_state(gen[2689])
		); 

/******************* CELL 2690 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2690 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2594]),
			.N(gen[2595]),
			.NE(gen[2596]),

			.O(gen[2689]),
			.E(gen[2691]),

			.SO(gen[2784]),
			.S(gen[2785]),
			.SE(gen[2786]),

			.SELF(gen[2690]),
			.cell_state(gen[2690])
		); 

/******************* CELL 2691 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2691 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2595]),
			.N(gen[2596]),
			.NE(gen[2597]),

			.O(gen[2690]),
			.E(gen[2692]),

			.SO(gen[2785]),
			.S(gen[2786]),
			.SE(gen[2787]),

			.SELF(gen[2691]),
			.cell_state(gen[2691])
		); 

/******************* CELL 2692 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2692 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2596]),
			.N(gen[2597]),
			.NE(gen[2598]),

			.O(gen[2691]),
			.E(gen[2693]),

			.SO(gen[2786]),
			.S(gen[2787]),
			.SE(gen[2788]),

			.SELF(gen[2692]),
			.cell_state(gen[2692])
		); 

/******************* CELL 2693 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2693 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2597]),
			.N(gen[2598]),
			.NE(gen[2599]),

			.O(gen[2692]),
			.E(gen[2694]),

			.SO(gen[2787]),
			.S(gen[2788]),
			.SE(gen[2789]),

			.SELF(gen[2693]),
			.cell_state(gen[2693])
		); 

/******************* CELL 2694 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2694 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2598]),
			.N(gen[2599]),
			.NE(gen[2600]),

			.O(gen[2693]),
			.E(gen[2695]),

			.SO(gen[2788]),
			.S(gen[2789]),
			.SE(gen[2790]),

			.SELF(gen[2694]),
			.cell_state(gen[2694])
		); 

/******************* CELL 2695 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2695 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2599]),
			.N(gen[2600]),
			.NE(gen[2601]),

			.O(gen[2694]),
			.E(gen[2696]),

			.SO(gen[2789]),
			.S(gen[2790]),
			.SE(gen[2791]),

			.SELF(gen[2695]),
			.cell_state(gen[2695])
		); 

/******************* CELL 2696 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2696 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2600]),
			.N(gen[2601]),
			.NE(gen[2602]),

			.O(gen[2695]),
			.E(gen[2697]),

			.SO(gen[2790]),
			.S(gen[2791]),
			.SE(gen[2792]),

			.SELF(gen[2696]),
			.cell_state(gen[2696])
		); 

/******************* CELL 2697 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2697 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2601]),
			.N(gen[2602]),
			.NE(gen[2603]),

			.O(gen[2696]),
			.E(gen[2698]),

			.SO(gen[2791]),
			.S(gen[2792]),
			.SE(gen[2793]),

			.SELF(gen[2697]),
			.cell_state(gen[2697])
		); 

/******************* CELL 2698 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2698 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2602]),
			.N(gen[2603]),
			.NE(gen[2604]),

			.O(gen[2697]),
			.E(gen[2699]),

			.SO(gen[2792]),
			.S(gen[2793]),
			.SE(gen[2794]),

			.SELF(gen[2698]),
			.cell_state(gen[2698])
		); 

/******************* CELL 2699 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2699 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2603]),
			.N(gen[2604]),
			.NE(gen[2605]),

			.O(gen[2698]),
			.E(gen[2700]),

			.SO(gen[2793]),
			.S(gen[2794]),
			.SE(gen[2795]),

			.SELF(gen[2699]),
			.cell_state(gen[2699])
		); 

/******************* CELL 2700 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2700 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2604]),
			.N(gen[2605]),
			.NE(gen[2606]),

			.O(gen[2699]),
			.E(gen[2701]),

			.SO(gen[2794]),
			.S(gen[2795]),
			.SE(gen[2796]),

			.SELF(gen[2700]),
			.cell_state(gen[2700])
		); 

/******************* CELL 2701 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2701 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2605]),
			.N(gen[2606]),
			.NE(gen[2607]),

			.O(gen[2700]),
			.E(gen[2702]),

			.SO(gen[2795]),
			.S(gen[2796]),
			.SE(gen[2797]),

			.SELF(gen[2701]),
			.cell_state(gen[2701])
		); 

/******************* CELL 2702 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2702 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2606]),
			.N(gen[2607]),
			.NE(gen[2608]),

			.O(gen[2701]),
			.E(gen[2703]),

			.SO(gen[2796]),
			.S(gen[2797]),
			.SE(gen[2798]),

			.SELF(gen[2702]),
			.cell_state(gen[2702])
		); 

/******************* CELL 2703 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2703 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2607]),
			.N(gen[2608]),
			.NE(gen[2609]),

			.O(gen[2702]),
			.E(gen[2704]),

			.SO(gen[2797]),
			.S(gen[2798]),
			.SE(gen[2799]),

			.SELF(gen[2703]),
			.cell_state(gen[2703])
		); 

/******************* CELL 2704 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2704 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2608]),
			.N(gen[2609]),
			.NE(gen[2610]),

			.O(gen[2703]),
			.E(gen[2705]),

			.SO(gen[2798]),
			.S(gen[2799]),
			.SE(gen[2800]),

			.SELF(gen[2704]),
			.cell_state(gen[2704])
		); 

/******************* CELL 2705 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2705 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2609]),
			.N(gen[2610]),
			.NE(gen[2611]),

			.O(gen[2704]),
			.E(gen[2706]),

			.SO(gen[2799]),
			.S(gen[2800]),
			.SE(gen[2801]),

			.SELF(gen[2705]),
			.cell_state(gen[2705])
		); 

/******************* CELL 2706 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2706 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2610]),
			.N(gen[2611]),
			.NE(gen[2612]),

			.O(gen[2705]),
			.E(gen[2707]),

			.SO(gen[2800]),
			.S(gen[2801]),
			.SE(gen[2802]),

			.SELF(gen[2706]),
			.cell_state(gen[2706])
		); 

/******************* CELL 2707 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2707 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2611]),
			.N(gen[2612]),
			.NE(gen[2613]),

			.O(gen[2706]),
			.E(gen[2708]),

			.SO(gen[2801]),
			.S(gen[2802]),
			.SE(gen[2803]),

			.SELF(gen[2707]),
			.cell_state(gen[2707])
		); 

/******************* CELL 2708 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2708 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2612]),
			.N(gen[2613]),
			.NE(gen[2614]),

			.O(gen[2707]),
			.E(gen[2709]),

			.SO(gen[2802]),
			.S(gen[2803]),
			.SE(gen[2804]),

			.SELF(gen[2708]),
			.cell_state(gen[2708])
		); 

/******************* CELL 2709 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2709 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2613]),
			.N(gen[2614]),
			.NE(gen[2615]),

			.O(gen[2708]),
			.E(gen[2710]),

			.SO(gen[2803]),
			.S(gen[2804]),
			.SE(gen[2805]),

			.SELF(gen[2709]),
			.cell_state(gen[2709])
		); 

/******************* CELL 2710 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2710 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2614]),
			.N(gen[2615]),
			.NE(gen[2616]),

			.O(gen[2709]),
			.E(gen[2711]),

			.SO(gen[2804]),
			.S(gen[2805]),
			.SE(gen[2806]),

			.SELF(gen[2710]),
			.cell_state(gen[2710])
		); 

/******************* CELL 2711 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2711 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2615]),
			.N(gen[2616]),
			.NE(gen[2617]),

			.O(gen[2710]),
			.E(gen[2712]),

			.SO(gen[2805]),
			.S(gen[2806]),
			.SE(gen[2807]),

			.SELF(gen[2711]),
			.cell_state(gen[2711])
		); 

/******************* CELL 2712 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2712 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2616]),
			.N(gen[2617]),
			.NE(gen[2618]),

			.O(gen[2711]),
			.E(gen[2713]),

			.SO(gen[2806]),
			.S(gen[2807]),
			.SE(gen[2808]),

			.SELF(gen[2712]),
			.cell_state(gen[2712])
		); 

/******************* CELL 2713 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2713 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2617]),
			.N(gen[2618]),
			.NE(gen[2619]),

			.O(gen[2712]),
			.E(gen[2714]),

			.SO(gen[2807]),
			.S(gen[2808]),
			.SE(gen[2809]),

			.SELF(gen[2713]),
			.cell_state(gen[2713])
		); 

/******************* CELL 2714 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2714 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2618]),
			.N(gen[2619]),
			.NE(gen[2620]),

			.O(gen[2713]),
			.E(gen[2715]),

			.SO(gen[2808]),
			.S(gen[2809]),
			.SE(gen[2810]),

			.SELF(gen[2714]),
			.cell_state(gen[2714])
		); 

/******************* CELL 2715 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2715 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2619]),
			.N(gen[2620]),
			.NE(gen[2621]),

			.O(gen[2714]),
			.E(gen[2716]),

			.SO(gen[2809]),
			.S(gen[2810]),
			.SE(gen[2811]),

			.SELF(gen[2715]),
			.cell_state(gen[2715])
		); 

/******************* CELL 2716 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2716 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2620]),
			.N(gen[2621]),
			.NE(gen[2622]),

			.O(gen[2715]),
			.E(gen[2717]),

			.SO(gen[2810]),
			.S(gen[2811]),
			.SE(gen[2812]),

			.SELF(gen[2716]),
			.cell_state(gen[2716])
		); 

/******************* CELL 2717 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2717 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2621]),
			.N(gen[2622]),
			.NE(gen[2623]),

			.O(gen[2716]),
			.E(gen[2718]),

			.SO(gen[2811]),
			.S(gen[2812]),
			.SE(gen[2813]),

			.SELF(gen[2717]),
			.cell_state(gen[2717])
		); 

/******************* CELL 2718 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2718 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2622]),
			.N(gen[2623]),
			.NE(gen[2624]),

			.O(gen[2717]),
			.E(gen[2719]),

			.SO(gen[2812]),
			.S(gen[2813]),
			.SE(gen[2814]),

			.SELF(gen[2718]),
			.cell_state(gen[2718])
		); 

/******************* CELL 2719 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2719 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2623]),
			.N(gen[2624]),
			.NE(gen[2625]),

			.O(gen[2718]),
			.E(gen[2720]),

			.SO(gen[2813]),
			.S(gen[2814]),
			.SE(gen[2815]),

			.SELF(gen[2719]),
			.cell_state(gen[2719])
		); 

/******************* CELL 2720 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2720 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2624]),
			.N(gen[2625]),
			.NE(gen[2626]),

			.O(gen[2719]),
			.E(gen[2721]),

			.SO(gen[2814]),
			.S(gen[2815]),
			.SE(gen[2816]),

			.SELF(gen[2720]),
			.cell_state(gen[2720])
		); 

/******************* CELL 2721 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2721 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2625]),
			.N(gen[2626]),
			.NE(gen[2627]),

			.O(gen[2720]),
			.E(gen[2722]),

			.SO(gen[2815]),
			.S(gen[2816]),
			.SE(gen[2817]),

			.SELF(gen[2721]),
			.cell_state(gen[2721])
		); 

/******************* CELL 2722 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2722 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2626]),
			.N(gen[2627]),
			.NE(gen[2628]),

			.O(gen[2721]),
			.E(gen[2723]),

			.SO(gen[2816]),
			.S(gen[2817]),
			.SE(gen[2818]),

			.SELF(gen[2722]),
			.cell_state(gen[2722])
		); 

/******************* CELL 2723 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2723 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2627]),
			.N(gen[2628]),
			.NE(gen[2629]),

			.O(gen[2722]),
			.E(gen[2724]),

			.SO(gen[2817]),
			.S(gen[2818]),
			.SE(gen[2819]),

			.SELF(gen[2723]),
			.cell_state(gen[2723])
		); 

/******************* CELL 2724 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2724 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2628]),
			.N(gen[2629]),
			.NE(gen[2630]),

			.O(gen[2723]),
			.E(gen[2725]),

			.SO(gen[2818]),
			.S(gen[2819]),
			.SE(gen[2820]),

			.SELF(gen[2724]),
			.cell_state(gen[2724])
		); 

/******************* CELL 2725 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2725 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2629]),
			.N(gen[2630]),
			.NE(gen[2631]),

			.O(gen[2724]),
			.E(gen[2726]),

			.SO(gen[2819]),
			.S(gen[2820]),
			.SE(gen[2821]),

			.SELF(gen[2725]),
			.cell_state(gen[2725])
		); 

/******************* CELL 2726 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2726 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2630]),
			.N(gen[2631]),
			.NE(gen[2632]),

			.O(gen[2725]),
			.E(gen[2727]),

			.SO(gen[2820]),
			.S(gen[2821]),
			.SE(gen[2822]),

			.SELF(gen[2726]),
			.cell_state(gen[2726])
		); 

/******************* CELL 2727 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2727 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2631]),
			.N(gen[2632]),
			.NE(gen[2633]),

			.O(gen[2726]),
			.E(gen[2728]),

			.SO(gen[2821]),
			.S(gen[2822]),
			.SE(gen[2823]),

			.SELF(gen[2727]),
			.cell_state(gen[2727])
		); 

/******************* CELL 2728 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2728 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2632]),
			.N(gen[2633]),
			.NE(gen[2634]),

			.O(gen[2727]),
			.E(gen[2729]),

			.SO(gen[2822]),
			.S(gen[2823]),
			.SE(gen[2824]),

			.SELF(gen[2728]),
			.cell_state(gen[2728])
		); 

/******************* CELL 2729 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2729 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2633]),
			.N(gen[2634]),
			.NE(gen[2635]),

			.O(gen[2728]),
			.E(gen[2730]),

			.SO(gen[2823]),
			.S(gen[2824]),
			.SE(gen[2825]),

			.SELF(gen[2729]),
			.cell_state(gen[2729])
		); 

/******************* CELL 2730 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2730 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2634]),
			.N(gen[2635]),
			.NE(gen[2636]),

			.O(gen[2729]),
			.E(gen[2731]),

			.SO(gen[2824]),
			.S(gen[2825]),
			.SE(gen[2826]),

			.SELF(gen[2730]),
			.cell_state(gen[2730])
		); 

/******************* CELL 2731 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2731 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2635]),
			.N(gen[2636]),
			.NE(gen[2637]),

			.O(gen[2730]),
			.E(gen[2732]),

			.SO(gen[2825]),
			.S(gen[2826]),
			.SE(gen[2827]),

			.SELF(gen[2731]),
			.cell_state(gen[2731])
		); 

/******************* CELL 2732 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2732 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2636]),
			.N(gen[2637]),
			.NE(gen[2638]),

			.O(gen[2731]),
			.E(gen[2733]),

			.SO(gen[2826]),
			.S(gen[2827]),
			.SE(gen[2828]),

			.SELF(gen[2732]),
			.cell_state(gen[2732])
		); 

/******************* CELL 2733 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2733 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2637]),
			.N(gen[2638]),
			.NE(gen[2639]),

			.O(gen[2732]),
			.E(gen[2734]),

			.SO(gen[2827]),
			.S(gen[2828]),
			.SE(gen[2829]),

			.SELF(gen[2733]),
			.cell_state(gen[2733])
		); 

/******************* CELL 2734 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2734 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2638]),
			.N(gen[2639]),
			.NE(gen[2640]),

			.O(gen[2733]),
			.E(gen[2735]),

			.SO(gen[2828]),
			.S(gen[2829]),
			.SE(gen[2830]),

			.SELF(gen[2734]),
			.cell_state(gen[2734])
		); 

/******************* CELL 2735 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2735 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2639]),
			.N(gen[2640]),
			.NE(gen[2641]),

			.O(gen[2734]),
			.E(gen[2736]),

			.SO(gen[2829]),
			.S(gen[2830]),
			.SE(gen[2831]),

			.SELF(gen[2735]),
			.cell_state(gen[2735])
		); 

/******************* CELL 2736 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2736 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2640]),
			.N(gen[2641]),
			.NE(gen[2642]),

			.O(gen[2735]),
			.E(gen[2737]),

			.SO(gen[2830]),
			.S(gen[2831]),
			.SE(gen[2832]),

			.SELF(gen[2736]),
			.cell_state(gen[2736])
		); 

/******************* CELL 2737 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2737 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2641]),
			.N(gen[2642]),
			.NE(gen[2643]),

			.O(gen[2736]),
			.E(gen[2738]),

			.SO(gen[2831]),
			.S(gen[2832]),
			.SE(gen[2833]),

			.SELF(gen[2737]),
			.cell_state(gen[2737])
		); 

/******************* CELL 2738 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2738 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2642]),
			.N(gen[2643]),
			.NE(gen[2644]),

			.O(gen[2737]),
			.E(gen[2739]),

			.SO(gen[2832]),
			.S(gen[2833]),
			.SE(gen[2834]),

			.SELF(gen[2738]),
			.cell_state(gen[2738])
		); 

/******************* CELL 2739 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2739 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2643]),
			.N(gen[2644]),
			.NE(gen[2645]),

			.O(gen[2738]),
			.E(gen[2740]),

			.SO(gen[2833]),
			.S(gen[2834]),
			.SE(gen[2835]),

			.SELF(gen[2739]),
			.cell_state(gen[2739])
		); 

/******************* CELL 2740 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2740 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2644]),
			.N(gen[2645]),
			.NE(gen[2646]),

			.O(gen[2739]),
			.E(gen[2741]),

			.SO(gen[2834]),
			.S(gen[2835]),
			.SE(gen[2836]),

			.SELF(gen[2740]),
			.cell_state(gen[2740])
		); 

/******************* CELL 2741 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2741 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2645]),
			.N(gen[2646]),
			.NE(gen[2647]),

			.O(gen[2740]),
			.E(gen[2742]),

			.SO(gen[2835]),
			.S(gen[2836]),
			.SE(gen[2837]),

			.SELF(gen[2741]),
			.cell_state(gen[2741])
		); 

/******************* CELL 2742 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2742 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2646]),
			.N(gen[2647]),
			.NE(gen[2648]),

			.O(gen[2741]),
			.E(gen[2743]),

			.SO(gen[2836]),
			.S(gen[2837]),
			.SE(gen[2838]),

			.SELF(gen[2742]),
			.cell_state(gen[2742])
		); 

/******************* CELL 2743 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2743 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2647]),
			.N(gen[2648]),
			.NE(gen[2649]),

			.O(gen[2742]),
			.E(gen[2744]),

			.SO(gen[2837]),
			.S(gen[2838]),
			.SE(gen[2839]),

			.SELF(gen[2743]),
			.cell_state(gen[2743])
		); 

/******************* CELL 2744 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2744 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2648]),
			.N(gen[2649]),
			.NE(gen[2650]),

			.O(gen[2743]),
			.E(gen[2745]),

			.SO(gen[2838]),
			.S(gen[2839]),
			.SE(gen[2840]),

			.SELF(gen[2744]),
			.cell_state(gen[2744])
		); 

/******************* CELL 2745 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2745 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2649]),
			.N(gen[2650]),
			.NE(gen[2651]),

			.O(gen[2744]),
			.E(gen[2746]),

			.SO(gen[2839]),
			.S(gen[2840]),
			.SE(gen[2841]),

			.SELF(gen[2745]),
			.cell_state(gen[2745])
		); 

/******************* CELL 2746 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2746 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2650]),
			.N(gen[2651]),
			.NE(gen[2652]),

			.O(gen[2745]),
			.E(gen[2747]),

			.SO(gen[2840]),
			.S(gen[2841]),
			.SE(gen[2842]),

			.SELF(gen[2746]),
			.cell_state(gen[2746])
		); 

/******************* CELL 2747 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2747 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2651]),
			.N(gen[2652]),
			.NE(gen[2653]),

			.O(gen[2746]),
			.E(gen[2748]),

			.SO(gen[2841]),
			.S(gen[2842]),
			.SE(gen[2843]),

			.SELF(gen[2747]),
			.cell_state(gen[2747])
		); 

/******************* CELL 2748 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2748 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2652]),
			.N(gen[2653]),
			.NE(gen[2654]),

			.O(gen[2747]),
			.E(gen[2749]),

			.SO(gen[2842]),
			.S(gen[2843]),
			.SE(gen[2844]),

			.SELF(gen[2748]),
			.cell_state(gen[2748])
		); 

/******************* CELL 2749 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2749 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2653]),
			.N(gen[2654]),
			.NE(gen[2655]),

			.O(gen[2748]),
			.E(gen[2750]),

			.SO(gen[2843]),
			.S(gen[2844]),
			.SE(gen[2845]),

			.SELF(gen[2749]),
			.cell_state(gen[2749])
		); 

/******************* CELL 2750 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2750 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2654]),
			.N(gen[2655]),
			.NE(gen[2656]),

			.O(gen[2749]),
			.E(gen[2751]),

			.SO(gen[2844]),
			.S(gen[2845]),
			.SE(gen[2846]),

			.SELF(gen[2750]),
			.cell_state(gen[2750])
		); 

/******************* CELL 2751 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2751 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2655]),
			.N(gen[2656]),
			.NE(gen[2657]),

			.O(gen[2750]),
			.E(gen[2752]),

			.SO(gen[2845]),
			.S(gen[2846]),
			.SE(gen[2847]),

			.SELF(gen[2751]),
			.cell_state(gen[2751])
		); 

/******************* CELL 2752 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2752 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2656]),
			.N(gen[2657]),
			.NE(gen[2658]),

			.O(gen[2751]),
			.E(gen[2753]),

			.SO(gen[2846]),
			.S(gen[2847]),
			.SE(gen[2848]),

			.SELF(gen[2752]),
			.cell_state(gen[2752])
		); 

/******************* CELL 2753 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2753 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2657]),
			.N(gen[2658]),
			.NE(gen[2659]),

			.O(gen[2752]),
			.E(gen[2754]),

			.SO(gen[2847]),
			.S(gen[2848]),
			.SE(gen[2849]),

			.SELF(gen[2753]),
			.cell_state(gen[2753])
		); 

/******************* CELL 2754 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2754 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2658]),
			.N(gen[2659]),
			.NE(gen[2658]),

			.O(gen[2753]),
			.E(gen[2753]),

			.SO(gen[2848]),
			.S(gen[2849]),
			.SE(gen[2848]),

			.SELF(gen[2754]),
			.cell_state(gen[2754])
		); 

/******************* CELL 2755 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2755 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2661]),
			.N(gen[2660]),
			.NE(gen[2661]),

			.O(gen[2756]),
			.E(gen[2756]),

			.SO(gen[2851]),
			.S(gen[2850]),
			.SE(gen[2851]),

			.SELF(gen[2755]),
			.cell_state(gen[2755])
		); 

/******************* CELL 2756 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2756 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2660]),
			.N(gen[2661]),
			.NE(gen[2662]),

			.O(gen[2755]),
			.E(gen[2757]),

			.SO(gen[2850]),
			.S(gen[2851]),
			.SE(gen[2852]),

			.SELF(gen[2756]),
			.cell_state(gen[2756])
		); 

/******************* CELL 2757 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2757 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2661]),
			.N(gen[2662]),
			.NE(gen[2663]),

			.O(gen[2756]),
			.E(gen[2758]),

			.SO(gen[2851]),
			.S(gen[2852]),
			.SE(gen[2853]),

			.SELF(gen[2757]),
			.cell_state(gen[2757])
		); 

/******************* CELL 2758 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2758 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2662]),
			.N(gen[2663]),
			.NE(gen[2664]),

			.O(gen[2757]),
			.E(gen[2759]),

			.SO(gen[2852]),
			.S(gen[2853]),
			.SE(gen[2854]),

			.SELF(gen[2758]),
			.cell_state(gen[2758])
		); 

/******************* CELL 2759 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2759 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2663]),
			.N(gen[2664]),
			.NE(gen[2665]),

			.O(gen[2758]),
			.E(gen[2760]),

			.SO(gen[2853]),
			.S(gen[2854]),
			.SE(gen[2855]),

			.SELF(gen[2759]),
			.cell_state(gen[2759])
		); 

/******************* CELL 2760 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2760 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2664]),
			.N(gen[2665]),
			.NE(gen[2666]),

			.O(gen[2759]),
			.E(gen[2761]),

			.SO(gen[2854]),
			.S(gen[2855]),
			.SE(gen[2856]),

			.SELF(gen[2760]),
			.cell_state(gen[2760])
		); 

/******************* CELL 2761 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2761 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2665]),
			.N(gen[2666]),
			.NE(gen[2667]),

			.O(gen[2760]),
			.E(gen[2762]),

			.SO(gen[2855]),
			.S(gen[2856]),
			.SE(gen[2857]),

			.SELF(gen[2761]),
			.cell_state(gen[2761])
		); 

/******************* CELL 2762 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2762 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2666]),
			.N(gen[2667]),
			.NE(gen[2668]),

			.O(gen[2761]),
			.E(gen[2763]),

			.SO(gen[2856]),
			.S(gen[2857]),
			.SE(gen[2858]),

			.SELF(gen[2762]),
			.cell_state(gen[2762])
		); 

/******************* CELL 2763 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2763 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2667]),
			.N(gen[2668]),
			.NE(gen[2669]),

			.O(gen[2762]),
			.E(gen[2764]),

			.SO(gen[2857]),
			.S(gen[2858]),
			.SE(gen[2859]),

			.SELF(gen[2763]),
			.cell_state(gen[2763])
		); 

/******************* CELL 2764 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2764 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2668]),
			.N(gen[2669]),
			.NE(gen[2670]),

			.O(gen[2763]),
			.E(gen[2765]),

			.SO(gen[2858]),
			.S(gen[2859]),
			.SE(gen[2860]),

			.SELF(gen[2764]),
			.cell_state(gen[2764])
		); 

/******************* CELL 2765 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2765 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2669]),
			.N(gen[2670]),
			.NE(gen[2671]),

			.O(gen[2764]),
			.E(gen[2766]),

			.SO(gen[2859]),
			.S(gen[2860]),
			.SE(gen[2861]),

			.SELF(gen[2765]),
			.cell_state(gen[2765])
		); 

/******************* CELL 2766 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2766 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2670]),
			.N(gen[2671]),
			.NE(gen[2672]),

			.O(gen[2765]),
			.E(gen[2767]),

			.SO(gen[2860]),
			.S(gen[2861]),
			.SE(gen[2862]),

			.SELF(gen[2766]),
			.cell_state(gen[2766])
		); 

/******************* CELL 2767 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2767 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2671]),
			.N(gen[2672]),
			.NE(gen[2673]),

			.O(gen[2766]),
			.E(gen[2768]),

			.SO(gen[2861]),
			.S(gen[2862]),
			.SE(gen[2863]),

			.SELF(gen[2767]),
			.cell_state(gen[2767])
		); 

/******************* CELL 2768 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2768 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2672]),
			.N(gen[2673]),
			.NE(gen[2674]),

			.O(gen[2767]),
			.E(gen[2769]),

			.SO(gen[2862]),
			.S(gen[2863]),
			.SE(gen[2864]),

			.SELF(gen[2768]),
			.cell_state(gen[2768])
		); 

/******************* CELL 2769 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2769 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2673]),
			.N(gen[2674]),
			.NE(gen[2675]),

			.O(gen[2768]),
			.E(gen[2770]),

			.SO(gen[2863]),
			.S(gen[2864]),
			.SE(gen[2865]),

			.SELF(gen[2769]),
			.cell_state(gen[2769])
		); 

/******************* CELL 2770 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2770 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2674]),
			.N(gen[2675]),
			.NE(gen[2676]),

			.O(gen[2769]),
			.E(gen[2771]),

			.SO(gen[2864]),
			.S(gen[2865]),
			.SE(gen[2866]),

			.SELF(gen[2770]),
			.cell_state(gen[2770])
		); 

/******************* CELL 2771 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2771 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2675]),
			.N(gen[2676]),
			.NE(gen[2677]),

			.O(gen[2770]),
			.E(gen[2772]),

			.SO(gen[2865]),
			.S(gen[2866]),
			.SE(gen[2867]),

			.SELF(gen[2771]),
			.cell_state(gen[2771])
		); 

/******************* CELL 2772 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2772 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2676]),
			.N(gen[2677]),
			.NE(gen[2678]),

			.O(gen[2771]),
			.E(gen[2773]),

			.SO(gen[2866]),
			.S(gen[2867]),
			.SE(gen[2868]),

			.SELF(gen[2772]),
			.cell_state(gen[2772])
		); 

/******************* CELL 2773 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2773 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2677]),
			.N(gen[2678]),
			.NE(gen[2679]),

			.O(gen[2772]),
			.E(gen[2774]),

			.SO(gen[2867]),
			.S(gen[2868]),
			.SE(gen[2869]),

			.SELF(gen[2773]),
			.cell_state(gen[2773])
		); 

/******************* CELL 2774 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2774 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2678]),
			.N(gen[2679]),
			.NE(gen[2680]),

			.O(gen[2773]),
			.E(gen[2775]),

			.SO(gen[2868]),
			.S(gen[2869]),
			.SE(gen[2870]),

			.SELF(gen[2774]),
			.cell_state(gen[2774])
		); 

/******************* CELL 2775 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2775 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2679]),
			.N(gen[2680]),
			.NE(gen[2681]),

			.O(gen[2774]),
			.E(gen[2776]),

			.SO(gen[2869]),
			.S(gen[2870]),
			.SE(gen[2871]),

			.SELF(gen[2775]),
			.cell_state(gen[2775])
		); 

/******************* CELL 2776 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2776 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2680]),
			.N(gen[2681]),
			.NE(gen[2682]),

			.O(gen[2775]),
			.E(gen[2777]),

			.SO(gen[2870]),
			.S(gen[2871]),
			.SE(gen[2872]),

			.SELF(gen[2776]),
			.cell_state(gen[2776])
		); 

/******************* CELL 2777 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2777 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2681]),
			.N(gen[2682]),
			.NE(gen[2683]),

			.O(gen[2776]),
			.E(gen[2778]),

			.SO(gen[2871]),
			.S(gen[2872]),
			.SE(gen[2873]),

			.SELF(gen[2777]),
			.cell_state(gen[2777])
		); 

/******************* CELL 2778 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2778 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2682]),
			.N(gen[2683]),
			.NE(gen[2684]),

			.O(gen[2777]),
			.E(gen[2779]),

			.SO(gen[2872]),
			.S(gen[2873]),
			.SE(gen[2874]),

			.SELF(gen[2778]),
			.cell_state(gen[2778])
		); 

/******************* CELL 2779 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2779 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2683]),
			.N(gen[2684]),
			.NE(gen[2685]),

			.O(gen[2778]),
			.E(gen[2780]),

			.SO(gen[2873]),
			.S(gen[2874]),
			.SE(gen[2875]),

			.SELF(gen[2779]),
			.cell_state(gen[2779])
		); 

/******************* CELL 2780 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2780 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2684]),
			.N(gen[2685]),
			.NE(gen[2686]),

			.O(gen[2779]),
			.E(gen[2781]),

			.SO(gen[2874]),
			.S(gen[2875]),
			.SE(gen[2876]),

			.SELF(gen[2780]),
			.cell_state(gen[2780])
		); 

/******************* CELL 2781 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2781 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2685]),
			.N(gen[2686]),
			.NE(gen[2687]),

			.O(gen[2780]),
			.E(gen[2782]),

			.SO(gen[2875]),
			.S(gen[2876]),
			.SE(gen[2877]),

			.SELF(gen[2781]),
			.cell_state(gen[2781])
		); 

/******************* CELL 2782 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2782 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2686]),
			.N(gen[2687]),
			.NE(gen[2688]),

			.O(gen[2781]),
			.E(gen[2783]),

			.SO(gen[2876]),
			.S(gen[2877]),
			.SE(gen[2878]),

			.SELF(gen[2782]),
			.cell_state(gen[2782])
		); 

/******************* CELL 2783 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2783 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2687]),
			.N(gen[2688]),
			.NE(gen[2689]),

			.O(gen[2782]),
			.E(gen[2784]),

			.SO(gen[2877]),
			.S(gen[2878]),
			.SE(gen[2879]),

			.SELF(gen[2783]),
			.cell_state(gen[2783])
		); 

/******************* CELL 2784 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2784 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2688]),
			.N(gen[2689]),
			.NE(gen[2690]),

			.O(gen[2783]),
			.E(gen[2785]),

			.SO(gen[2878]),
			.S(gen[2879]),
			.SE(gen[2880]),

			.SELF(gen[2784]),
			.cell_state(gen[2784])
		); 

/******************* CELL 2785 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2785 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2689]),
			.N(gen[2690]),
			.NE(gen[2691]),

			.O(gen[2784]),
			.E(gen[2786]),

			.SO(gen[2879]),
			.S(gen[2880]),
			.SE(gen[2881]),

			.SELF(gen[2785]),
			.cell_state(gen[2785])
		); 

/******************* CELL 2786 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2786 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2690]),
			.N(gen[2691]),
			.NE(gen[2692]),

			.O(gen[2785]),
			.E(gen[2787]),

			.SO(gen[2880]),
			.S(gen[2881]),
			.SE(gen[2882]),

			.SELF(gen[2786]),
			.cell_state(gen[2786])
		); 

/******************* CELL 2787 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2787 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2691]),
			.N(gen[2692]),
			.NE(gen[2693]),

			.O(gen[2786]),
			.E(gen[2788]),

			.SO(gen[2881]),
			.S(gen[2882]),
			.SE(gen[2883]),

			.SELF(gen[2787]),
			.cell_state(gen[2787])
		); 

/******************* CELL 2788 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2788 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2692]),
			.N(gen[2693]),
			.NE(gen[2694]),

			.O(gen[2787]),
			.E(gen[2789]),

			.SO(gen[2882]),
			.S(gen[2883]),
			.SE(gen[2884]),

			.SELF(gen[2788]),
			.cell_state(gen[2788])
		); 

/******************* CELL 2789 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2789 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2693]),
			.N(gen[2694]),
			.NE(gen[2695]),

			.O(gen[2788]),
			.E(gen[2790]),

			.SO(gen[2883]),
			.S(gen[2884]),
			.SE(gen[2885]),

			.SELF(gen[2789]),
			.cell_state(gen[2789])
		); 

/******************* CELL 2790 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2790 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2694]),
			.N(gen[2695]),
			.NE(gen[2696]),

			.O(gen[2789]),
			.E(gen[2791]),

			.SO(gen[2884]),
			.S(gen[2885]),
			.SE(gen[2886]),

			.SELF(gen[2790]),
			.cell_state(gen[2790])
		); 

/******************* CELL 2791 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2791 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2695]),
			.N(gen[2696]),
			.NE(gen[2697]),

			.O(gen[2790]),
			.E(gen[2792]),

			.SO(gen[2885]),
			.S(gen[2886]),
			.SE(gen[2887]),

			.SELF(gen[2791]),
			.cell_state(gen[2791])
		); 

/******************* CELL 2792 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2792 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2696]),
			.N(gen[2697]),
			.NE(gen[2698]),

			.O(gen[2791]),
			.E(gen[2793]),

			.SO(gen[2886]),
			.S(gen[2887]),
			.SE(gen[2888]),

			.SELF(gen[2792]),
			.cell_state(gen[2792])
		); 

/******************* CELL 2793 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2793 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2697]),
			.N(gen[2698]),
			.NE(gen[2699]),

			.O(gen[2792]),
			.E(gen[2794]),

			.SO(gen[2887]),
			.S(gen[2888]),
			.SE(gen[2889]),

			.SELF(gen[2793]),
			.cell_state(gen[2793])
		); 

/******************* CELL 2794 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2794 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2698]),
			.N(gen[2699]),
			.NE(gen[2700]),

			.O(gen[2793]),
			.E(gen[2795]),

			.SO(gen[2888]),
			.S(gen[2889]),
			.SE(gen[2890]),

			.SELF(gen[2794]),
			.cell_state(gen[2794])
		); 

/******************* CELL 2795 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2795 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2699]),
			.N(gen[2700]),
			.NE(gen[2701]),

			.O(gen[2794]),
			.E(gen[2796]),

			.SO(gen[2889]),
			.S(gen[2890]),
			.SE(gen[2891]),

			.SELF(gen[2795]),
			.cell_state(gen[2795])
		); 

/******************* CELL 2796 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2796 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2700]),
			.N(gen[2701]),
			.NE(gen[2702]),

			.O(gen[2795]),
			.E(gen[2797]),

			.SO(gen[2890]),
			.S(gen[2891]),
			.SE(gen[2892]),

			.SELF(gen[2796]),
			.cell_state(gen[2796])
		); 

/******************* CELL 2797 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2797 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2701]),
			.N(gen[2702]),
			.NE(gen[2703]),

			.O(gen[2796]),
			.E(gen[2798]),

			.SO(gen[2891]),
			.S(gen[2892]),
			.SE(gen[2893]),

			.SELF(gen[2797]),
			.cell_state(gen[2797])
		); 

/******************* CELL 2798 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2798 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2702]),
			.N(gen[2703]),
			.NE(gen[2704]),

			.O(gen[2797]),
			.E(gen[2799]),

			.SO(gen[2892]),
			.S(gen[2893]),
			.SE(gen[2894]),

			.SELF(gen[2798]),
			.cell_state(gen[2798])
		); 

/******************* CELL 2799 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2799 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2703]),
			.N(gen[2704]),
			.NE(gen[2705]),

			.O(gen[2798]),
			.E(gen[2800]),

			.SO(gen[2893]),
			.S(gen[2894]),
			.SE(gen[2895]),

			.SELF(gen[2799]),
			.cell_state(gen[2799])
		); 

/******************* CELL 2800 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2800 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2704]),
			.N(gen[2705]),
			.NE(gen[2706]),

			.O(gen[2799]),
			.E(gen[2801]),

			.SO(gen[2894]),
			.S(gen[2895]),
			.SE(gen[2896]),

			.SELF(gen[2800]),
			.cell_state(gen[2800])
		); 

/******************* CELL 2801 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2801 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2705]),
			.N(gen[2706]),
			.NE(gen[2707]),

			.O(gen[2800]),
			.E(gen[2802]),

			.SO(gen[2895]),
			.S(gen[2896]),
			.SE(gen[2897]),

			.SELF(gen[2801]),
			.cell_state(gen[2801])
		); 

/******************* CELL 2802 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2802 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2706]),
			.N(gen[2707]),
			.NE(gen[2708]),

			.O(gen[2801]),
			.E(gen[2803]),

			.SO(gen[2896]),
			.S(gen[2897]),
			.SE(gen[2898]),

			.SELF(gen[2802]),
			.cell_state(gen[2802])
		); 

/******************* CELL 2803 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2803 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2707]),
			.N(gen[2708]),
			.NE(gen[2709]),

			.O(gen[2802]),
			.E(gen[2804]),

			.SO(gen[2897]),
			.S(gen[2898]),
			.SE(gen[2899]),

			.SELF(gen[2803]),
			.cell_state(gen[2803])
		); 

/******************* CELL 2804 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2804 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2708]),
			.N(gen[2709]),
			.NE(gen[2710]),

			.O(gen[2803]),
			.E(gen[2805]),

			.SO(gen[2898]),
			.S(gen[2899]),
			.SE(gen[2900]),

			.SELF(gen[2804]),
			.cell_state(gen[2804])
		); 

/******************* CELL 2805 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2805 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2709]),
			.N(gen[2710]),
			.NE(gen[2711]),

			.O(gen[2804]),
			.E(gen[2806]),

			.SO(gen[2899]),
			.S(gen[2900]),
			.SE(gen[2901]),

			.SELF(gen[2805]),
			.cell_state(gen[2805])
		); 

/******************* CELL 2806 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2806 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2710]),
			.N(gen[2711]),
			.NE(gen[2712]),

			.O(gen[2805]),
			.E(gen[2807]),

			.SO(gen[2900]),
			.S(gen[2901]),
			.SE(gen[2902]),

			.SELF(gen[2806]),
			.cell_state(gen[2806])
		); 

/******************* CELL 2807 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2807 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2711]),
			.N(gen[2712]),
			.NE(gen[2713]),

			.O(gen[2806]),
			.E(gen[2808]),

			.SO(gen[2901]),
			.S(gen[2902]),
			.SE(gen[2903]),

			.SELF(gen[2807]),
			.cell_state(gen[2807])
		); 

/******************* CELL 2808 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2808 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2712]),
			.N(gen[2713]),
			.NE(gen[2714]),

			.O(gen[2807]),
			.E(gen[2809]),

			.SO(gen[2902]),
			.S(gen[2903]),
			.SE(gen[2904]),

			.SELF(gen[2808]),
			.cell_state(gen[2808])
		); 

/******************* CELL 2809 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2809 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2713]),
			.N(gen[2714]),
			.NE(gen[2715]),

			.O(gen[2808]),
			.E(gen[2810]),

			.SO(gen[2903]),
			.S(gen[2904]),
			.SE(gen[2905]),

			.SELF(gen[2809]),
			.cell_state(gen[2809])
		); 

/******************* CELL 2810 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2810 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2714]),
			.N(gen[2715]),
			.NE(gen[2716]),

			.O(gen[2809]),
			.E(gen[2811]),

			.SO(gen[2904]),
			.S(gen[2905]),
			.SE(gen[2906]),

			.SELF(gen[2810]),
			.cell_state(gen[2810])
		); 

/******************* CELL 2811 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2811 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2715]),
			.N(gen[2716]),
			.NE(gen[2717]),

			.O(gen[2810]),
			.E(gen[2812]),

			.SO(gen[2905]),
			.S(gen[2906]),
			.SE(gen[2907]),

			.SELF(gen[2811]),
			.cell_state(gen[2811])
		); 

/******************* CELL 2812 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2812 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2716]),
			.N(gen[2717]),
			.NE(gen[2718]),

			.O(gen[2811]),
			.E(gen[2813]),

			.SO(gen[2906]),
			.S(gen[2907]),
			.SE(gen[2908]),

			.SELF(gen[2812]),
			.cell_state(gen[2812])
		); 

/******************* CELL 2813 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2813 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2717]),
			.N(gen[2718]),
			.NE(gen[2719]),

			.O(gen[2812]),
			.E(gen[2814]),

			.SO(gen[2907]),
			.S(gen[2908]),
			.SE(gen[2909]),

			.SELF(gen[2813]),
			.cell_state(gen[2813])
		); 

/******************* CELL 2814 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2814 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2718]),
			.N(gen[2719]),
			.NE(gen[2720]),

			.O(gen[2813]),
			.E(gen[2815]),

			.SO(gen[2908]),
			.S(gen[2909]),
			.SE(gen[2910]),

			.SELF(gen[2814]),
			.cell_state(gen[2814])
		); 

/******************* CELL 2815 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2815 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2719]),
			.N(gen[2720]),
			.NE(gen[2721]),

			.O(gen[2814]),
			.E(gen[2816]),

			.SO(gen[2909]),
			.S(gen[2910]),
			.SE(gen[2911]),

			.SELF(gen[2815]),
			.cell_state(gen[2815])
		); 

/******************* CELL 2816 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2816 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2720]),
			.N(gen[2721]),
			.NE(gen[2722]),

			.O(gen[2815]),
			.E(gen[2817]),

			.SO(gen[2910]),
			.S(gen[2911]),
			.SE(gen[2912]),

			.SELF(gen[2816]),
			.cell_state(gen[2816])
		); 

/******************* CELL 2817 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2817 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2721]),
			.N(gen[2722]),
			.NE(gen[2723]),

			.O(gen[2816]),
			.E(gen[2818]),

			.SO(gen[2911]),
			.S(gen[2912]),
			.SE(gen[2913]),

			.SELF(gen[2817]),
			.cell_state(gen[2817])
		); 

/******************* CELL 2818 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2818 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2722]),
			.N(gen[2723]),
			.NE(gen[2724]),

			.O(gen[2817]),
			.E(gen[2819]),

			.SO(gen[2912]),
			.S(gen[2913]),
			.SE(gen[2914]),

			.SELF(gen[2818]),
			.cell_state(gen[2818])
		); 

/******************* CELL 2819 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2819 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2723]),
			.N(gen[2724]),
			.NE(gen[2725]),

			.O(gen[2818]),
			.E(gen[2820]),

			.SO(gen[2913]),
			.S(gen[2914]),
			.SE(gen[2915]),

			.SELF(gen[2819]),
			.cell_state(gen[2819])
		); 

/******************* CELL 2820 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2820 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2724]),
			.N(gen[2725]),
			.NE(gen[2726]),

			.O(gen[2819]),
			.E(gen[2821]),

			.SO(gen[2914]),
			.S(gen[2915]),
			.SE(gen[2916]),

			.SELF(gen[2820]),
			.cell_state(gen[2820])
		); 

/******************* CELL 2821 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2821 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2725]),
			.N(gen[2726]),
			.NE(gen[2727]),

			.O(gen[2820]),
			.E(gen[2822]),

			.SO(gen[2915]),
			.S(gen[2916]),
			.SE(gen[2917]),

			.SELF(gen[2821]),
			.cell_state(gen[2821])
		); 

/******************* CELL 2822 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2822 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2726]),
			.N(gen[2727]),
			.NE(gen[2728]),

			.O(gen[2821]),
			.E(gen[2823]),

			.SO(gen[2916]),
			.S(gen[2917]),
			.SE(gen[2918]),

			.SELF(gen[2822]),
			.cell_state(gen[2822])
		); 

/******************* CELL 2823 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2823 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2727]),
			.N(gen[2728]),
			.NE(gen[2729]),

			.O(gen[2822]),
			.E(gen[2824]),

			.SO(gen[2917]),
			.S(gen[2918]),
			.SE(gen[2919]),

			.SELF(gen[2823]),
			.cell_state(gen[2823])
		); 

/******************* CELL 2824 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2824 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2728]),
			.N(gen[2729]),
			.NE(gen[2730]),

			.O(gen[2823]),
			.E(gen[2825]),

			.SO(gen[2918]),
			.S(gen[2919]),
			.SE(gen[2920]),

			.SELF(gen[2824]),
			.cell_state(gen[2824])
		); 

/******************* CELL 2825 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2825 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2729]),
			.N(gen[2730]),
			.NE(gen[2731]),

			.O(gen[2824]),
			.E(gen[2826]),

			.SO(gen[2919]),
			.S(gen[2920]),
			.SE(gen[2921]),

			.SELF(gen[2825]),
			.cell_state(gen[2825])
		); 

/******************* CELL 2826 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2826 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2730]),
			.N(gen[2731]),
			.NE(gen[2732]),

			.O(gen[2825]),
			.E(gen[2827]),

			.SO(gen[2920]),
			.S(gen[2921]),
			.SE(gen[2922]),

			.SELF(gen[2826]),
			.cell_state(gen[2826])
		); 

/******************* CELL 2827 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2827 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2731]),
			.N(gen[2732]),
			.NE(gen[2733]),

			.O(gen[2826]),
			.E(gen[2828]),

			.SO(gen[2921]),
			.S(gen[2922]),
			.SE(gen[2923]),

			.SELF(gen[2827]),
			.cell_state(gen[2827])
		); 

/******************* CELL 2828 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2828 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2732]),
			.N(gen[2733]),
			.NE(gen[2734]),

			.O(gen[2827]),
			.E(gen[2829]),

			.SO(gen[2922]),
			.S(gen[2923]),
			.SE(gen[2924]),

			.SELF(gen[2828]),
			.cell_state(gen[2828])
		); 

/******************* CELL 2829 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2829 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2733]),
			.N(gen[2734]),
			.NE(gen[2735]),

			.O(gen[2828]),
			.E(gen[2830]),

			.SO(gen[2923]),
			.S(gen[2924]),
			.SE(gen[2925]),

			.SELF(gen[2829]),
			.cell_state(gen[2829])
		); 

/******************* CELL 2830 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2830 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2734]),
			.N(gen[2735]),
			.NE(gen[2736]),

			.O(gen[2829]),
			.E(gen[2831]),

			.SO(gen[2924]),
			.S(gen[2925]),
			.SE(gen[2926]),

			.SELF(gen[2830]),
			.cell_state(gen[2830])
		); 

/******************* CELL 2831 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2831 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2735]),
			.N(gen[2736]),
			.NE(gen[2737]),

			.O(gen[2830]),
			.E(gen[2832]),

			.SO(gen[2925]),
			.S(gen[2926]),
			.SE(gen[2927]),

			.SELF(gen[2831]),
			.cell_state(gen[2831])
		); 

/******************* CELL 2832 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2832 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2736]),
			.N(gen[2737]),
			.NE(gen[2738]),

			.O(gen[2831]),
			.E(gen[2833]),

			.SO(gen[2926]),
			.S(gen[2927]),
			.SE(gen[2928]),

			.SELF(gen[2832]),
			.cell_state(gen[2832])
		); 

/******************* CELL 2833 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2833 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2737]),
			.N(gen[2738]),
			.NE(gen[2739]),

			.O(gen[2832]),
			.E(gen[2834]),

			.SO(gen[2927]),
			.S(gen[2928]),
			.SE(gen[2929]),

			.SELF(gen[2833]),
			.cell_state(gen[2833])
		); 

/******************* CELL 2834 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2834 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2738]),
			.N(gen[2739]),
			.NE(gen[2740]),

			.O(gen[2833]),
			.E(gen[2835]),

			.SO(gen[2928]),
			.S(gen[2929]),
			.SE(gen[2930]),

			.SELF(gen[2834]),
			.cell_state(gen[2834])
		); 

/******************* CELL 2835 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2835 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2739]),
			.N(gen[2740]),
			.NE(gen[2741]),

			.O(gen[2834]),
			.E(gen[2836]),

			.SO(gen[2929]),
			.S(gen[2930]),
			.SE(gen[2931]),

			.SELF(gen[2835]),
			.cell_state(gen[2835])
		); 

/******************* CELL 2836 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2836 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2740]),
			.N(gen[2741]),
			.NE(gen[2742]),

			.O(gen[2835]),
			.E(gen[2837]),

			.SO(gen[2930]),
			.S(gen[2931]),
			.SE(gen[2932]),

			.SELF(gen[2836]),
			.cell_state(gen[2836])
		); 

/******************* CELL 2837 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2837 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2741]),
			.N(gen[2742]),
			.NE(gen[2743]),

			.O(gen[2836]),
			.E(gen[2838]),

			.SO(gen[2931]),
			.S(gen[2932]),
			.SE(gen[2933]),

			.SELF(gen[2837]),
			.cell_state(gen[2837])
		); 

/******************* CELL 2838 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2838 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2742]),
			.N(gen[2743]),
			.NE(gen[2744]),

			.O(gen[2837]),
			.E(gen[2839]),

			.SO(gen[2932]),
			.S(gen[2933]),
			.SE(gen[2934]),

			.SELF(gen[2838]),
			.cell_state(gen[2838])
		); 

/******************* CELL 2839 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2839 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2743]),
			.N(gen[2744]),
			.NE(gen[2745]),

			.O(gen[2838]),
			.E(gen[2840]),

			.SO(gen[2933]),
			.S(gen[2934]),
			.SE(gen[2935]),

			.SELF(gen[2839]),
			.cell_state(gen[2839])
		); 

/******************* CELL 2840 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2840 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2744]),
			.N(gen[2745]),
			.NE(gen[2746]),

			.O(gen[2839]),
			.E(gen[2841]),

			.SO(gen[2934]),
			.S(gen[2935]),
			.SE(gen[2936]),

			.SELF(gen[2840]),
			.cell_state(gen[2840])
		); 

/******************* CELL 2841 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2841 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2745]),
			.N(gen[2746]),
			.NE(gen[2747]),

			.O(gen[2840]),
			.E(gen[2842]),

			.SO(gen[2935]),
			.S(gen[2936]),
			.SE(gen[2937]),

			.SELF(gen[2841]),
			.cell_state(gen[2841])
		); 

/******************* CELL 2842 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2842 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2746]),
			.N(gen[2747]),
			.NE(gen[2748]),

			.O(gen[2841]),
			.E(gen[2843]),

			.SO(gen[2936]),
			.S(gen[2937]),
			.SE(gen[2938]),

			.SELF(gen[2842]),
			.cell_state(gen[2842])
		); 

/******************* CELL 2843 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2843 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2747]),
			.N(gen[2748]),
			.NE(gen[2749]),

			.O(gen[2842]),
			.E(gen[2844]),

			.SO(gen[2937]),
			.S(gen[2938]),
			.SE(gen[2939]),

			.SELF(gen[2843]),
			.cell_state(gen[2843])
		); 

/******************* CELL 2844 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2844 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2748]),
			.N(gen[2749]),
			.NE(gen[2750]),

			.O(gen[2843]),
			.E(gen[2845]),

			.SO(gen[2938]),
			.S(gen[2939]),
			.SE(gen[2940]),

			.SELF(gen[2844]),
			.cell_state(gen[2844])
		); 

/******************* CELL 2845 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2845 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2749]),
			.N(gen[2750]),
			.NE(gen[2751]),

			.O(gen[2844]),
			.E(gen[2846]),

			.SO(gen[2939]),
			.S(gen[2940]),
			.SE(gen[2941]),

			.SELF(gen[2845]),
			.cell_state(gen[2845])
		); 

/******************* CELL 2846 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2846 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2750]),
			.N(gen[2751]),
			.NE(gen[2752]),

			.O(gen[2845]),
			.E(gen[2847]),

			.SO(gen[2940]),
			.S(gen[2941]),
			.SE(gen[2942]),

			.SELF(gen[2846]),
			.cell_state(gen[2846])
		); 

/******************* CELL 2847 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2847 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2751]),
			.N(gen[2752]),
			.NE(gen[2753]),

			.O(gen[2846]),
			.E(gen[2848]),

			.SO(gen[2941]),
			.S(gen[2942]),
			.SE(gen[2943]),

			.SELF(gen[2847]),
			.cell_state(gen[2847])
		); 

/******************* CELL 2848 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2848 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2752]),
			.N(gen[2753]),
			.NE(gen[2754]),

			.O(gen[2847]),
			.E(gen[2849]),

			.SO(gen[2942]),
			.S(gen[2943]),
			.SE(gen[2944]),

			.SELF(gen[2848]),
			.cell_state(gen[2848])
		); 

/******************* CELL 2849 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2849 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2753]),
			.N(gen[2754]),
			.NE(gen[2753]),

			.O(gen[2848]),
			.E(gen[2848]),

			.SO(gen[2943]),
			.S(gen[2944]),
			.SE(gen[2943]),

			.SELF(gen[2849]),
			.cell_state(gen[2849])
		); 

/******************* CELL 2850 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2850 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2756]),
			.N(gen[2755]),
			.NE(gen[2756]),

			.O(gen[2851]),
			.E(gen[2851]),

			.SO(gen[2946]),
			.S(gen[2945]),
			.SE(gen[2946]),

			.SELF(gen[2850]),
			.cell_state(gen[2850])
		); 

/******************* CELL 2851 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2851 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2755]),
			.N(gen[2756]),
			.NE(gen[2757]),

			.O(gen[2850]),
			.E(gen[2852]),

			.SO(gen[2945]),
			.S(gen[2946]),
			.SE(gen[2947]),

			.SELF(gen[2851]),
			.cell_state(gen[2851])
		); 

/******************* CELL 2852 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2852 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2756]),
			.N(gen[2757]),
			.NE(gen[2758]),

			.O(gen[2851]),
			.E(gen[2853]),

			.SO(gen[2946]),
			.S(gen[2947]),
			.SE(gen[2948]),

			.SELF(gen[2852]),
			.cell_state(gen[2852])
		); 

/******************* CELL 2853 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2853 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2757]),
			.N(gen[2758]),
			.NE(gen[2759]),

			.O(gen[2852]),
			.E(gen[2854]),

			.SO(gen[2947]),
			.S(gen[2948]),
			.SE(gen[2949]),

			.SELF(gen[2853]),
			.cell_state(gen[2853])
		); 

/******************* CELL 2854 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2854 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2758]),
			.N(gen[2759]),
			.NE(gen[2760]),

			.O(gen[2853]),
			.E(gen[2855]),

			.SO(gen[2948]),
			.S(gen[2949]),
			.SE(gen[2950]),

			.SELF(gen[2854]),
			.cell_state(gen[2854])
		); 

/******************* CELL 2855 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2855 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2759]),
			.N(gen[2760]),
			.NE(gen[2761]),

			.O(gen[2854]),
			.E(gen[2856]),

			.SO(gen[2949]),
			.S(gen[2950]),
			.SE(gen[2951]),

			.SELF(gen[2855]),
			.cell_state(gen[2855])
		); 

/******************* CELL 2856 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2856 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2760]),
			.N(gen[2761]),
			.NE(gen[2762]),

			.O(gen[2855]),
			.E(gen[2857]),

			.SO(gen[2950]),
			.S(gen[2951]),
			.SE(gen[2952]),

			.SELF(gen[2856]),
			.cell_state(gen[2856])
		); 

/******************* CELL 2857 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2857 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2761]),
			.N(gen[2762]),
			.NE(gen[2763]),

			.O(gen[2856]),
			.E(gen[2858]),

			.SO(gen[2951]),
			.S(gen[2952]),
			.SE(gen[2953]),

			.SELF(gen[2857]),
			.cell_state(gen[2857])
		); 

/******************* CELL 2858 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2858 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2762]),
			.N(gen[2763]),
			.NE(gen[2764]),

			.O(gen[2857]),
			.E(gen[2859]),

			.SO(gen[2952]),
			.S(gen[2953]),
			.SE(gen[2954]),

			.SELF(gen[2858]),
			.cell_state(gen[2858])
		); 

/******************* CELL 2859 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2859 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2763]),
			.N(gen[2764]),
			.NE(gen[2765]),

			.O(gen[2858]),
			.E(gen[2860]),

			.SO(gen[2953]),
			.S(gen[2954]),
			.SE(gen[2955]),

			.SELF(gen[2859]),
			.cell_state(gen[2859])
		); 

/******************* CELL 2860 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2860 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2764]),
			.N(gen[2765]),
			.NE(gen[2766]),

			.O(gen[2859]),
			.E(gen[2861]),

			.SO(gen[2954]),
			.S(gen[2955]),
			.SE(gen[2956]),

			.SELF(gen[2860]),
			.cell_state(gen[2860])
		); 

/******************* CELL 2861 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2861 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2765]),
			.N(gen[2766]),
			.NE(gen[2767]),

			.O(gen[2860]),
			.E(gen[2862]),

			.SO(gen[2955]),
			.S(gen[2956]),
			.SE(gen[2957]),

			.SELF(gen[2861]),
			.cell_state(gen[2861])
		); 

/******************* CELL 2862 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2862 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2766]),
			.N(gen[2767]),
			.NE(gen[2768]),

			.O(gen[2861]),
			.E(gen[2863]),

			.SO(gen[2956]),
			.S(gen[2957]),
			.SE(gen[2958]),

			.SELF(gen[2862]),
			.cell_state(gen[2862])
		); 

/******************* CELL 2863 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2863 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2767]),
			.N(gen[2768]),
			.NE(gen[2769]),

			.O(gen[2862]),
			.E(gen[2864]),

			.SO(gen[2957]),
			.S(gen[2958]),
			.SE(gen[2959]),

			.SELF(gen[2863]),
			.cell_state(gen[2863])
		); 

/******************* CELL 2864 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2864 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2768]),
			.N(gen[2769]),
			.NE(gen[2770]),

			.O(gen[2863]),
			.E(gen[2865]),

			.SO(gen[2958]),
			.S(gen[2959]),
			.SE(gen[2960]),

			.SELF(gen[2864]),
			.cell_state(gen[2864])
		); 

/******************* CELL 2865 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2865 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2769]),
			.N(gen[2770]),
			.NE(gen[2771]),

			.O(gen[2864]),
			.E(gen[2866]),

			.SO(gen[2959]),
			.S(gen[2960]),
			.SE(gen[2961]),

			.SELF(gen[2865]),
			.cell_state(gen[2865])
		); 

/******************* CELL 2866 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2866 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2770]),
			.N(gen[2771]),
			.NE(gen[2772]),

			.O(gen[2865]),
			.E(gen[2867]),

			.SO(gen[2960]),
			.S(gen[2961]),
			.SE(gen[2962]),

			.SELF(gen[2866]),
			.cell_state(gen[2866])
		); 

/******************* CELL 2867 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2867 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2771]),
			.N(gen[2772]),
			.NE(gen[2773]),

			.O(gen[2866]),
			.E(gen[2868]),

			.SO(gen[2961]),
			.S(gen[2962]),
			.SE(gen[2963]),

			.SELF(gen[2867]),
			.cell_state(gen[2867])
		); 

/******************* CELL 2868 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2868 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2772]),
			.N(gen[2773]),
			.NE(gen[2774]),

			.O(gen[2867]),
			.E(gen[2869]),

			.SO(gen[2962]),
			.S(gen[2963]),
			.SE(gen[2964]),

			.SELF(gen[2868]),
			.cell_state(gen[2868])
		); 

/******************* CELL 2869 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2869 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2773]),
			.N(gen[2774]),
			.NE(gen[2775]),

			.O(gen[2868]),
			.E(gen[2870]),

			.SO(gen[2963]),
			.S(gen[2964]),
			.SE(gen[2965]),

			.SELF(gen[2869]),
			.cell_state(gen[2869])
		); 

/******************* CELL 2870 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2870 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2774]),
			.N(gen[2775]),
			.NE(gen[2776]),

			.O(gen[2869]),
			.E(gen[2871]),

			.SO(gen[2964]),
			.S(gen[2965]),
			.SE(gen[2966]),

			.SELF(gen[2870]),
			.cell_state(gen[2870])
		); 

/******************* CELL 2871 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2871 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2775]),
			.N(gen[2776]),
			.NE(gen[2777]),

			.O(gen[2870]),
			.E(gen[2872]),

			.SO(gen[2965]),
			.S(gen[2966]),
			.SE(gen[2967]),

			.SELF(gen[2871]),
			.cell_state(gen[2871])
		); 

/******************* CELL 2872 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2872 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2776]),
			.N(gen[2777]),
			.NE(gen[2778]),

			.O(gen[2871]),
			.E(gen[2873]),

			.SO(gen[2966]),
			.S(gen[2967]),
			.SE(gen[2968]),

			.SELF(gen[2872]),
			.cell_state(gen[2872])
		); 

/******************* CELL 2873 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2873 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2777]),
			.N(gen[2778]),
			.NE(gen[2779]),

			.O(gen[2872]),
			.E(gen[2874]),

			.SO(gen[2967]),
			.S(gen[2968]),
			.SE(gen[2969]),

			.SELF(gen[2873]),
			.cell_state(gen[2873])
		); 

/******************* CELL 2874 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2874 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2778]),
			.N(gen[2779]),
			.NE(gen[2780]),

			.O(gen[2873]),
			.E(gen[2875]),

			.SO(gen[2968]),
			.S(gen[2969]),
			.SE(gen[2970]),

			.SELF(gen[2874]),
			.cell_state(gen[2874])
		); 

/******************* CELL 2875 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2875 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2779]),
			.N(gen[2780]),
			.NE(gen[2781]),

			.O(gen[2874]),
			.E(gen[2876]),

			.SO(gen[2969]),
			.S(gen[2970]),
			.SE(gen[2971]),

			.SELF(gen[2875]),
			.cell_state(gen[2875])
		); 

/******************* CELL 2876 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2876 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2780]),
			.N(gen[2781]),
			.NE(gen[2782]),

			.O(gen[2875]),
			.E(gen[2877]),

			.SO(gen[2970]),
			.S(gen[2971]),
			.SE(gen[2972]),

			.SELF(gen[2876]),
			.cell_state(gen[2876])
		); 

/******************* CELL 2877 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2877 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2781]),
			.N(gen[2782]),
			.NE(gen[2783]),

			.O(gen[2876]),
			.E(gen[2878]),

			.SO(gen[2971]),
			.S(gen[2972]),
			.SE(gen[2973]),

			.SELF(gen[2877]),
			.cell_state(gen[2877])
		); 

/******************* CELL 2878 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2878 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2782]),
			.N(gen[2783]),
			.NE(gen[2784]),

			.O(gen[2877]),
			.E(gen[2879]),

			.SO(gen[2972]),
			.S(gen[2973]),
			.SE(gen[2974]),

			.SELF(gen[2878]),
			.cell_state(gen[2878])
		); 

/******************* CELL 2879 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2879 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2783]),
			.N(gen[2784]),
			.NE(gen[2785]),

			.O(gen[2878]),
			.E(gen[2880]),

			.SO(gen[2973]),
			.S(gen[2974]),
			.SE(gen[2975]),

			.SELF(gen[2879]),
			.cell_state(gen[2879])
		); 

/******************* CELL 2880 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2880 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2784]),
			.N(gen[2785]),
			.NE(gen[2786]),

			.O(gen[2879]),
			.E(gen[2881]),

			.SO(gen[2974]),
			.S(gen[2975]),
			.SE(gen[2976]),

			.SELF(gen[2880]),
			.cell_state(gen[2880])
		); 

/******************* CELL 2881 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2881 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2785]),
			.N(gen[2786]),
			.NE(gen[2787]),

			.O(gen[2880]),
			.E(gen[2882]),

			.SO(gen[2975]),
			.S(gen[2976]),
			.SE(gen[2977]),

			.SELF(gen[2881]),
			.cell_state(gen[2881])
		); 

/******************* CELL 2882 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2882 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2786]),
			.N(gen[2787]),
			.NE(gen[2788]),

			.O(gen[2881]),
			.E(gen[2883]),

			.SO(gen[2976]),
			.S(gen[2977]),
			.SE(gen[2978]),

			.SELF(gen[2882]),
			.cell_state(gen[2882])
		); 

/******************* CELL 2883 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2883 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2787]),
			.N(gen[2788]),
			.NE(gen[2789]),

			.O(gen[2882]),
			.E(gen[2884]),

			.SO(gen[2977]),
			.S(gen[2978]),
			.SE(gen[2979]),

			.SELF(gen[2883]),
			.cell_state(gen[2883])
		); 

/******************* CELL 2884 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2884 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2788]),
			.N(gen[2789]),
			.NE(gen[2790]),

			.O(gen[2883]),
			.E(gen[2885]),

			.SO(gen[2978]),
			.S(gen[2979]),
			.SE(gen[2980]),

			.SELF(gen[2884]),
			.cell_state(gen[2884])
		); 

/******************* CELL 2885 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2885 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2789]),
			.N(gen[2790]),
			.NE(gen[2791]),

			.O(gen[2884]),
			.E(gen[2886]),

			.SO(gen[2979]),
			.S(gen[2980]),
			.SE(gen[2981]),

			.SELF(gen[2885]),
			.cell_state(gen[2885])
		); 

/******************* CELL 2886 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2886 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2790]),
			.N(gen[2791]),
			.NE(gen[2792]),

			.O(gen[2885]),
			.E(gen[2887]),

			.SO(gen[2980]),
			.S(gen[2981]),
			.SE(gen[2982]),

			.SELF(gen[2886]),
			.cell_state(gen[2886])
		); 

/******************* CELL 2887 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2887 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2791]),
			.N(gen[2792]),
			.NE(gen[2793]),

			.O(gen[2886]),
			.E(gen[2888]),

			.SO(gen[2981]),
			.S(gen[2982]),
			.SE(gen[2983]),

			.SELF(gen[2887]),
			.cell_state(gen[2887])
		); 

/******************* CELL 2888 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2888 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2792]),
			.N(gen[2793]),
			.NE(gen[2794]),

			.O(gen[2887]),
			.E(gen[2889]),

			.SO(gen[2982]),
			.S(gen[2983]),
			.SE(gen[2984]),

			.SELF(gen[2888]),
			.cell_state(gen[2888])
		); 

/******************* CELL 2889 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2889 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2793]),
			.N(gen[2794]),
			.NE(gen[2795]),

			.O(gen[2888]),
			.E(gen[2890]),

			.SO(gen[2983]),
			.S(gen[2984]),
			.SE(gen[2985]),

			.SELF(gen[2889]),
			.cell_state(gen[2889])
		); 

/******************* CELL 2890 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2890 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2794]),
			.N(gen[2795]),
			.NE(gen[2796]),

			.O(gen[2889]),
			.E(gen[2891]),

			.SO(gen[2984]),
			.S(gen[2985]),
			.SE(gen[2986]),

			.SELF(gen[2890]),
			.cell_state(gen[2890])
		); 

/******************* CELL 2891 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2891 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2795]),
			.N(gen[2796]),
			.NE(gen[2797]),

			.O(gen[2890]),
			.E(gen[2892]),

			.SO(gen[2985]),
			.S(gen[2986]),
			.SE(gen[2987]),

			.SELF(gen[2891]),
			.cell_state(gen[2891])
		); 

/******************* CELL 2892 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2892 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2796]),
			.N(gen[2797]),
			.NE(gen[2798]),

			.O(gen[2891]),
			.E(gen[2893]),

			.SO(gen[2986]),
			.S(gen[2987]),
			.SE(gen[2988]),

			.SELF(gen[2892]),
			.cell_state(gen[2892])
		); 

/******************* CELL 2893 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2893 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2797]),
			.N(gen[2798]),
			.NE(gen[2799]),

			.O(gen[2892]),
			.E(gen[2894]),

			.SO(gen[2987]),
			.S(gen[2988]),
			.SE(gen[2989]),

			.SELF(gen[2893]),
			.cell_state(gen[2893])
		); 

/******************* CELL 2894 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2894 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2798]),
			.N(gen[2799]),
			.NE(gen[2800]),

			.O(gen[2893]),
			.E(gen[2895]),

			.SO(gen[2988]),
			.S(gen[2989]),
			.SE(gen[2990]),

			.SELF(gen[2894]),
			.cell_state(gen[2894])
		); 

/******************* CELL 2895 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2895 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2799]),
			.N(gen[2800]),
			.NE(gen[2801]),

			.O(gen[2894]),
			.E(gen[2896]),

			.SO(gen[2989]),
			.S(gen[2990]),
			.SE(gen[2991]),

			.SELF(gen[2895]),
			.cell_state(gen[2895])
		); 

/******************* CELL 2896 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2896 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2800]),
			.N(gen[2801]),
			.NE(gen[2802]),

			.O(gen[2895]),
			.E(gen[2897]),

			.SO(gen[2990]),
			.S(gen[2991]),
			.SE(gen[2992]),

			.SELF(gen[2896]),
			.cell_state(gen[2896])
		); 

/******************* CELL 2897 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2897 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2801]),
			.N(gen[2802]),
			.NE(gen[2803]),

			.O(gen[2896]),
			.E(gen[2898]),

			.SO(gen[2991]),
			.S(gen[2992]),
			.SE(gen[2993]),

			.SELF(gen[2897]),
			.cell_state(gen[2897])
		); 

/******************* CELL 2898 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2898 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2802]),
			.N(gen[2803]),
			.NE(gen[2804]),

			.O(gen[2897]),
			.E(gen[2899]),

			.SO(gen[2992]),
			.S(gen[2993]),
			.SE(gen[2994]),

			.SELF(gen[2898]),
			.cell_state(gen[2898])
		); 

/******************* CELL 2899 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2899 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2803]),
			.N(gen[2804]),
			.NE(gen[2805]),

			.O(gen[2898]),
			.E(gen[2900]),

			.SO(gen[2993]),
			.S(gen[2994]),
			.SE(gen[2995]),

			.SELF(gen[2899]),
			.cell_state(gen[2899])
		); 

/******************* CELL 2900 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2900 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2804]),
			.N(gen[2805]),
			.NE(gen[2806]),

			.O(gen[2899]),
			.E(gen[2901]),

			.SO(gen[2994]),
			.S(gen[2995]),
			.SE(gen[2996]),

			.SELF(gen[2900]),
			.cell_state(gen[2900])
		); 

/******************* CELL 2901 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2901 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2805]),
			.N(gen[2806]),
			.NE(gen[2807]),

			.O(gen[2900]),
			.E(gen[2902]),

			.SO(gen[2995]),
			.S(gen[2996]),
			.SE(gen[2997]),

			.SELF(gen[2901]),
			.cell_state(gen[2901])
		); 

/******************* CELL 2902 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2902 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2806]),
			.N(gen[2807]),
			.NE(gen[2808]),

			.O(gen[2901]),
			.E(gen[2903]),

			.SO(gen[2996]),
			.S(gen[2997]),
			.SE(gen[2998]),

			.SELF(gen[2902]),
			.cell_state(gen[2902])
		); 

/******************* CELL 2903 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2903 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2807]),
			.N(gen[2808]),
			.NE(gen[2809]),

			.O(gen[2902]),
			.E(gen[2904]),

			.SO(gen[2997]),
			.S(gen[2998]),
			.SE(gen[2999]),

			.SELF(gen[2903]),
			.cell_state(gen[2903])
		); 

/******************* CELL 2904 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2904 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2808]),
			.N(gen[2809]),
			.NE(gen[2810]),

			.O(gen[2903]),
			.E(gen[2905]),

			.SO(gen[2998]),
			.S(gen[2999]),
			.SE(gen[3000]),

			.SELF(gen[2904]),
			.cell_state(gen[2904])
		); 

/******************* CELL 2905 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2905 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2809]),
			.N(gen[2810]),
			.NE(gen[2811]),

			.O(gen[2904]),
			.E(gen[2906]),

			.SO(gen[2999]),
			.S(gen[3000]),
			.SE(gen[3001]),

			.SELF(gen[2905]),
			.cell_state(gen[2905])
		); 

/******************* CELL 2906 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2906 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2810]),
			.N(gen[2811]),
			.NE(gen[2812]),

			.O(gen[2905]),
			.E(gen[2907]),

			.SO(gen[3000]),
			.S(gen[3001]),
			.SE(gen[3002]),

			.SELF(gen[2906]),
			.cell_state(gen[2906])
		); 

/******************* CELL 2907 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2907 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2811]),
			.N(gen[2812]),
			.NE(gen[2813]),

			.O(gen[2906]),
			.E(gen[2908]),

			.SO(gen[3001]),
			.S(gen[3002]),
			.SE(gen[3003]),

			.SELF(gen[2907]),
			.cell_state(gen[2907])
		); 

/******************* CELL 2908 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2908 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2812]),
			.N(gen[2813]),
			.NE(gen[2814]),

			.O(gen[2907]),
			.E(gen[2909]),

			.SO(gen[3002]),
			.S(gen[3003]),
			.SE(gen[3004]),

			.SELF(gen[2908]),
			.cell_state(gen[2908])
		); 

/******************* CELL 2909 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2909 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2813]),
			.N(gen[2814]),
			.NE(gen[2815]),

			.O(gen[2908]),
			.E(gen[2910]),

			.SO(gen[3003]),
			.S(gen[3004]),
			.SE(gen[3005]),

			.SELF(gen[2909]),
			.cell_state(gen[2909])
		); 

/******************* CELL 2910 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2910 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2814]),
			.N(gen[2815]),
			.NE(gen[2816]),

			.O(gen[2909]),
			.E(gen[2911]),

			.SO(gen[3004]),
			.S(gen[3005]),
			.SE(gen[3006]),

			.SELF(gen[2910]),
			.cell_state(gen[2910])
		); 

/******************* CELL 2911 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2911 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2815]),
			.N(gen[2816]),
			.NE(gen[2817]),

			.O(gen[2910]),
			.E(gen[2912]),

			.SO(gen[3005]),
			.S(gen[3006]),
			.SE(gen[3007]),

			.SELF(gen[2911]),
			.cell_state(gen[2911])
		); 

/******************* CELL 2912 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2912 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2816]),
			.N(gen[2817]),
			.NE(gen[2818]),

			.O(gen[2911]),
			.E(gen[2913]),

			.SO(gen[3006]),
			.S(gen[3007]),
			.SE(gen[3008]),

			.SELF(gen[2912]),
			.cell_state(gen[2912])
		); 

/******************* CELL 2913 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2913 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2817]),
			.N(gen[2818]),
			.NE(gen[2819]),

			.O(gen[2912]),
			.E(gen[2914]),

			.SO(gen[3007]),
			.S(gen[3008]),
			.SE(gen[3009]),

			.SELF(gen[2913]),
			.cell_state(gen[2913])
		); 

/******************* CELL 2914 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2914 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2818]),
			.N(gen[2819]),
			.NE(gen[2820]),

			.O(gen[2913]),
			.E(gen[2915]),

			.SO(gen[3008]),
			.S(gen[3009]),
			.SE(gen[3010]),

			.SELF(gen[2914]),
			.cell_state(gen[2914])
		); 

/******************* CELL 2915 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2915 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2819]),
			.N(gen[2820]),
			.NE(gen[2821]),

			.O(gen[2914]),
			.E(gen[2916]),

			.SO(gen[3009]),
			.S(gen[3010]),
			.SE(gen[3011]),

			.SELF(gen[2915]),
			.cell_state(gen[2915])
		); 

/******************* CELL 2916 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2916 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2820]),
			.N(gen[2821]),
			.NE(gen[2822]),

			.O(gen[2915]),
			.E(gen[2917]),

			.SO(gen[3010]),
			.S(gen[3011]),
			.SE(gen[3012]),

			.SELF(gen[2916]),
			.cell_state(gen[2916])
		); 

/******************* CELL 2917 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2917 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2821]),
			.N(gen[2822]),
			.NE(gen[2823]),

			.O(gen[2916]),
			.E(gen[2918]),

			.SO(gen[3011]),
			.S(gen[3012]),
			.SE(gen[3013]),

			.SELF(gen[2917]),
			.cell_state(gen[2917])
		); 

/******************* CELL 2918 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2918 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2822]),
			.N(gen[2823]),
			.NE(gen[2824]),

			.O(gen[2917]),
			.E(gen[2919]),

			.SO(gen[3012]),
			.S(gen[3013]),
			.SE(gen[3014]),

			.SELF(gen[2918]),
			.cell_state(gen[2918])
		); 

/******************* CELL 2919 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2919 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2823]),
			.N(gen[2824]),
			.NE(gen[2825]),

			.O(gen[2918]),
			.E(gen[2920]),

			.SO(gen[3013]),
			.S(gen[3014]),
			.SE(gen[3015]),

			.SELF(gen[2919]),
			.cell_state(gen[2919])
		); 

/******************* CELL 2920 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2920 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2824]),
			.N(gen[2825]),
			.NE(gen[2826]),

			.O(gen[2919]),
			.E(gen[2921]),

			.SO(gen[3014]),
			.S(gen[3015]),
			.SE(gen[3016]),

			.SELF(gen[2920]),
			.cell_state(gen[2920])
		); 

/******************* CELL 2921 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2921 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2825]),
			.N(gen[2826]),
			.NE(gen[2827]),

			.O(gen[2920]),
			.E(gen[2922]),

			.SO(gen[3015]),
			.S(gen[3016]),
			.SE(gen[3017]),

			.SELF(gen[2921]),
			.cell_state(gen[2921])
		); 

/******************* CELL 2922 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2922 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2826]),
			.N(gen[2827]),
			.NE(gen[2828]),

			.O(gen[2921]),
			.E(gen[2923]),

			.SO(gen[3016]),
			.S(gen[3017]),
			.SE(gen[3018]),

			.SELF(gen[2922]),
			.cell_state(gen[2922])
		); 

/******************* CELL 2923 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2923 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2827]),
			.N(gen[2828]),
			.NE(gen[2829]),

			.O(gen[2922]),
			.E(gen[2924]),

			.SO(gen[3017]),
			.S(gen[3018]),
			.SE(gen[3019]),

			.SELF(gen[2923]),
			.cell_state(gen[2923])
		); 

/******************* CELL 2924 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2924 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2828]),
			.N(gen[2829]),
			.NE(gen[2830]),

			.O(gen[2923]),
			.E(gen[2925]),

			.SO(gen[3018]),
			.S(gen[3019]),
			.SE(gen[3020]),

			.SELF(gen[2924]),
			.cell_state(gen[2924])
		); 

/******************* CELL 2925 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2925 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2829]),
			.N(gen[2830]),
			.NE(gen[2831]),

			.O(gen[2924]),
			.E(gen[2926]),

			.SO(gen[3019]),
			.S(gen[3020]),
			.SE(gen[3021]),

			.SELF(gen[2925]),
			.cell_state(gen[2925])
		); 

/******************* CELL 2926 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2926 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2830]),
			.N(gen[2831]),
			.NE(gen[2832]),

			.O(gen[2925]),
			.E(gen[2927]),

			.SO(gen[3020]),
			.S(gen[3021]),
			.SE(gen[3022]),

			.SELF(gen[2926]),
			.cell_state(gen[2926])
		); 

/******************* CELL 2927 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2927 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2831]),
			.N(gen[2832]),
			.NE(gen[2833]),

			.O(gen[2926]),
			.E(gen[2928]),

			.SO(gen[3021]),
			.S(gen[3022]),
			.SE(gen[3023]),

			.SELF(gen[2927]),
			.cell_state(gen[2927])
		); 

/******************* CELL 2928 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2928 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2832]),
			.N(gen[2833]),
			.NE(gen[2834]),

			.O(gen[2927]),
			.E(gen[2929]),

			.SO(gen[3022]),
			.S(gen[3023]),
			.SE(gen[3024]),

			.SELF(gen[2928]),
			.cell_state(gen[2928])
		); 

/******************* CELL 2929 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2929 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2833]),
			.N(gen[2834]),
			.NE(gen[2835]),

			.O(gen[2928]),
			.E(gen[2930]),

			.SO(gen[3023]),
			.S(gen[3024]),
			.SE(gen[3025]),

			.SELF(gen[2929]),
			.cell_state(gen[2929])
		); 

/******************* CELL 2930 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2930 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2834]),
			.N(gen[2835]),
			.NE(gen[2836]),

			.O(gen[2929]),
			.E(gen[2931]),

			.SO(gen[3024]),
			.S(gen[3025]),
			.SE(gen[3026]),

			.SELF(gen[2930]),
			.cell_state(gen[2930])
		); 

/******************* CELL 2931 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2931 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2835]),
			.N(gen[2836]),
			.NE(gen[2837]),

			.O(gen[2930]),
			.E(gen[2932]),

			.SO(gen[3025]),
			.S(gen[3026]),
			.SE(gen[3027]),

			.SELF(gen[2931]),
			.cell_state(gen[2931])
		); 

/******************* CELL 2932 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2932 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2836]),
			.N(gen[2837]),
			.NE(gen[2838]),

			.O(gen[2931]),
			.E(gen[2933]),

			.SO(gen[3026]),
			.S(gen[3027]),
			.SE(gen[3028]),

			.SELF(gen[2932]),
			.cell_state(gen[2932])
		); 

/******************* CELL 2933 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2933 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2837]),
			.N(gen[2838]),
			.NE(gen[2839]),

			.O(gen[2932]),
			.E(gen[2934]),

			.SO(gen[3027]),
			.S(gen[3028]),
			.SE(gen[3029]),

			.SELF(gen[2933]),
			.cell_state(gen[2933])
		); 

/******************* CELL 2934 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2934 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2838]),
			.N(gen[2839]),
			.NE(gen[2840]),

			.O(gen[2933]),
			.E(gen[2935]),

			.SO(gen[3028]),
			.S(gen[3029]),
			.SE(gen[3030]),

			.SELF(gen[2934]),
			.cell_state(gen[2934])
		); 

/******************* CELL 2935 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2935 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2839]),
			.N(gen[2840]),
			.NE(gen[2841]),

			.O(gen[2934]),
			.E(gen[2936]),

			.SO(gen[3029]),
			.S(gen[3030]),
			.SE(gen[3031]),

			.SELF(gen[2935]),
			.cell_state(gen[2935])
		); 

/******************* CELL 2936 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2936 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2840]),
			.N(gen[2841]),
			.NE(gen[2842]),

			.O(gen[2935]),
			.E(gen[2937]),

			.SO(gen[3030]),
			.S(gen[3031]),
			.SE(gen[3032]),

			.SELF(gen[2936]),
			.cell_state(gen[2936])
		); 

/******************* CELL 2937 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2937 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2841]),
			.N(gen[2842]),
			.NE(gen[2843]),

			.O(gen[2936]),
			.E(gen[2938]),

			.SO(gen[3031]),
			.S(gen[3032]),
			.SE(gen[3033]),

			.SELF(gen[2937]),
			.cell_state(gen[2937])
		); 

/******************* CELL 2938 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2938 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2842]),
			.N(gen[2843]),
			.NE(gen[2844]),

			.O(gen[2937]),
			.E(gen[2939]),

			.SO(gen[3032]),
			.S(gen[3033]),
			.SE(gen[3034]),

			.SELF(gen[2938]),
			.cell_state(gen[2938])
		); 

/******************* CELL 2939 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2939 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2843]),
			.N(gen[2844]),
			.NE(gen[2845]),

			.O(gen[2938]),
			.E(gen[2940]),

			.SO(gen[3033]),
			.S(gen[3034]),
			.SE(gen[3035]),

			.SELF(gen[2939]),
			.cell_state(gen[2939])
		); 

/******************* CELL 2940 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2940 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2844]),
			.N(gen[2845]),
			.NE(gen[2846]),

			.O(gen[2939]),
			.E(gen[2941]),

			.SO(gen[3034]),
			.S(gen[3035]),
			.SE(gen[3036]),

			.SELF(gen[2940]),
			.cell_state(gen[2940])
		); 

/******************* CELL 2941 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2941 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2845]),
			.N(gen[2846]),
			.NE(gen[2847]),

			.O(gen[2940]),
			.E(gen[2942]),

			.SO(gen[3035]),
			.S(gen[3036]),
			.SE(gen[3037]),

			.SELF(gen[2941]),
			.cell_state(gen[2941])
		); 

/******************* CELL 2942 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2942 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2846]),
			.N(gen[2847]),
			.NE(gen[2848]),

			.O(gen[2941]),
			.E(gen[2943]),

			.SO(gen[3036]),
			.S(gen[3037]),
			.SE(gen[3038]),

			.SELF(gen[2942]),
			.cell_state(gen[2942])
		); 

/******************* CELL 2943 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2943 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2847]),
			.N(gen[2848]),
			.NE(gen[2849]),

			.O(gen[2942]),
			.E(gen[2944]),

			.SO(gen[3037]),
			.S(gen[3038]),
			.SE(gen[3039]),

			.SELF(gen[2943]),
			.cell_state(gen[2943])
		); 

/******************* CELL 2944 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2944 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2848]),
			.N(gen[2849]),
			.NE(gen[2848]),

			.O(gen[2943]),
			.E(gen[2943]),

			.SO(gen[3038]),
			.S(gen[3039]),
			.SE(gen[3038]),

			.SELF(gen[2944]),
			.cell_state(gen[2944])
		); 

/******************* CELL 2945 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2945 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2851]),
			.N(gen[2850]),
			.NE(gen[2851]),

			.O(gen[2946]),
			.E(gen[2946]),

			.SO(gen[3041]),
			.S(gen[3040]),
			.SE(gen[3041]),

			.SELF(gen[2945]),
			.cell_state(gen[2945])
		); 

/******************* CELL 2946 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2946 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2850]),
			.N(gen[2851]),
			.NE(gen[2852]),

			.O(gen[2945]),
			.E(gen[2947]),

			.SO(gen[3040]),
			.S(gen[3041]),
			.SE(gen[3042]),

			.SELF(gen[2946]),
			.cell_state(gen[2946])
		); 

/******************* CELL 2947 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2947 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2851]),
			.N(gen[2852]),
			.NE(gen[2853]),

			.O(gen[2946]),
			.E(gen[2948]),

			.SO(gen[3041]),
			.S(gen[3042]),
			.SE(gen[3043]),

			.SELF(gen[2947]),
			.cell_state(gen[2947])
		); 

/******************* CELL 2948 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2948 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2852]),
			.N(gen[2853]),
			.NE(gen[2854]),

			.O(gen[2947]),
			.E(gen[2949]),

			.SO(gen[3042]),
			.S(gen[3043]),
			.SE(gen[3044]),

			.SELF(gen[2948]),
			.cell_state(gen[2948])
		); 

/******************* CELL 2949 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2949 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2853]),
			.N(gen[2854]),
			.NE(gen[2855]),

			.O(gen[2948]),
			.E(gen[2950]),

			.SO(gen[3043]),
			.S(gen[3044]),
			.SE(gen[3045]),

			.SELF(gen[2949]),
			.cell_state(gen[2949])
		); 

/******************* CELL 2950 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2950 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2854]),
			.N(gen[2855]),
			.NE(gen[2856]),

			.O(gen[2949]),
			.E(gen[2951]),

			.SO(gen[3044]),
			.S(gen[3045]),
			.SE(gen[3046]),

			.SELF(gen[2950]),
			.cell_state(gen[2950])
		); 

/******************* CELL 2951 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2951 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2855]),
			.N(gen[2856]),
			.NE(gen[2857]),

			.O(gen[2950]),
			.E(gen[2952]),

			.SO(gen[3045]),
			.S(gen[3046]),
			.SE(gen[3047]),

			.SELF(gen[2951]),
			.cell_state(gen[2951])
		); 

/******************* CELL 2952 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2952 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2856]),
			.N(gen[2857]),
			.NE(gen[2858]),

			.O(gen[2951]),
			.E(gen[2953]),

			.SO(gen[3046]),
			.S(gen[3047]),
			.SE(gen[3048]),

			.SELF(gen[2952]),
			.cell_state(gen[2952])
		); 

/******************* CELL 2953 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2953 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2857]),
			.N(gen[2858]),
			.NE(gen[2859]),

			.O(gen[2952]),
			.E(gen[2954]),

			.SO(gen[3047]),
			.S(gen[3048]),
			.SE(gen[3049]),

			.SELF(gen[2953]),
			.cell_state(gen[2953])
		); 

/******************* CELL 2954 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2954 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2858]),
			.N(gen[2859]),
			.NE(gen[2860]),

			.O(gen[2953]),
			.E(gen[2955]),

			.SO(gen[3048]),
			.S(gen[3049]),
			.SE(gen[3050]),

			.SELF(gen[2954]),
			.cell_state(gen[2954])
		); 

/******************* CELL 2955 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2955 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2859]),
			.N(gen[2860]),
			.NE(gen[2861]),

			.O(gen[2954]),
			.E(gen[2956]),

			.SO(gen[3049]),
			.S(gen[3050]),
			.SE(gen[3051]),

			.SELF(gen[2955]),
			.cell_state(gen[2955])
		); 

/******************* CELL 2956 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2956 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2860]),
			.N(gen[2861]),
			.NE(gen[2862]),

			.O(gen[2955]),
			.E(gen[2957]),

			.SO(gen[3050]),
			.S(gen[3051]),
			.SE(gen[3052]),

			.SELF(gen[2956]),
			.cell_state(gen[2956])
		); 

/******************* CELL 2957 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2957 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2861]),
			.N(gen[2862]),
			.NE(gen[2863]),

			.O(gen[2956]),
			.E(gen[2958]),

			.SO(gen[3051]),
			.S(gen[3052]),
			.SE(gen[3053]),

			.SELF(gen[2957]),
			.cell_state(gen[2957])
		); 

/******************* CELL 2958 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2958 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2862]),
			.N(gen[2863]),
			.NE(gen[2864]),

			.O(gen[2957]),
			.E(gen[2959]),

			.SO(gen[3052]),
			.S(gen[3053]),
			.SE(gen[3054]),

			.SELF(gen[2958]),
			.cell_state(gen[2958])
		); 

/******************* CELL 2959 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2959 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2863]),
			.N(gen[2864]),
			.NE(gen[2865]),

			.O(gen[2958]),
			.E(gen[2960]),

			.SO(gen[3053]),
			.S(gen[3054]),
			.SE(gen[3055]),

			.SELF(gen[2959]),
			.cell_state(gen[2959])
		); 

/******************* CELL 2960 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2960 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2864]),
			.N(gen[2865]),
			.NE(gen[2866]),

			.O(gen[2959]),
			.E(gen[2961]),

			.SO(gen[3054]),
			.S(gen[3055]),
			.SE(gen[3056]),

			.SELF(gen[2960]),
			.cell_state(gen[2960])
		); 

/******************* CELL 2961 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2961 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2865]),
			.N(gen[2866]),
			.NE(gen[2867]),

			.O(gen[2960]),
			.E(gen[2962]),

			.SO(gen[3055]),
			.S(gen[3056]),
			.SE(gen[3057]),

			.SELF(gen[2961]),
			.cell_state(gen[2961])
		); 

/******************* CELL 2962 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2962 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2866]),
			.N(gen[2867]),
			.NE(gen[2868]),

			.O(gen[2961]),
			.E(gen[2963]),

			.SO(gen[3056]),
			.S(gen[3057]),
			.SE(gen[3058]),

			.SELF(gen[2962]),
			.cell_state(gen[2962])
		); 

/******************* CELL 2963 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2963 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2867]),
			.N(gen[2868]),
			.NE(gen[2869]),

			.O(gen[2962]),
			.E(gen[2964]),

			.SO(gen[3057]),
			.S(gen[3058]),
			.SE(gen[3059]),

			.SELF(gen[2963]),
			.cell_state(gen[2963])
		); 

/******************* CELL 2964 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2964 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2868]),
			.N(gen[2869]),
			.NE(gen[2870]),

			.O(gen[2963]),
			.E(gen[2965]),

			.SO(gen[3058]),
			.S(gen[3059]),
			.SE(gen[3060]),

			.SELF(gen[2964]),
			.cell_state(gen[2964])
		); 

/******************* CELL 2965 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2965 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2869]),
			.N(gen[2870]),
			.NE(gen[2871]),

			.O(gen[2964]),
			.E(gen[2966]),

			.SO(gen[3059]),
			.S(gen[3060]),
			.SE(gen[3061]),

			.SELF(gen[2965]),
			.cell_state(gen[2965])
		); 

/******************* CELL 2966 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2966 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2870]),
			.N(gen[2871]),
			.NE(gen[2872]),

			.O(gen[2965]),
			.E(gen[2967]),

			.SO(gen[3060]),
			.S(gen[3061]),
			.SE(gen[3062]),

			.SELF(gen[2966]),
			.cell_state(gen[2966])
		); 

/******************* CELL 2967 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2967 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2871]),
			.N(gen[2872]),
			.NE(gen[2873]),

			.O(gen[2966]),
			.E(gen[2968]),

			.SO(gen[3061]),
			.S(gen[3062]),
			.SE(gen[3063]),

			.SELF(gen[2967]),
			.cell_state(gen[2967])
		); 

/******************* CELL 2968 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2968 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2872]),
			.N(gen[2873]),
			.NE(gen[2874]),

			.O(gen[2967]),
			.E(gen[2969]),

			.SO(gen[3062]),
			.S(gen[3063]),
			.SE(gen[3064]),

			.SELF(gen[2968]),
			.cell_state(gen[2968])
		); 

/******************* CELL 2969 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2969 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2873]),
			.N(gen[2874]),
			.NE(gen[2875]),

			.O(gen[2968]),
			.E(gen[2970]),

			.SO(gen[3063]),
			.S(gen[3064]),
			.SE(gen[3065]),

			.SELF(gen[2969]),
			.cell_state(gen[2969])
		); 

/******************* CELL 2970 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2970 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2874]),
			.N(gen[2875]),
			.NE(gen[2876]),

			.O(gen[2969]),
			.E(gen[2971]),

			.SO(gen[3064]),
			.S(gen[3065]),
			.SE(gen[3066]),

			.SELF(gen[2970]),
			.cell_state(gen[2970])
		); 

/******************* CELL 2971 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2971 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2875]),
			.N(gen[2876]),
			.NE(gen[2877]),

			.O(gen[2970]),
			.E(gen[2972]),

			.SO(gen[3065]),
			.S(gen[3066]),
			.SE(gen[3067]),

			.SELF(gen[2971]),
			.cell_state(gen[2971])
		); 

/******************* CELL 2972 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2972 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2876]),
			.N(gen[2877]),
			.NE(gen[2878]),

			.O(gen[2971]),
			.E(gen[2973]),

			.SO(gen[3066]),
			.S(gen[3067]),
			.SE(gen[3068]),

			.SELF(gen[2972]),
			.cell_state(gen[2972])
		); 

/******************* CELL 2973 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2973 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2877]),
			.N(gen[2878]),
			.NE(gen[2879]),

			.O(gen[2972]),
			.E(gen[2974]),

			.SO(gen[3067]),
			.S(gen[3068]),
			.SE(gen[3069]),

			.SELF(gen[2973]),
			.cell_state(gen[2973])
		); 

/******************* CELL 2974 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2974 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2878]),
			.N(gen[2879]),
			.NE(gen[2880]),

			.O(gen[2973]),
			.E(gen[2975]),

			.SO(gen[3068]),
			.S(gen[3069]),
			.SE(gen[3070]),

			.SELF(gen[2974]),
			.cell_state(gen[2974])
		); 

/******************* CELL 2975 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2975 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2879]),
			.N(gen[2880]),
			.NE(gen[2881]),

			.O(gen[2974]),
			.E(gen[2976]),

			.SO(gen[3069]),
			.S(gen[3070]),
			.SE(gen[3071]),

			.SELF(gen[2975]),
			.cell_state(gen[2975])
		); 

/******************* CELL 2976 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2976 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2880]),
			.N(gen[2881]),
			.NE(gen[2882]),

			.O(gen[2975]),
			.E(gen[2977]),

			.SO(gen[3070]),
			.S(gen[3071]),
			.SE(gen[3072]),

			.SELF(gen[2976]),
			.cell_state(gen[2976])
		); 

/******************* CELL 2977 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2977 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2881]),
			.N(gen[2882]),
			.NE(gen[2883]),

			.O(gen[2976]),
			.E(gen[2978]),

			.SO(gen[3071]),
			.S(gen[3072]),
			.SE(gen[3073]),

			.SELF(gen[2977]),
			.cell_state(gen[2977])
		); 

/******************* CELL 2978 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2978 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2882]),
			.N(gen[2883]),
			.NE(gen[2884]),

			.O(gen[2977]),
			.E(gen[2979]),

			.SO(gen[3072]),
			.S(gen[3073]),
			.SE(gen[3074]),

			.SELF(gen[2978]),
			.cell_state(gen[2978])
		); 

/******************* CELL 2979 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2979 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2883]),
			.N(gen[2884]),
			.NE(gen[2885]),

			.O(gen[2978]),
			.E(gen[2980]),

			.SO(gen[3073]),
			.S(gen[3074]),
			.SE(gen[3075]),

			.SELF(gen[2979]),
			.cell_state(gen[2979])
		); 

/******************* CELL 2980 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2980 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2884]),
			.N(gen[2885]),
			.NE(gen[2886]),

			.O(gen[2979]),
			.E(gen[2981]),

			.SO(gen[3074]),
			.S(gen[3075]),
			.SE(gen[3076]),

			.SELF(gen[2980]),
			.cell_state(gen[2980])
		); 

/******************* CELL 2981 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2981 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2885]),
			.N(gen[2886]),
			.NE(gen[2887]),

			.O(gen[2980]),
			.E(gen[2982]),

			.SO(gen[3075]),
			.S(gen[3076]),
			.SE(gen[3077]),

			.SELF(gen[2981]),
			.cell_state(gen[2981])
		); 

/******************* CELL 2982 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2982 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2886]),
			.N(gen[2887]),
			.NE(gen[2888]),

			.O(gen[2981]),
			.E(gen[2983]),

			.SO(gen[3076]),
			.S(gen[3077]),
			.SE(gen[3078]),

			.SELF(gen[2982]),
			.cell_state(gen[2982])
		); 

/******************* CELL 2983 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2983 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2887]),
			.N(gen[2888]),
			.NE(gen[2889]),

			.O(gen[2982]),
			.E(gen[2984]),

			.SO(gen[3077]),
			.S(gen[3078]),
			.SE(gen[3079]),

			.SELF(gen[2983]),
			.cell_state(gen[2983])
		); 

/******************* CELL 2984 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2984 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2888]),
			.N(gen[2889]),
			.NE(gen[2890]),

			.O(gen[2983]),
			.E(gen[2985]),

			.SO(gen[3078]),
			.S(gen[3079]),
			.SE(gen[3080]),

			.SELF(gen[2984]),
			.cell_state(gen[2984])
		); 

/******************* CELL 2985 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2985 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2889]),
			.N(gen[2890]),
			.NE(gen[2891]),

			.O(gen[2984]),
			.E(gen[2986]),

			.SO(gen[3079]),
			.S(gen[3080]),
			.SE(gen[3081]),

			.SELF(gen[2985]),
			.cell_state(gen[2985])
		); 

/******************* CELL 2986 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2986 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2890]),
			.N(gen[2891]),
			.NE(gen[2892]),

			.O(gen[2985]),
			.E(gen[2987]),

			.SO(gen[3080]),
			.S(gen[3081]),
			.SE(gen[3082]),

			.SELF(gen[2986]),
			.cell_state(gen[2986])
		); 

/******************* CELL 2987 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2987 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2891]),
			.N(gen[2892]),
			.NE(gen[2893]),

			.O(gen[2986]),
			.E(gen[2988]),

			.SO(gen[3081]),
			.S(gen[3082]),
			.SE(gen[3083]),

			.SELF(gen[2987]),
			.cell_state(gen[2987])
		); 

/******************* CELL 2988 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2988 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2892]),
			.N(gen[2893]),
			.NE(gen[2894]),

			.O(gen[2987]),
			.E(gen[2989]),

			.SO(gen[3082]),
			.S(gen[3083]),
			.SE(gen[3084]),

			.SELF(gen[2988]),
			.cell_state(gen[2988])
		); 

/******************* CELL 2989 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2989 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2893]),
			.N(gen[2894]),
			.NE(gen[2895]),

			.O(gen[2988]),
			.E(gen[2990]),

			.SO(gen[3083]),
			.S(gen[3084]),
			.SE(gen[3085]),

			.SELF(gen[2989]),
			.cell_state(gen[2989])
		); 

/******************* CELL 2990 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2990 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2894]),
			.N(gen[2895]),
			.NE(gen[2896]),

			.O(gen[2989]),
			.E(gen[2991]),

			.SO(gen[3084]),
			.S(gen[3085]),
			.SE(gen[3086]),

			.SELF(gen[2990]),
			.cell_state(gen[2990])
		); 

/******************* CELL 2991 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2991 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2895]),
			.N(gen[2896]),
			.NE(gen[2897]),

			.O(gen[2990]),
			.E(gen[2992]),

			.SO(gen[3085]),
			.S(gen[3086]),
			.SE(gen[3087]),

			.SELF(gen[2991]),
			.cell_state(gen[2991])
		); 

/******************* CELL 2992 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2992 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2896]),
			.N(gen[2897]),
			.NE(gen[2898]),

			.O(gen[2991]),
			.E(gen[2993]),

			.SO(gen[3086]),
			.S(gen[3087]),
			.SE(gen[3088]),

			.SELF(gen[2992]),
			.cell_state(gen[2992])
		); 

/******************* CELL 2993 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2993 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2897]),
			.N(gen[2898]),
			.NE(gen[2899]),

			.O(gen[2992]),
			.E(gen[2994]),

			.SO(gen[3087]),
			.S(gen[3088]),
			.SE(gen[3089]),

			.SELF(gen[2993]),
			.cell_state(gen[2993])
		); 

/******************* CELL 2994 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2994 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2898]),
			.N(gen[2899]),
			.NE(gen[2900]),

			.O(gen[2993]),
			.E(gen[2995]),

			.SO(gen[3088]),
			.S(gen[3089]),
			.SE(gen[3090]),

			.SELF(gen[2994]),
			.cell_state(gen[2994])
		); 

/******************* CELL 2995 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2995 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2899]),
			.N(gen[2900]),
			.NE(gen[2901]),

			.O(gen[2994]),
			.E(gen[2996]),

			.SO(gen[3089]),
			.S(gen[3090]),
			.SE(gen[3091]),

			.SELF(gen[2995]),
			.cell_state(gen[2995])
		); 

/******************* CELL 2996 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2996 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2900]),
			.N(gen[2901]),
			.NE(gen[2902]),

			.O(gen[2995]),
			.E(gen[2997]),

			.SO(gen[3090]),
			.S(gen[3091]),
			.SE(gen[3092]),

			.SELF(gen[2996]),
			.cell_state(gen[2996])
		); 

/******************* CELL 2997 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2997 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2901]),
			.N(gen[2902]),
			.NE(gen[2903]),

			.O(gen[2996]),
			.E(gen[2998]),

			.SO(gen[3091]),
			.S(gen[3092]),
			.SE(gen[3093]),

			.SELF(gen[2997]),
			.cell_state(gen[2997])
		); 

/******************* CELL 2998 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2998 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2902]),
			.N(gen[2903]),
			.NE(gen[2904]),

			.O(gen[2997]),
			.E(gen[2999]),

			.SO(gen[3092]),
			.S(gen[3093]),
			.SE(gen[3094]),

			.SELF(gen[2998]),
			.cell_state(gen[2998])
		); 

/******************* CELL 2999 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2999 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2903]),
			.N(gen[2904]),
			.NE(gen[2905]),

			.O(gen[2998]),
			.E(gen[3000]),

			.SO(gen[3093]),
			.S(gen[3094]),
			.SE(gen[3095]),

			.SELF(gen[2999]),
			.cell_state(gen[2999])
		); 

/******************* CELL 3000 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3000 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2904]),
			.N(gen[2905]),
			.NE(gen[2906]),

			.O(gen[2999]),
			.E(gen[3001]),

			.SO(gen[3094]),
			.S(gen[3095]),
			.SE(gen[3096]),

			.SELF(gen[3000]),
			.cell_state(gen[3000])
		); 

/******************* CELL 3001 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3001 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2905]),
			.N(gen[2906]),
			.NE(gen[2907]),

			.O(gen[3000]),
			.E(gen[3002]),

			.SO(gen[3095]),
			.S(gen[3096]),
			.SE(gen[3097]),

			.SELF(gen[3001]),
			.cell_state(gen[3001])
		); 

/******************* CELL 3002 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3002 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2906]),
			.N(gen[2907]),
			.NE(gen[2908]),

			.O(gen[3001]),
			.E(gen[3003]),

			.SO(gen[3096]),
			.S(gen[3097]),
			.SE(gen[3098]),

			.SELF(gen[3002]),
			.cell_state(gen[3002])
		); 

/******************* CELL 3003 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3003 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2907]),
			.N(gen[2908]),
			.NE(gen[2909]),

			.O(gen[3002]),
			.E(gen[3004]),

			.SO(gen[3097]),
			.S(gen[3098]),
			.SE(gen[3099]),

			.SELF(gen[3003]),
			.cell_state(gen[3003])
		); 

/******************* CELL 3004 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3004 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2908]),
			.N(gen[2909]),
			.NE(gen[2910]),

			.O(gen[3003]),
			.E(gen[3005]),

			.SO(gen[3098]),
			.S(gen[3099]),
			.SE(gen[3100]),

			.SELF(gen[3004]),
			.cell_state(gen[3004])
		); 

/******************* CELL 3005 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3005 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2909]),
			.N(gen[2910]),
			.NE(gen[2911]),

			.O(gen[3004]),
			.E(gen[3006]),

			.SO(gen[3099]),
			.S(gen[3100]),
			.SE(gen[3101]),

			.SELF(gen[3005]),
			.cell_state(gen[3005])
		); 

/******************* CELL 3006 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3006 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2910]),
			.N(gen[2911]),
			.NE(gen[2912]),

			.O(gen[3005]),
			.E(gen[3007]),

			.SO(gen[3100]),
			.S(gen[3101]),
			.SE(gen[3102]),

			.SELF(gen[3006]),
			.cell_state(gen[3006])
		); 

/******************* CELL 3007 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3007 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2911]),
			.N(gen[2912]),
			.NE(gen[2913]),

			.O(gen[3006]),
			.E(gen[3008]),

			.SO(gen[3101]),
			.S(gen[3102]),
			.SE(gen[3103]),

			.SELF(gen[3007]),
			.cell_state(gen[3007])
		); 

/******************* CELL 3008 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3008 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2912]),
			.N(gen[2913]),
			.NE(gen[2914]),

			.O(gen[3007]),
			.E(gen[3009]),

			.SO(gen[3102]),
			.S(gen[3103]),
			.SE(gen[3104]),

			.SELF(gen[3008]),
			.cell_state(gen[3008])
		); 

/******************* CELL 3009 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3009 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2913]),
			.N(gen[2914]),
			.NE(gen[2915]),

			.O(gen[3008]),
			.E(gen[3010]),

			.SO(gen[3103]),
			.S(gen[3104]),
			.SE(gen[3105]),

			.SELF(gen[3009]),
			.cell_state(gen[3009])
		); 

/******************* CELL 3010 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3010 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2914]),
			.N(gen[2915]),
			.NE(gen[2916]),

			.O(gen[3009]),
			.E(gen[3011]),

			.SO(gen[3104]),
			.S(gen[3105]),
			.SE(gen[3106]),

			.SELF(gen[3010]),
			.cell_state(gen[3010])
		); 

/******************* CELL 3011 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3011 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2915]),
			.N(gen[2916]),
			.NE(gen[2917]),

			.O(gen[3010]),
			.E(gen[3012]),

			.SO(gen[3105]),
			.S(gen[3106]),
			.SE(gen[3107]),

			.SELF(gen[3011]),
			.cell_state(gen[3011])
		); 

/******************* CELL 3012 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3012 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2916]),
			.N(gen[2917]),
			.NE(gen[2918]),

			.O(gen[3011]),
			.E(gen[3013]),

			.SO(gen[3106]),
			.S(gen[3107]),
			.SE(gen[3108]),

			.SELF(gen[3012]),
			.cell_state(gen[3012])
		); 

/******************* CELL 3013 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3013 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2917]),
			.N(gen[2918]),
			.NE(gen[2919]),

			.O(gen[3012]),
			.E(gen[3014]),

			.SO(gen[3107]),
			.S(gen[3108]),
			.SE(gen[3109]),

			.SELF(gen[3013]),
			.cell_state(gen[3013])
		); 

/******************* CELL 3014 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3014 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2918]),
			.N(gen[2919]),
			.NE(gen[2920]),

			.O(gen[3013]),
			.E(gen[3015]),

			.SO(gen[3108]),
			.S(gen[3109]),
			.SE(gen[3110]),

			.SELF(gen[3014]),
			.cell_state(gen[3014])
		); 

/******************* CELL 3015 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3015 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2919]),
			.N(gen[2920]),
			.NE(gen[2921]),

			.O(gen[3014]),
			.E(gen[3016]),

			.SO(gen[3109]),
			.S(gen[3110]),
			.SE(gen[3111]),

			.SELF(gen[3015]),
			.cell_state(gen[3015])
		); 

/******************* CELL 3016 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3016 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2920]),
			.N(gen[2921]),
			.NE(gen[2922]),

			.O(gen[3015]),
			.E(gen[3017]),

			.SO(gen[3110]),
			.S(gen[3111]),
			.SE(gen[3112]),

			.SELF(gen[3016]),
			.cell_state(gen[3016])
		); 

/******************* CELL 3017 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3017 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2921]),
			.N(gen[2922]),
			.NE(gen[2923]),

			.O(gen[3016]),
			.E(gen[3018]),

			.SO(gen[3111]),
			.S(gen[3112]),
			.SE(gen[3113]),

			.SELF(gen[3017]),
			.cell_state(gen[3017])
		); 

/******************* CELL 3018 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3018 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2922]),
			.N(gen[2923]),
			.NE(gen[2924]),

			.O(gen[3017]),
			.E(gen[3019]),

			.SO(gen[3112]),
			.S(gen[3113]),
			.SE(gen[3114]),

			.SELF(gen[3018]),
			.cell_state(gen[3018])
		); 

/******************* CELL 3019 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3019 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2923]),
			.N(gen[2924]),
			.NE(gen[2925]),

			.O(gen[3018]),
			.E(gen[3020]),

			.SO(gen[3113]),
			.S(gen[3114]),
			.SE(gen[3115]),

			.SELF(gen[3019]),
			.cell_state(gen[3019])
		); 

/******************* CELL 3020 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3020 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2924]),
			.N(gen[2925]),
			.NE(gen[2926]),

			.O(gen[3019]),
			.E(gen[3021]),

			.SO(gen[3114]),
			.S(gen[3115]),
			.SE(gen[3116]),

			.SELF(gen[3020]),
			.cell_state(gen[3020])
		); 

/******************* CELL 3021 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3021 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2925]),
			.N(gen[2926]),
			.NE(gen[2927]),

			.O(gen[3020]),
			.E(gen[3022]),

			.SO(gen[3115]),
			.S(gen[3116]),
			.SE(gen[3117]),

			.SELF(gen[3021]),
			.cell_state(gen[3021])
		); 

/******************* CELL 3022 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3022 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2926]),
			.N(gen[2927]),
			.NE(gen[2928]),

			.O(gen[3021]),
			.E(gen[3023]),

			.SO(gen[3116]),
			.S(gen[3117]),
			.SE(gen[3118]),

			.SELF(gen[3022]),
			.cell_state(gen[3022])
		); 

/******************* CELL 3023 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3023 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2927]),
			.N(gen[2928]),
			.NE(gen[2929]),

			.O(gen[3022]),
			.E(gen[3024]),

			.SO(gen[3117]),
			.S(gen[3118]),
			.SE(gen[3119]),

			.SELF(gen[3023]),
			.cell_state(gen[3023])
		); 

/******************* CELL 3024 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3024 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2928]),
			.N(gen[2929]),
			.NE(gen[2930]),

			.O(gen[3023]),
			.E(gen[3025]),

			.SO(gen[3118]),
			.S(gen[3119]),
			.SE(gen[3120]),

			.SELF(gen[3024]),
			.cell_state(gen[3024])
		); 

/******************* CELL 3025 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3025 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2929]),
			.N(gen[2930]),
			.NE(gen[2931]),

			.O(gen[3024]),
			.E(gen[3026]),

			.SO(gen[3119]),
			.S(gen[3120]),
			.SE(gen[3121]),

			.SELF(gen[3025]),
			.cell_state(gen[3025])
		); 

/******************* CELL 3026 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3026 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2930]),
			.N(gen[2931]),
			.NE(gen[2932]),

			.O(gen[3025]),
			.E(gen[3027]),

			.SO(gen[3120]),
			.S(gen[3121]),
			.SE(gen[3122]),

			.SELF(gen[3026]),
			.cell_state(gen[3026])
		); 

/******************* CELL 3027 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3027 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2931]),
			.N(gen[2932]),
			.NE(gen[2933]),

			.O(gen[3026]),
			.E(gen[3028]),

			.SO(gen[3121]),
			.S(gen[3122]),
			.SE(gen[3123]),

			.SELF(gen[3027]),
			.cell_state(gen[3027])
		); 

/******************* CELL 3028 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3028 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2932]),
			.N(gen[2933]),
			.NE(gen[2934]),

			.O(gen[3027]),
			.E(gen[3029]),

			.SO(gen[3122]),
			.S(gen[3123]),
			.SE(gen[3124]),

			.SELF(gen[3028]),
			.cell_state(gen[3028])
		); 

/******************* CELL 3029 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3029 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2933]),
			.N(gen[2934]),
			.NE(gen[2935]),

			.O(gen[3028]),
			.E(gen[3030]),

			.SO(gen[3123]),
			.S(gen[3124]),
			.SE(gen[3125]),

			.SELF(gen[3029]),
			.cell_state(gen[3029])
		); 

/******************* CELL 3030 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3030 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2934]),
			.N(gen[2935]),
			.NE(gen[2936]),

			.O(gen[3029]),
			.E(gen[3031]),

			.SO(gen[3124]),
			.S(gen[3125]),
			.SE(gen[3126]),

			.SELF(gen[3030]),
			.cell_state(gen[3030])
		); 

/******************* CELL 3031 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3031 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2935]),
			.N(gen[2936]),
			.NE(gen[2937]),

			.O(gen[3030]),
			.E(gen[3032]),

			.SO(gen[3125]),
			.S(gen[3126]),
			.SE(gen[3127]),

			.SELF(gen[3031]),
			.cell_state(gen[3031])
		); 

/******************* CELL 3032 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3032 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2936]),
			.N(gen[2937]),
			.NE(gen[2938]),

			.O(gen[3031]),
			.E(gen[3033]),

			.SO(gen[3126]),
			.S(gen[3127]),
			.SE(gen[3128]),

			.SELF(gen[3032]),
			.cell_state(gen[3032])
		); 

/******************* CELL 3033 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3033 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2937]),
			.N(gen[2938]),
			.NE(gen[2939]),

			.O(gen[3032]),
			.E(gen[3034]),

			.SO(gen[3127]),
			.S(gen[3128]),
			.SE(gen[3129]),

			.SELF(gen[3033]),
			.cell_state(gen[3033])
		); 

/******************* CELL 3034 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3034 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2938]),
			.N(gen[2939]),
			.NE(gen[2940]),

			.O(gen[3033]),
			.E(gen[3035]),

			.SO(gen[3128]),
			.S(gen[3129]),
			.SE(gen[3130]),

			.SELF(gen[3034]),
			.cell_state(gen[3034])
		); 

/******************* CELL 3035 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3035 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2939]),
			.N(gen[2940]),
			.NE(gen[2941]),

			.O(gen[3034]),
			.E(gen[3036]),

			.SO(gen[3129]),
			.S(gen[3130]),
			.SE(gen[3131]),

			.SELF(gen[3035]),
			.cell_state(gen[3035])
		); 

/******************* CELL 3036 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3036 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2940]),
			.N(gen[2941]),
			.NE(gen[2942]),

			.O(gen[3035]),
			.E(gen[3037]),

			.SO(gen[3130]),
			.S(gen[3131]),
			.SE(gen[3132]),

			.SELF(gen[3036]),
			.cell_state(gen[3036])
		); 

/******************* CELL 3037 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3037 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2941]),
			.N(gen[2942]),
			.NE(gen[2943]),

			.O(gen[3036]),
			.E(gen[3038]),

			.SO(gen[3131]),
			.S(gen[3132]),
			.SE(gen[3133]),

			.SELF(gen[3037]),
			.cell_state(gen[3037])
		); 

/******************* CELL 3038 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3038 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2942]),
			.N(gen[2943]),
			.NE(gen[2944]),

			.O(gen[3037]),
			.E(gen[3039]),

			.SO(gen[3132]),
			.S(gen[3133]),
			.SE(gen[3134]),

			.SELF(gen[3038]),
			.cell_state(gen[3038])
		); 

/******************* CELL 3039 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3039 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2943]),
			.N(gen[2944]),
			.NE(gen[2943]),

			.O(gen[3038]),
			.E(gen[3038]),

			.SO(gen[3133]),
			.S(gen[3134]),
			.SE(gen[3133]),

			.SELF(gen[3039]),
			.cell_state(gen[3039])
		); 

/******************* CELL 3040 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3040 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2946]),
			.N(gen[2945]),
			.NE(gen[2946]),

			.O(gen[3041]),
			.E(gen[3041]),

			.SO(gen[3136]),
			.S(gen[3135]),
			.SE(gen[3136]),

			.SELF(gen[3040]),
			.cell_state(gen[3040])
		); 

/******************* CELL 3041 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3041 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2945]),
			.N(gen[2946]),
			.NE(gen[2947]),

			.O(gen[3040]),
			.E(gen[3042]),

			.SO(gen[3135]),
			.S(gen[3136]),
			.SE(gen[3137]),

			.SELF(gen[3041]),
			.cell_state(gen[3041])
		); 

/******************* CELL 3042 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3042 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2946]),
			.N(gen[2947]),
			.NE(gen[2948]),

			.O(gen[3041]),
			.E(gen[3043]),

			.SO(gen[3136]),
			.S(gen[3137]),
			.SE(gen[3138]),

			.SELF(gen[3042]),
			.cell_state(gen[3042])
		); 

/******************* CELL 3043 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3043 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2947]),
			.N(gen[2948]),
			.NE(gen[2949]),

			.O(gen[3042]),
			.E(gen[3044]),

			.SO(gen[3137]),
			.S(gen[3138]),
			.SE(gen[3139]),

			.SELF(gen[3043]),
			.cell_state(gen[3043])
		); 

/******************* CELL 3044 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3044 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2948]),
			.N(gen[2949]),
			.NE(gen[2950]),

			.O(gen[3043]),
			.E(gen[3045]),

			.SO(gen[3138]),
			.S(gen[3139]),
			.SE(gen[3140]),

			.SELF(gen[3044]),
			.cell_state(gen[3044])
		); 

/******************* CELL 3045 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3045 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2949]),
			.N(gen[2950]),
			.NE(gen[2951]),

			.O(gen[3044]),
			.E(gen[3046]),

			.SO(gen[3139]),
			.S(gen[3140]),
			.SE(gen[3141]),

			.SELF(gen[3045]),
			.cell_state(gen[3045])
		); 

/******************* CELL 3046 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3046 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2950]),
			.N(gen[2951]),
			.NE(gen[2952]),

			.O(gen[3045]),
			.E(gen[3047]),

			.SO(gen[3140]),
			.S(gen[3141]),
			.SE(gen[3142]),

			.SELF(gen[3046]),
			.cell_state(gen[3046])
		); 

/******************* CELL 3047 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3047 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2951]),
			.N(gen[2952]),
			.NE(gen[2953]),

			.O(gen[3046]),
			.E(gen[3048]),

			.SO(gen[3141]),
			.S(gen[3142]),
			.SE(gen[3143]),

			.SELF(gen[3047]),
			.cell_state(gen[3047])
		); 

/******************* CELL 3048 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3048 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2952]),
			.N(gen[2953]),
			.NE(gen[2954]),

			.O(gen[3047]),
			.E(gen[3049]),

			.SO(gen[3142]),
			.S(gen[3143]),
			.SE(gen[3144]),

			.SELF(gen[3048]),
			.cell_state(gen[3048])
		); 

/******************* CELL 3049 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3049 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2953]),
			.N(gen[2954]),
			.NE(gen[2955]),

			.O(gen[3048]),
			.E(gen[3050]),

			.SO(gen[3143]),
			.S(gen[3144]),
			.SE(gen[3145]),

			.SELF(gen[3049]),
			.cell_state(gen[3049])
		); 

/******************* CELL 3050 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3050 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2954]),
			.N(gen[2955]),
			.NE(gen[2956]),

			.O(gen[3049]),
			.E(gen[3051]),

			.SO(gen[3144]),
			.S(gen[3145]),
			.SE(gen[3146]),

			.SELF(gen[3050]),
			.cell_state(gen[3050])
		); 

/******************* CELL 3051 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3051 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2955]),
			.N(gen[2956]),
			.NE(gen[2957]),

			.O(gen[3050]),
			.E(gen[3052]),

			.SO(gen[3145]),
			.S(gen[3146]),
			.SE(gen[3147]),

			.SELF(gen[3051]),
			.cell_state(gen[3051])
		); 

/******************* CELL 3052 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3052 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2956]),
			.N(gen[2957]),
			.NE(gen[2958]),

			.O(gen[3051]),
			.E(gen[3053]),

			.SO(gen[3146]),
			.S(gen[3147]),
			.SE(gen[3148]),

			.SELF(gen[3052]),
			.cell_state(gen[3052])
		); 

/******************* CELL 3053 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3053 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2957]),
			.N(gen[2958]),
			.NE(gen[2959]),

			.O(gen[3052]),
			.E(gen[3054]),

			.SO(gen[3147]),
			.S(gen[3148]),
			.SE(gen[3149]),

			.SELF(gen[3053]),
			.cell_state(gen[3053])
		); 

/******************* CELL 3054 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3054 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2958]),
			.N(gen[2959]),
			.NE(gen[2960]),

			.O(gen[3053]),
			.E(gen[3055]),

			.SO(gen[3148]),
			.S(gen[3149]),
			.SE(gen[3150]),

			.SELF(gen[3054]),
			.cell_state(gen[3054])
		); 

/******************* CELL 3055 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3055 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2959]),
			.N(gen[2960]),
			.NE(gen[2961]),

			.O(gen[3054]),
			.E(gen[3056]),

			.SO(gen[3149]),
			.S(gen[3150]),
			.SE(gen[3151]),

			.SELF(gen[3055]),
			.cell_state(gen[3055])
		); 

/******************* CELL 3056 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3056 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2960]),
			.N(gen[2961]),
			.NE(gen[2962]),

			.O(gen[3055]),
			.E(gen[3057]),

			.SO(gen[3150]),
			.S(gen[3151]),
			.SE(gen[3152]),

			.SELF(gen[3056]),
			.cell_state(gen[3056])
		); 

/******************* CELL 3057 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3057 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2961]),
			.N(gen[2962]),
			.NE(gen[2963]),

			.O(gen[3056]),
			.E(gen[3058]),

			.SO(gen[3151]),
			.S(gen[3152]),
			.SE(gen[3153]),

			.SELF(gen[3057]),
			.cell_state(gen[3057])
		); 

/******************* CELL 3058 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3058 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2962]),
			.N(gen[2963]),
			.NE(gen[2964]),

			.O(gen[3057]),
			.E(gen[3059]),

			.SO(gen[3152]),
			.S(gen[3153]),
			.SE(gen[3154]),

			.SELF(gen[3058]),
			.cell_state(gen[3058])
		); 

/******************* CELL 3059 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3059 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2963]),
			.N(gen[2964]),
			.NE(gen[2965]),

			.O(gen[3058]),
			.E(gen[3060]),

			.SO(gen[3153]),
			.S(gen[3154]),
			.SE(gen[3155]),

			.SELF(gen[3059]),
			.cell_state(gen[3059])
		); 

/******************* CELL 3060 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3060 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2964]),
			.N(gen[2965]),
			.NE(gen[2966]),

			.O(gen[3059]),
			.E(gen[3061]),

			.SO(gen[3154]),
			.S(gen[3155]),
			.SE(gen[3156]),

			.SELF(gen[3060]),
			.cell_state(gen[3060])
		); 

/******************* CELL 3061 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3061 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2965]),
			.N(gen[2966]),
			.NE(gen[2967]),

			.O(gen[3060]),
			.E(gen[3062]),

			.SO(gen[3155]),
			.S(gen[3156]),
			.SE(gen[3157]),

			.SELF(gen[3061]),
			.cell_state(gen[3061])
		); 

/******************* CELL 3062 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3062 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2966]),
			.N(gen[2967]),
			.NE(gen[2968]),

			.O(gen[3061]),
			.E(gen[3063]),

			.SO(gen[3156]),
			.S(gen[3157]),
			.SE(gen[3158]),

			.SELF(gen[3062]),
			.cell_state(gen[3062])
		); 

/******************* CELL 3063 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3063 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2967]),
			.N(gen[2968]),
			.NE(gen[2969]),

			.O(gen[3062]),
			.E(gen[3064]),

			.SO(gen[3157]),
			.S(gen[3158]),
			.SE(gen[3159]),

			.SELF(gen[3063]),
			.cell_state(gen[3063])
		); 

/******************* CELL 3064 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3064 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2968]),
			.N(gen[2969]),
			.NE(gen[2970]),

			.O(gen[3063]),
			.E(gen[3065]),

			.SO(gen[3158]),
			.S(gen[3159]),
			.SE(gen[3160]),

			.SELF(gen[3064]),
			.cell_state(gen[3064])
		); 

/******************* CELL 3065 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3065 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2969]),
			.N(gen[2970]),
			.NE(gen[2971]),

			.O(gen[3064]),
			.E(gen[3066]),

			.SO(gen[3159]),
			.S(gen[3160]),
			.SE(gen[3161]),

			.SELF(gen[3065]),
			.cell_state(gen[3065])
		); 

/******************* CELL 3066 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3066 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2970]),
			.N(gen[2971]),
			.NE(gen[2972]),

			.O(gen[3065]),
			.E(gen[3067]),

			.SO(gen[3160]),
			.S(gen[3161]),
			.SE(gen[3162]),

			.SELF(gen[3066]),
			.cell_state(gen[3066])
		); 

/******************* CELL 3067 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3067 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2971]),
			.N(gen[2972]),
			.NE(gen[2973]),

			.O(gen[3066]),
			.E(gen[3068]),

			.SO(gen[3161]),
			.S(gen[3162]),
			.SE(gen[3163]),

			.SELF(gen[3067]),
			.cell_state(gen[3067])
		); 

/******************* CELL 3068 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3068 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2972]),
			.N(gen[2973]),
			.NE(gen[2974]),

			.O(gen[3067]),
			.E(gen[3069]),

			.SO(gen[3162]),
			.S(gen[3163]),
			.SE(gen[3164]),

			.SELF(gen[3068]),
			.cell_state(gen[3068])
		); 

/******************* CELL 3069 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3069 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2973]),
			.N(gen[2974]),
			.NE(gen[2975]),

			.O(gen[3068]),
			.E(gen[3070]),

			.SO(gen[3163]),
			.S(gen[3164]),
			.SE(gen[3165]),

			.SELF(gen[3069]),
			.cell_state(gen[3069])
		); 

/******************* CELL 3070 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3070 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2974]),
			.N(gen[2975]),
			.NE(gen[2976]),

			.O(gen[3069]),
			.E(gen[3071]),

			.SO(gen[3164]),
			.S(gen[3165]),
			.SE(gen[3166]),

			.SELF(gen[3070]),
			.cell_state(gen[3070])
		); 

/******************* CELL 3071 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3071 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2975]),
			.N(gen[2976]),
			.NE(gen[2977]),

			.O(gen[3070]),
			.E(gen[3072]),

			.SO(gen[3165]),
			.S(gen[3166]),
			.SE(gen[3167]),

			.SELF(gen[3071]),
			.cell_state(gen[3071])
		); 

/******************* CELL 3072 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3072 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2976]),
			.N(gen[2977]),
			.NE(gen[2978]),

			.O(gen[3071]),
			.E(gen[3073]),

			.SO(gen[3166]),
			.S(gen[3167]),
			.SE(gen[3168]),

			.SELF(gen[3072]),
			.cell_state(gen[3072])
		); 

/******************* CELL 3073 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3073 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2977]),
			.N(gen[2978]),
			.NE(gen[2979]),

			.O(gen[3072]),
			.E(gen[3074]),

			.SO(gen[3167]),
			.S(gen[3168]),
			.SE(gen[3169]),

			.SELF(gen[3073]),
			.cell_state(gen[3073])
		); 

/******************* CELL 3074 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3074 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2978]),
			.N(gen[2979]),
			.NE(gen[2980]),

			.O(gen[3073]),
			.E(gen[3075]),

			.SO(gen[3168]),
			.S(gen[3169]),
			.SE(gen[3170]),

			.SELF(gen[3074]),
			.cell_state(gen[3074])
		); 

/******************* CELL 3075 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3075 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2979]),
			.N(gen[2980]),
			.NE(gen[2981]),

			.O(gen[3074]),
			.E(gen[3076]),

			.SO(gen[3169]),
			.S(gen[3170]),
			.SE(gen[3171]),

			.SELF(gen[3075]),
			.cell_state(gen[3075])
		); 

/******************* CELL 3076 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3076 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2980]),
			.N(gen[2981]),
			.NE(gen[2982]),

			.O(gen[3075]),
			.E(gen[3077]),

			.SO(gen[3170]),
			.S(gen[3171]),
			.SE(gen[3172]),

			.SELF(gen[3076]),
			.cell_state(gen[3076])
		); 

/******************* CELL 3077 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3077 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2981]),
			.N(gen[2982]),
			.NE(gen[2983]),

			.O(gen[3076]),
			.E(gen[3078]),

			.SO(gen[3171]),
			.S(gen[3172]),
			.SE(gen[3173]),

			.SELF(gen[3077]),
			.cell_state(gen[3077])
		); 

/******************* CELL 3078 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3078 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2982]),
			.N(gen[2983]),
			.NE(gen[2984]),

			.O(gen[3077]),
			.E(gen[3079]),

			.SO(gen[3172]),
			.S(gen[3173]),
			.SE(gen[3174]),

			.SELF(gen[3078]),
			.cell_state(gen[3078])
		); 

/******************* CELL 3079 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3079 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2983]),
			.N(gen[2984]),
			.NE(gen[2985]),

			.O(gen[3078]),
			.E(gen[3080]),

			.SO(gen[3173]),
			.S(gen[3174]),
			.SE(gen[3175]),

			.SELF(gen[3079]),
			.cell_state(gen[3079])
		); 

/******************* CELL 3080 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3080 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2984]),
			.N(gen[2985]),
			.NE(gen[2986]),

			.O(gen[3079]),
			.E(gen[3081]),

			.SO(gen[3174]),
			.S(gen[3175]),
			.SE(gen[3176]),

			.SELF(gen[3080]),
			.cell_state(gen[3080])
		); 

/******************* CELL 3081 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3081 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2985]),
			.N(gen[2986]),
			.NE(gen[2987]),

			.O(gen[3080]),
			.E(gen[3082]),

			.SO(gen[3175]),
			.S(gen[3176]),
			.SE(gen[3177]),

			.SELF(gen[3081]),
			.cell_state(gen[3081])
		); 

/******************* CELL 3082 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3082 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2986]),
			.N(gen[2987]),
			.NE(gen[2988]),

			.O(gen[3081]),
			.E(gen[3083]),

			.SO(gen[3176]),
			.S(gen[3177]),
			.SE(gen[3178]),

			.SELF(gen[3082]),
			.cell_state(gen[3082])
		); 

/******************* CELL 3083 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3083 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2987]),
			.N(gen[2988]),
			.NE(gen[2989]),

			.O(gen[3082]),
			.E(gen[3084]),

			.SO(gen[3177]),
			.S(gen[3178]),
			.SE(gen[3179]),

			.SELF(gen[3083]),
			.cell_state(gen[3083])
		); 

/******************* CELL 3084 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3084 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2988]),
			.N(gen[2989]),
			.NE(gen[2990]),

			.O(gen[3083]),
			.E(gen[3085]),

			.SO(gen[3178]),
			.S(gen[3179]),
			.SE(gen[3180]),

			.SELF(gen[3084]),
			.cell_state(gen[3084])
		); 

/******************* CELL 3085 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3085 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2989]),
			.N(gen[2990]),
			.NE(gen[2991]),

			.O(gen[3084]),
			.E(gen[3086]),

			.SO(gen[3179]),
			.S(gen[3180]),
			.SE(gen[3181]),

			.SELF(gen[3085]),
			.cell_state(gen[3085])
		); 

/******************* CELL 3086 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3086 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2990]),
			.N(gen[2991]),
			.NE(gen[2992]),

			.O(gen[3085]),
			.E(gen[3087]),

			.SO(gen[3180]),
			.S(gen[3181]),
			.SE(gen[3182]),

			.SELF(gen[3086]),
			.cell_state(gen[3086])
		); 

/******************* CELL 3087 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3087 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2991]),
			.N(gen[2992]),
			.NE(gen[2993]),

			.O(gen[3086]),
			.E(gen[3088]),

			.SO(gen[3181]),
			.S(gen[3182]),
			.SE(gen[3183]),

			.SELF(gen[3087]),
			.cell_state(gen[3087])
		); 

/******************* CELL 3088 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3088 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2992]),
			.N(gen[2993]),
			.NE(gen[2994]),

			.O(gen[3087]),
			.E(gen[3089]),

			.SO(gen[3182]),
			.S(gen[3183]),
			.SE(gen[3184]),

			.SELF(gen[3088]),
			.cell_state(gen[3088])
		); 

/******************* CELL 3089 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3089 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2993]),
			.N(gen[2994]),
			.NE(gen[2995]),

			.O(gen[3088]),
			.E(gen[3090]),

			.SO(gen[3183]),
			.S(gen[3184]),
			.SE(gen[3185]),

			.SELF(gen[3089]),
			.cell_state(gen[3089])
		); 

/******************* CELL 3090 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3090 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2994]),
			.N(gen[2995]),
			.NE(gen[2996]),

			.O(gen[3089]),
			.E(gen[3091]),

			.SO(gen[3184]),
			.S(gen[3185]),
			.SE(gen[3186]),

			.SELF(gen[3090]),
			.cell_state(gen[3090])
		); 

/******************* CELL 3091 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3091 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2995]),
			.N(gen[2996]),
			.NE(gen[2997]),

			.O(gen[3090]),
			.E(gen[3092]),

			.SO(gen[3185]),
			.S(gen[3186]),
			.SE(gen[3187]),

			.SELF(gen[3091]),
			.cell_state(gen[3091])
		); 

/******************* CELL 3092 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3092 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2996]),
			.N(gen[2997]),
			.NE(gen[2998]),

			.O(gen[3091]),
			.E(gen[3093]),

			.SO(gen[3186]),
			.S(gen[3187]),
			.SE(gen[3188]),

			.SELF(gen[3092]),
			.cell_state(gen[3092])
		); 

/******************* CELL 3093 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3093 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2997]),
			.N(gen[2998]),
			.NE(gen[2999]),

			.O(gen[3092]),
			.E(gen[3094]),

			.SO(gen[3187]),
			.S(gen[3188]),
			.SE(gen[3189]),

			.SELF(gen[3093]),
			.cell_state(gen[3093])
		); 

/******************* CELL 3094 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3094 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2998]),
			.N(gen[2999]),
			.NE(gen[3000]),

			.O(gen[3093]),
			.E(gen[3095]),

			.SO(gen[3188]),
			.S(gen[3189]),
			.SE(gen[3190]),

			.SELF(gen[3094]),
			.cell_state(gen[3094])
		); 

/******************* CELL 3095 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3095 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2999]),
			.N(gen[3000]),
			.NE(gen[3001]),

			.O(gen[3094]),
			.E(gen[3096]),

			.SO(gen[3189]),
			.S(gen[3190]),
			.SE(gen[3191]),

			.SELF(gen[3095]),
			.cell_state(gen[3095])
		); 

/******************* CELL 3096 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3096 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3000]),
			.N(gen[3001]),
			.NE(gen[3002]),

			.O(gen[3095]),
			.E(gen[3097]),

			.SO(gen[3190]),
			.S(gen[3191]),
			.SE(gen[3192]),

			.SELF(gen[3096]),
			.cell_state(gen[3096])
		); 

/******************* CELL 3097 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3097 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3001]),
			.N(gen[3002]),
			.NE(gen[3003]),

			.O(gen[3096]),
			.E(gen[3098]),

			.SO(gen[3191]),
			.S(gen[3192]),
			.SE(gen[3193]),

			.SELF(gen[3097]),
			.cell_state(gen[3097])
		); 

/******************* CELL 3098 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3098 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3002]),
			.N(gen[3003]),
			.NE(gen[3004]),

			.O(gen[3097]),
			.E(gen[3099]),

			.SO(gen[3192]),
			.S(gen[3193]),
			.SE(gen[3194]),

			.SELF(gen[3098]),
			.cell_state(gen[3098])
		); 

/******************* CELL 3099 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3099 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3003]),
			.N(gen[3004]),
			.NE(gen[3005]),

			.O(gen[3098]),
			.E(gen[3100]),

			.SO(gen[3193]),
			.S(gen[3194]),
			.SE(gen[3195]),

			.SELF(gen[3099]),
			.cell_state(gen[3099])
		); 

/******************* CELL 3100 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3100 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3004]),
			.N(gen[3005]),
			.NE(gen[3006]),

			.O(gen[3099]),
			.E(gen[3101]),

			.SO(gen[3194]),
			.S(gen[3195]),
			.SE(gen[3196]),

			.SELF(gen[3100]),
			.cell_state(gen[3100])
		); 

/******************* CELL 3101 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3101 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3005]),
			.N(gen[3006]),
			.NE(gen[3007]),

			.O(gen[3100]),
			.E(gen[3102]),

			.SO(gen[3195]),
			.S(gen[3196]),
			.SE(gen[3197]),

			.SELF(gen[3101]),
			.cell_state(gen[3101])
		); 

/******************* CELL 3102 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3102 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3006]),
			.N(gen[3007]),
			.NE(gen[3008]),

			.O(gen[3101]),
			.E(gen[3103]),

			.SO(gen[3196]),
			.S(gen[3197]),
			.SE(gen[3198]),

			.SELF(gen[3102]),
			.cell_state(gen[3102])
		); 

/******************* CELL 3103 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3103 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3007]),
			.N(gen[3008]),
			.NE(gen[3009]),

			.O(gen[3102]),
			.E(gen[3104]),

			.SO(gen[3197]),
			.S(gen[3198]),
			.SE(gen[3199]),

			.SELF(gen[3103]),
			.cell_state(gen[3103])
		); 

/******************* CELL 3104 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3104 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3008]),
			.N(gen[3009]),
			.NE(gen[3010]),

			.O(gen[3103]),
			.E(gen[3105]),

			.SO(gen[3198]),
			.S(gen[3199]),
			.SE(gen[3200]),

			.SELF(gen[3104]),
			.cell_state(gen[3104])
		); 

/******************* CELL 3105 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3105 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3009]),
			.N(gen[3010]),
			.NE(gen[3011]),

			.O(gen[3104]),
			.E(gen[3106]),

			.SO(gen[3199]),
			.S(gen[3200]),
			.SE(gen[3201]),

			.SELF(gen[3105]),
			.cell_state(gen[3105])
		); 

/******************* CELL 3106 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3106 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3010]),
			.N(gen[3011]),
			.NE(gen[3012]),

			.O(gen[3105]),
			.E(gen[3107]),

			.SO(gen[3200]),
			.S(gen[3201]),
			.SE(gen[3202]),

			.SELF(gen[3106]),
			.cell_state(gen[3106])
		); 

/******************* CELL 3107 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3107 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3011]),
			.N(gen[3012]),
			.NE(gen[3013]),

			.O(gen[3106]),
			.E(gen[3108]),

			.SO(gen[3201]),
			.S(gen[3202]),
			.SE(gen[3203]),

			.SELF(gen[3107]),
			.cell_state(gen[3107])
		); 

/******************* CELL 3108 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3108 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3012]),
			.N(gen[3013]),
			.NE(gen[3014]),

			.O(gen[3107]),
			.E(gen[3109]),

			.SO(gen[3202]),
			.S(gen[3203]),
			.SE(gen[3204]),

			.SELF(gen[3108]),
			.cell_state(gen[3108])
		); 

/******************* CELL 3109 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3109 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3013]),
			.N(gen[3014]),
			.NE(gen[3015]),

			.O(gen[3108]),
			.E(gen[3110]),

			.SO(gen[3203]),
			.S(gen[3204]),
			.SE(gen[3205]),

			.SELF(gen[3109]),
			.cell_state(gen[3109])
		); 

/******************* CELL 3110 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3110 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3014]),
			.N(gen[3015]),
			.NE(gen[3016]),

			.O(gen[3109]),
			.E(gen[3111]),

			.SO(gen[3204]),
			.S(gen[3205]),
			.SE(gen[3206]),

			.SELF(gen[3110]),
			.cell_state(gen[3110])
		); 

/******************* CELL 3111 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3111 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3015]),
			.N(gen[3016]),
			.NE(gen[3017]),

			.O(gen[3110]),
			.E(gen[3112]),

			.SO(gen[3205]),
			.S(gen[3206]),
			.SE(gen[3207]),

			.SELF(gen[3111]),
			.cell_state(gen[3111])
		); 

/******************* CELL 3112 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3112 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3016]),
			.N(gen[3017]),
			.NE(gen[3018]),

			.O(gen[3111]),
			.E(gen[3113]),

			.SO(gen[3206]),
			.S(gen[3207]),
			.SE(gen[3208]),

			.SELF(gen[3112]),
			.cell_state(gen[3112])
		); 

/******************* CELL 3113 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3113 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3017]),
			.N(gen[3018]),
			.NE(gen[3019]),

			.O(gen[3112]),
			.E(gen[3114]),

			.SO(gen[3207]),
			.S(gen[3208]),
			.SE(gen[3209]),

			.SELF(gen[3113]),
			.cell_state(gen[3113])
		); 

/******************* CELL 3114 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3114 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3018]),
			.N(gen[3019]),
			.NE(gen[3020]),

			.O(gen[3113]),
			.E(gen[3115]),

			.SO(gen[3208]),
			.S(gen[3209]),
			.SE(gen[3210]),

			.SELF(gen[3114]),
			.cell_state(gen[3114])
		); 

/******************* CELL 3115 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3115 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3019]),
			.N(gen[3020]),
			.NE(gen[3021]),

			.O(gen[3114]),
			.E(gen[3116]),

			.SO(gen[3209]),
			.S(gen[3210]),
			.SE(gen[3211]),

			.SELF(gen[3115]),
			.cell_state(gen[3115])
		); 

/******************* CELL 3116 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3116 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3020]),
			.N(gen[3021]),
			.NE(gen[3022]),

			.O(gen[3115]),
			.E(gen[3117]),

			.SO(gen[3210]),
			.S(gen[3211]),
			.SE(gen[3212]),

			.SELF(gen[3116]),
			.cell_state(gen[3116])
		); 

/******************* CELL 3117 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3117 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3021]),
			.N(gen[3022]),
			.NE(gen[3023]),

			.O(gen[3116]),
			.E(gen[3118]),

			.SO(gen[3211]),
			.S(gen[3212]),
			.SE(gen[3213]),

			.SELF(gen[3117]),
			.cell_state(gen[3117])
		); 

/******************* CELL 3118 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3118 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3022]),
			.N(gen[3023]),
			.NE(gen[3024]),

			.O(gen[3117]),
			.E(gen[3119]),

			.SO(gen[3212]),
			.S(gen[3213]),
			.SE(gen[3214]),

			.SELF(gen[3118]),
			.cell_state(gen[3118])
		); 

/******************* CELL 3119 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3119 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3023]),
			.N(gen[3024]),
			.NE(gen[3025]),

			.O(gen[3118]),
			.E(gen[3120]),

			.SO(gen[3213]),
			.S(gen[3214]),
			.SE(gen[3215]),

			.SELF(gen[3119]),
			.cell_state(gen[3119])
		); 

/******************* CELL 3120 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3120 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3024]),
			.N(gen[3025]),
			.NE(gen[3026]),

			.O(gen[3119]),
			.E(gen[3121]),

			.SO(gen[3214]),
			.S(gen[3215]),
			.SE(gen[3216]),

			.SELF(gen[3120]),
			.cell_state(gen[3120])
		); 

/******************* CELL 3121 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3121 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3025]),
			.N(gen[3026]),
			.NE(gen[3027]),

			.O(gen[3120]),
			.E(gen[3122]),

			.SO(gen[3215]),
			.S(gen[3216]),
			.SE(gen[3217]),

			.SELF(gen[3121]),
			.cell_state(gen[3121])
		); 

/******************* CELL 3122 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3122 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3026]),
			.N(gen[3027]),
			.NE(gen[3028]),

			.O(gen[3121]),
			.E(gen[3123]),

			.SO(gen[3216]),
			.S(gen[3217]),
			.SE(gen[3218]),

			.SELF(gen[3122]),
			.cell_state(gen[3122])
		); 

/******************* CELL 3123 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3123 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3027]),
			.N(gen[3028]),
			.NE(gen[3029]),

			.O(gen[3122]),
			.E(gen[3124]),

			.SO(gen[3217]),
			.S(gen[3218]),
			.SE(gen[3219]),

			.SELF(gen[3123]),
			.cell_state(gen[3123])
		); 

/******************* CELL 3124 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3124 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3028]),
			.N(gen[3029]),
			.NE(gen[3030]),

			.O(gen[3123]),
			.E(gen[3125]),

			.SO(gen[3218]),
			.S(gen[3219]),
			.SE(gen[3220]),

			.SELF(gen[3124]),
			.cell_state(gen[3124])
		); 

/******************* CELL 3125 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3125 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3029]),
			.N(gen[3030]),
			.NE(gen[3031]),

			.O(gen[3124]),
			.E(gen[3126]),

			.SO(gen[3219]),
			.S(gen[3220]),
			.SE(gen[3221]),

			.SELF(gen[3125]),
			.cell_state(gen[3125])
		); 

/******************* CELL 3126 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3126 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3030]),
			.N(gen[3031]),
			.NE(gen[3032]),

			.O(gen[3125]),
			.E(gen[3127]),

			.SO(gen[3220]),
			.S(gen[3221]),
			.SE(gen[3222]),

			.SELF(gen[3126]),
			.cell_state(gen[3126])
		); 

/******************* CELL 3127 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3127 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3031]),
			.N(gen[3032]),
			.NE(gen[3033]),

			.O(gen[3126]),
			.E(gen[3128]),

			.SO(gen[3221]),
			.S(gen[3222]),
			.SE(gen[3223]),

			.SELF(gen[3127]),
			.cell_state(gen[3127])
		); 

/******************* CELL 3128 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3128 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3032]),
			.N(gen[3033]),
			.NE(gen[3034]),

			.O(gen[3127]),
			.E(gen[3129]),

			.SO(gen[3222]),
			.S(gen[3223]),
			.SE(gen[3224]),

			.SELF(gen[3128]),
			.cell_state(gen[3128])
		); 

/******************* CELL 3129 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3129 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3033]),
			.N(gen[3034]),
			.NE(gen[3035]),

			.O(gen[3128]),
			.E(gen[3130]),

			.SO(gen[3223]),
			.S(gen[3224]),
			.SE(gen[3225]),

			.SELF(gen[3129]),
			.cell_state(gen[3129])
		); 

/******************* CELL 3130 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3130 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3034]),
			.N(gen[3035]),
			.NE(gen[3036]),

			.O(gen[3129]),
			.E(gen[3131]),

			.SO(gen[3224]),
			.S(gen[3225]),
			.SE(gen[3226]),

			.SELF(gen[3130]),
			.cell_state(gen[3130])
		); 

/******************* CELL 3131 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3131 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3035]),
			.N(gen[3036]),
			.NE(gen[3037]),

			.O(gen[3130]),
			.E(gen[3132]),

			.SO(gen[3225]),
			.S(gen[3226]),
			.SE(gen[3227]),

			.SELF(gen[3131]),
			.cell_state(gen[3131])
		); 

/******************* CELL 3132 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3132 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3036]),
			.N(gen[3037]),
			.NE(gen[3038]),

			.O(gen[3131]),
			.E(gen[3133]),

			.SO(gen[3226]),
			.S(gen[3227]),
			.SE(gen[3228]),

			.SELF(gen[3132]),
			.cell_state(gen[3132])
		); 

/******************* CELL 3133 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3133 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3037]),
			.N(gen[3038]),
			.NE(gen[3039]),

			.O(gen[3132]),
			.E(gen[3134]),

			.SO(gen[3227]),
			.S(gen[3228]),
			.SE(gen[3229]),

			.SELF(gen[3133]),
			.cell_state(gen[3133])
		); 

/******************* CELL 3134 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3134 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3038]),
			.N(gen[3039]),
			.NE(gen[3038]),

			.O(gen[3133]),
			.E(gen[3133]),

			.SO(gen[3228]),
			.S(gen[3229]),
			.SE(gen[3228]),

			.SELF(gen[3134]),
			.cell_state(gen[3134])
		); 

/******************* CELL 3135 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3135 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3041]),
			.N(gen[3040]),
			.NE(gen[3041]),

			.O(gen[3136]),
			.E(gen[3136]),

			.SO(gen[3231]),
			.S(gen[3230]),
			.SE(gen[3231]),

			.SELF(gen[3135]),
			.cell_state(gen[3135])
		); 

/******************* CELL 3136 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3136 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3040]),
			.N(gen[3041]),
			.NE(gen[3042]),

			.O(gen[3135]),
			.E(gen[3137]),

			.SO(gen[3230]),
			.S(gen[3231]),
			.SE(gen[3232]),

			.SELF(gen[3136]),
			.cell_state(gen[3136])
		); 

/******************* CELL 3137 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3137 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3041]),
			.N(gen[3042]),
			.NE(gen[3043]),

			.O(gen[3136]),
			.E(gen[3138]),

			.SO(gen[3231]),
			.S(gen[3232]),
			.SE(gen[3233]),

			.SELF(gen[3137]),
			.cell_state(gen[3137])
		); 

/******************* CELL 3138 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3138 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3042]),
			.N(gen[3043]),
			.NE(gen[3044]),

			.O(gen[3137]),
			.E(gen[3139]),

			.SO(gen[3232]),
			.S(gen[3233]),
			.SE(gen[3234]),

			.SELF(gen[3138]),
			.cell_state(gen[3138])
		); 

/******************* CELL 3139 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3139 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3043]),
			.N(gen[3044]),
			.NE(gen[3045]),

			.O(gen[3138]),
			.E(gen[3140]),

			.SO(gen[3233]),
			.S(gen[3234]),
			.SE(gen[3235]),

			.SELF(gen[3139]),
			.cell_state(gen[3139])
		); 

/******************* CELL 3140 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3140 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3044]),
			.N(gen[3045]),
			.NE(gen[3046]),

			.O(gen[3139]),
			.E(gen[3141]),

			.SO(gen[3234]),
			.S(gen[3235]),
			.SE(gen[3236]),

			.SELF(gen[3140]),
			.cell_state(gen[3140])
		); 

/******************* CELL 3141 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3141 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3045]),
			.N(gen[3046]),
			.NE(gen[3047]),

			.O(gen[3140]),
			.E(gen[3142]),

			.SO(gen[3235]),
			.S(gen[3236]),
			.SE(gen[3237]),

			.SELF(gen[3141]),
			.cell_state(gen[3141])
		); 

/******************* CELL 3142 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3142 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3046]),
			.N(gen[3047]),
			.NE(gen[3048]),

			.O(gen[3141]),
			.E(gen[3143]),

			.SO(gen[3236]),
			.S(gen[3237]),
			.SE(gen[3238]),

			.SELF(gen[3142]),
			.cell_state(gen[3142])
		); 

/******************* CELL 3143 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3143 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3047]),
			.N(gen[3048]),
			.NE(gen[3049]),

			.O(gen[3142]),
			.E(gen[3144]),

			.SO(gen[3237]),
			.S(gen[3238]),
			.SE(gen[3239]),

			.SELF(gen[3143]),
			.cell_state(gen[3143])
		); 

/******************* CELL 3144 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3144 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3048]),
			.N(gen[3049]),
			.NE(gen[3050]),

			.O(gen[3143]),
			.E(gen[3145]),

			.SO(gen[3238]),
			.S(gen[3239]),
			.SE(gen[3240]),

			.SELF(gen[3144]),
			.cell_state(gen[3144])
		); 

/******************* CELL 3145 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3145 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3049]),
			.N(gen[3050]),
			.NE(gen[3051]),

			.O(gen[3144]),
			.E(gen[3146]),

			.SO(gen[3239]),
			.S(gen[3240]),
			.SE(gen[3241]),

			.SELF(gen[3145]),
			.cell_state(gen[3145])
		); 

/******************* CELL 3146 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3146 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3050]),
			.N(gen[3051]),
			.NE(gen[3052]),

			.O(gen[3145]),
			.E(gen[3147]),

			.SO(gen[3240]),
			.S(gen[3241]),
			.SE(gen[3242]),

			.SELF(gen[3146]),
			.cell_state(gen[3146])
		); 

/******************* CELL 3147 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3147 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3051]),
			.N(gen[3052]),
			.NE(gen[3053]),

			.O(gen[3146]),
			.E(gen[3148]),

			.SO(gen[3241]),
			.S(gen[3242]),
			.SE(gen[3243]),

			.SELF(gen[3147]),
			.cell_state(gen[3147])
		); 

/******************* CELL 3148 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3148 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3052]),
			.N(gen[3053]),
			.NE(gen[3054]),

			.O(gen[3147]),
			.E(gen[3149]),

			.SO(gen[3242]),
			.S(gen[3243]),
			.SE(gen[3244]),

			.SELF(gen[3148]),
			.cell_state(gen[3148])
		); 

/******************* CELL 3149 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3149 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3053]),
			.N(gen[3054]),
			.NE(gen[3055]),

			.O(gen[3148]),
			.E(gen[3150]),

			.SO(gen[3243]),
			.S(gen[3244]),
			.SE(gen[3245]),

			.SELF(gen[3149]),
			.cell_state(gen[3149])
		); 

/******************* CELL 3150 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3150 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3054]),
			.N(gen[3055]),
			.NE(gen[3056]),

			.O(gen[3149]),
			.E(gen[3151]),

			.SO(gen[3244]),
			.S(gen[3245]),
			.SE(gen[3246]),

			.SELF(gen[3150]),
			.cell_state(gen[3150])
		); 

/******************* CELL 3151 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3151 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3055]),
			.N(gen[3056]),
			.NE(gen[3057]),

			.O(gen[3150]),
			.E(gen[3152]),

			.SO(gen[3245]),
			.S(gen[3246]),
			.SE(gen[3247]),

			.SELF(gen[3151]),
			.cell_state(gen[3151])
		); 

/******************* CELL 3152 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3152 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3056]),
			.N(gen[3057]),
			.NE(gen[3058]),

			.O(gen[3151]),
			.E(gen[3153]),

			.SO(gen[3246]),
			.S(gen[3247]),
			.SE(gen[3248]),

			.SELF(gen[3152]),
			.cell_state(gen[3152])
		); 

/******************* CELL 3153 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3153 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3057]),
			.N(gen[3058]),
			.NE(gen[3059]),

			.O(gen[3152]),
			.E(gen[3154]),

			.SO(gen[3247]),
			.S(gen[3248]),
			.SE(gen[3249]),

			.SELF(gen[3153]),
			.cell_state(gen[3153])
		); 

/******************* CELL 3154 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3154 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3058]),
			.N(gen[3059]),
			.NE(gen[3060]),

			.O(gen[3153]),
			.E(gen[3155]),

			.SO(gen[3248]),
			.S(gen[3249]),
			.SE(gen[3250]),

			.SELF(gen[3154]),
			.cell_state(gen[3154])
		); 

/******************* CELL 3155 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3155 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3059]),
			.N(gen[3060]),
			.NE(gen[3061]),

			.O(gen[3154]),
			.E(gen[3156]),

			.SO(gen[3249]),
			.S(gen[3250]),
			.SE(gen[3251]),

			.SELF(gen[3155]),
			.cell_state(gen[3155])
		); 

/******************* CELL 3156 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3156 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3060]),
			.N(gen[3061]),
			.NE(gen[3062]),

			.O(gen[3155]),
			.E(gen[3157]),

			.SO(gen[3250]),
			.S(gen[3251]),
			.SE(gen[3252]),

			.SELF(gen[3156]),
			.cell_state(gen[3156])
		); 

/******************* CELL 3157 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3157 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3061]),
			.N(gen[3062]),
			.NE(gen[3063]),

			.O(gen[3156]),
			.E(gen[3158]),

			.SO(gen[3251]),
			.S(gen[3252]),
			.SE(gen[3253]),

			.SELF(gen[3157]),
			.cell_state(gen[3157])
		); 

/******************* CELL 3158 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3158 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3062]),
			.N(gen[3063]),
			.NE(gen[3064]),

			.O(gen[3157]),
			.E(gen[3159]),

			.SO(gen[3252]),
			.S(gen[3253]),
			.SE(gen[3254]),

			.SELF(gen[3158]),
			.cell_state(gen[3158])
		); 

/******************* CELL 3159 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3159 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3063]),
			.N(gen[3064]),
			.NE(gen[3065]),

			.O(gen[3158]),
			.E(gen[3160]),

			.SO(gen[3253]),
			.S(gen[3254]),
			.SE(gen[3255]),

			.SELF(gen[3159]),
			.cell_state(gen[3159])
		); 

/******************* CELL 3160 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3160 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3064]),
			.N(gen[3065]),
			.NE(gen[3066]),

			.O(gen[3159]),
			.E(gen[3161]),

			.SO(gen[3254]),
			.S(gen[3255]),
			.SE(gen[3256]),

			.SELF(gen[3160]),
			.cell_state(gen[3160])
		); 

/******************* CELL 3161 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3161 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3065]),
			.N(gen[3066]),
			.NE(gen[3067]),

			.O(gen[3160]),
			.E(gen[3162]),

			.SO(gen[3255]),
			.S(gen[3256]),
			.SE(gen[3257]),

			.SELF(gen[3161]),
			.cell_state(gen[3161])
		); 

/******************* CELL 3162 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3162 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3066]),
			.N(gen[3067]),
			.NE(gen[3068]),

			.O(gen[3161]),
			.E(gen[3163]),

			.SO(gen[3256]),
			.S(gen[3257]),
			.SE(gen[3258]),

			.SELF(gen[3162]),
			.cell_state(gen[3162])
		); 

/******************* CELL 3163 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3163 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3067]),
			.N(gen[3068]),
			.NE(gen[3069]),

			.O(gen[3162]),
			.E(gen[3164]),

			.SO(gen[3257]),
			.S(gen[3258]),
			.SE(gen[3259]),

			.SELF(gen[3163]),
			.cell_state(gen[3163])
		); 

/******************* CELL 3164 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3164 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3068]),
			.N(gen[3069]),
			.NE(gen[3070]),

			.O(gen[3163]),
			.E(gen[3165]),

			.SO(gen[3258]),
			.S(gen[3259]),
			.SE(gen[3260]),

			.SELF(gen[3164]),
			.cell_state(gen[3164])
		); 

/******************* CELL 3165 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3165 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3069]),
			.N(gen[3070]),
			.NE(gen[3071]),

			.O(gen[3164]),
			.E(gen[3166]),

			.SO(gen[3259]),
			.S(gen[3260]),
			.SE(gen[3261]),

			.SELF(gen[3165]),
			.cell_state(gen[3165])
		); 

/******************* CELL 3166 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3166 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3070]),
			.N(gen[3071]),
			.NE(gen[3072]),

			.O(gen[3165]),
			.E(gen[3167]),

			.SO(gen[3260]),
			.S(gen[3261]),
			.SE(gen[3262]),

			.SELF(gen[3166]),
			.cell_state(gen[3166])
		); 

/******************* CELL 3167 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3167 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3071]),
			.N(gen[3072]),
			.NE(gen[3073]),

			.O(gen[3166]),
			.E(gen[3168]),

			.SO(gen[3261]),
			.S(gen[3262]),
			.SE(gen[3263]),

			.SELF(gen[3167]),
			.cell_state(gen[3167])
		); 

/******************* CELL 3168 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3168 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3072]),
			.N(gen[3073]),
			.NE(gen[3074]),

			.O(gen[3167]),
			.E(gen[3169]),

			.SO(gen[3262]),
			.S(gen[3263]),
			.SE(gen[3264]),

			.SELF(gen[3168]),
			.cell_state(gen[3168])
		); 

/******************* CELL 3169 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3169 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3073]),
			.N(gen[3074]),
			.NE(gen[3075]),

			.O(gen[3168]),
			.E(gen[3170]),

			.SO(gen[3263]),
			.S(gen[3264]),
			.SE(gen[3265]),

			.SELF(gen[3169]),
			.cell_state(gen[3169])
		); 

/******************* CELL 3170 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3170 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3074]),
			.N(gen[3075]),
			.NE(gen[3076]),

			.O(gen[3169]),
			.E(gen[3171]),

			.SO(gen[3264]),
			.S(gen[3265]),
			.SE(gen[3266]),

			.SELF(gen[3170]),
			.cell_state(gen[3170])
		); 

/******************* CELL 3171 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3171 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3075]),
			.N(gen[3076]),
			.NE(gen[3077]),

			.O(gen[3170]),
			.E(gen[3172]),

			.SO(gen[3265]),
			.S(gen[3266]),
			.SE(gen[3267]),

			.SELF(gen[3171]),
			.cell_state(gen[3171])
		); 

/******************* CELL 3172 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3172 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3076]),
			.N(gen[3077]),
			.NE(gen[3078]),

			.O(gen[3171]),
			.E(gen[3173]),

			.SO(gen[3266]),
			.S(gen[3267]),
			.SE(gen[3268]),

			.SELF(gen[3172]),
			.cell_state(gen[3172])
		); 

/******************* CELL 3173 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3173 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3077]),
			.N(gen[3078]),
			.NE(gen[3079]),

			.O(gen[3172]),
			.E(gen[3174]),

			.SO(gen[3267]),
			.S(gen[3268]),
			.SE(gen[3269]),

			.SELF(gen[3173]),
			.cell_state(gen[3173])
		); 

/******************* CELL 3174 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3174 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3078]),
			.N(gen[3079]),
			.NE(gen[3080]),

			.O(gen[3173]),
			.E(gen[3175]),

			.SO(gen[3268]),
			.S(gen[3269]),
			.SE(gen[3270]),

			.SELF(gen[3174]),
			.cell_state(gen[3174])
		); 

/******************* CELL 3175 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3175 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3079]),
			.N(gen[3080]),
			.NE(gen[3081]),

			.O(gen[3174]),
			.E(gen[3176]),

			.SO(gen[3269]),
			.S(gen[3270]),
			.SE(gen[3271]),

			.SELF(gen[3175]),
			.cell_state(gen[3175])
		); 

/******************* CELL 3176 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3176 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3080]),
			.N(gen[3081]),
			.NE(gen[3082]),

			.O(gen[3175]),
			.E(gen[3177]),

			.SO(gen[3270]),
			.S(gen[3271]),
			.SE(gen[3272]),

			.SELF(gen[3176]),
			.cell_state(gen[3176])
		); 

/******************* CELL 3177 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3177 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3081]),
			.N(gen[3082]),
			.NE(gen[3083]),

			.O(gen[3176]),
			.E(gen[3178]),

			.SO(gen[3271]),
			.S(gen[3272]),
			.SE(gen[3273]),

			.SELF(gen[3177]),
			.cell_state(gen[3177])
		); 

/******************* CELL 3178 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3178 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3082]),
			.N(gen[3083]),
			.NE(gen[3084]),

			.O(gen[3177]),
			.E(gen[3179]),

			.SO(gen[3272]),
			.S(gen[3273]),
			.SE(gen[3274]),

			.SELF(gen[3178]),
			.cell_state(gen[3178])
		); 

/******************* CELL 3179 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3179 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3083]),
			.N(gen[3084]),
			.NE(gen[3085]),

			.O(gen[3178]),
			.E(gen[3180]),

			.SO(gen[3273]),
			.S(gen[3274]),
			.SE(gen[3275]),

			.SELF(gen[3179]),
			.cell_state(gen[3179])
		); 

/******************* CELL 3180 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3180 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3084]),
			.N(gen[3085]),
			.NE(gen[3086]),

			.O(gen[3179]),
			.E(gen[3181]),

			.SO(gen[3274]),
			.S(gen[3275]),
			.SE(gen[3276]),

			.SELF(gen[3180]),
			.cell_state(gen[3180])
		); 

/******************* CELL 3181 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3181 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3085]),
			.N(gen[3086]),
			.NE(gen[3087]),

			.O(gen[3180]),
			.E(gen[3182]),

			.SO(gen[3275]),
			.S(gen[3276]),
			.SE(gen[3277]),

			.SELF(gen[3181]),
			.cell_state(gen[3181])
		); 

/******************* CELL 3182 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3182 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3086]),
			.N(gen[3087]),
			.NE(gen[3088]),

			.O(gen[3181]),
			.E(gen[3183]),

			.SO(gen[3276]),
			.S(gen[3277]),
			.SE(gen[3278]),

			.SELF(gen[3182]),
			.cell_state(gen[3182])
		); 

/******************* CELL 3183 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3183 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3087]),
			.N(gen[3088]),
			.NE(gen[3089]),

			.O(gen[3182]),
			.E(gen[3184]),

			.SO(gen[3277]),
			.S(gen[3278]),
			.SE(gen[3279]),

			.SELF(gen[3183]),
			.cell_state(gen[3183])
		); 

/******************* CELL 3184 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3184 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3088]),
			.N(gen[3089]),
			.NE(gen[3090]),

			.O(gen[3183]),
			.E(gen[3185]),

			.SO(gen[3278]),
			.S(gen[3279]),
			.SE(gen[3280]),

			.SELF(gen[3184]),
			.cell_state(gen[3184])
		); 

/******************* CELL 3185 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3185 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3089]),
			.N(gen[3090]),
			.NE(gen[3091]),

			.O(gen[3184]),
			.E(gen[3186]),

			.SO(gen[3279]),
			.S(gen[3280]),
			.SE(gen[3281]),

			.SELF(gen[3185]),
			.cell_state(gen[3185])
		); 

/******************* CELL 3186 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3186 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3090]),
			.N(gen[3091]),
			.NE(gen[3092]),

			.O(gen[3185]),
			.E(gen[3187]),

			.SO(gen[3280]),
			.S(gen[3281]),
			.SE(gen[3282]),

			.SELF(gen[3186]),
			.cell_state(gen[3186])
		); 

/******************* CELL 3187 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3187 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3091]),
			.N(gen[3092]),
			.NE(gen[3093]),

			.O(gen[3186]),
			.E(gen[3188]),

			.SO(gen[3281]),
			.S(gen[3282]),
			.SE(gen[3283]),

			.SELF(gen[3187]),
			.cell_state(gen[3187])
		); 

/******************* CELL 3188 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3188 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3092]),
			.N(gen[3093]),
			.NE(gen[3094]),

			.O(gen[3187]),
			.E(gen[3189]),

			.SO(gen[3282]),
			.S(gen[3283]),
			.SE(gen[3284]),

			.SELF(gen[3188]),
			.cell_state(gen[3188])
		); 

/******************* CELL 3189 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3189 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3093]),
			.N(gen[3094]),
			.NE(gen[3095]),

			.O(gen[3188]),
			.E(gen[3190]),

			.SO(gen[3283]),
			.S(gen[3284]),
			.SE(gen[3285]),

			.SELF(gen[3189]),
			.cell_state(gen[3189])
		); 

/******************* CELL 3190 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3190 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3094]),
			.N(gen[3095]),
			.NE(gen[3096]),

			.O(gen[3189]),
			.E(gen[3191]),

			.SO(gen[3284]),
			.S(gen[3285]),
			.SE(gen[3286]),

			.SELF(gen[3190]),
			.cell_state(gen[3190])
		); 

/******************* CELL 3191 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3191 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3095]),
			.N(gen[3096]),
			.NE(gen[3097]),

			.O(gen[3190]),
			.E(gen[3192]),

			.SO(gen[3285]),
			.S(gen[3286]),
			.SE(gen[3287]),

			.SELF(gen[3191]),
			.cell_state(gen[3191])
		); 

/******************* CELL 3192 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3192 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3096]),
			.N(gen[3097]),
			.NE(gen[3098]),

			.O(gen[3191]),
			.E(gen[3193]),

			.SO(gen[3286]),
			.S(gen[3287]),
			.SE(gen[3288]),

			.SELF(gen[3192]),
			.cell_state(gen[3192])
		); 

/******************* CELL 3193 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3193 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3097]),
			.N(gen[3098]),
			.NE(gen[3099]),

			.O(gen[3192]),
			.E(gen[3194]),

			.SO(gen[3287]),
			.S(gen[3288]),
			.SE(gen[3289]),

			.SELF(gen[3193]),
			.cell_state(gen[3193])
		); 

/******************* CELL 3194 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3194 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3098]),
			.N(gen[3099]),
			.NE(gen[3100]),

			.O(gen[3193]),
			.E(gen[3195]),

			.SO(gen[3288]),
			.S(gen[3289]),
			.SE(gen[3290]),

			.SELF(gen[3194]),
			.cell_state(gen[3194])
		); 

/******************* CELL 3195 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3195 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3099]),
			.N(gen[3100]),
			.NE(gen[3101]),

			.O(gen[3194]),
			.E(gen[3196]),

			.SO(gen[3289]),
			.S(gen[3290]),
			.SE(gen[3291]),

			.SELF(gen[3195]),
			.cell_state(gen[3195])
		); 

/******************* CELL 3196 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3196 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3100]),
			.N(gen[3101]),
			.NE(gen[3102]),

			.O(gen[3195]),
			.E(gen[3197]),

			.SO(gen[3290]),
			.S(gen[3291]),
			.SE(gen[3292]),

			.SELF(gen[3196]),
			.cell_state(gen[3196])
		); 

/******************* CELL 3197 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3197 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3101]),
			.N(gen[3102]),
			.NE(gen[3103]),

			.O(gen[3196]),
			.E(gen[3198]),

			.SO(gen[3291]),
			.S(gen[3292]),
			.SE(gen[3293]),

			.SELF(gen[3197]),
			.cell_state(gen[3197])
		); 

/******************* CELL 3198 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3198 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3102]),
			.N(gen[3103]),
			.NE(gen[3104]),

			.O(gen[3197]),
			.E(gen[3199]),

			.SO(gen[3292]),
			.S(gen[3293]),
			.SE(gen[3294]),

			.SELF(gen[3198]),
			.cell_state(gen[3198])
		); 

/******************* CELL 3199 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3199 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3103]),
			.N(gen[3104]),
			.NE(gen[3105]),

			.O(gen[3198]),
			.E(gen[3200]),

			.SO(gen[3293]),
			.S(gen[3294]),
			.SE(gen[3295]),

			.SELF(gen[3199]),
			.cell_state(gen[3199])
		); 

/******************* CELL 3200 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3200 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3104]),
			.N(gen[3105]),
			.NE(gen[3106]),

			.O(gen[3199]),
			.E(gen[3201]),

			.SO(gen[3294]),
			.S(gen[3295]),
			.SE(gen[3296]),

			.SELF(gen[3200]),
			.cell_state(gen[3200])
		); 

/******************* CELL 3201 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3201 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3105]),
			.N(gen[3106]),
			.NE(gen[3107]),

			.O(gen[3200]),
			.E(gen[3202]),

			.SO(gen[3295]),
			.S(gen[3296]),
			.SE(gen[3297]),

			.SELF(gen[3201]),
			.cell_state(gen[3201])
		); 

/******************* CELL 3202 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3202 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3106]),
			.N(gen[3107]),
			.NE(gen[3108]),

			.O(gen[3201]),
			.E(gen[3203]),

			.SO(gen[3296]),
			.S(gen[3297]),
			.SE(gen[3298]),

			.SELF(gen[3202]),
			.cell_state(gen[3202])
		); 

/******************* CELL 3203 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3203 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3107]),
			.N(gen[3108]),
			.NE(gen[3109]),

			.O(gen[3202]),
			.E(gen[3204]),

			.SO(gen[3297]),
			.S(gen[3298]),
			.SE(gen[3299]),

			.SELF(gen[3203]),
			.cell_state(gen[3203])
		); 

/******************* CELL 3204 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3204 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3108]),
			.N(gen[3109]),
			.NE(gen[3110]),

			.O(gen[3203]),
			.E(gen[3205]),

			.SO(gen[3298]),
			.S(gen[3299]),
			.SE(gen[3300]),

			.SELF(gen[3204]),
			.cell_state(gen[3204])
		); 

/******************* CELL 3205 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3205 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3109]),
			.N(gen[3110]),
			.NE(gen[3111]),

			.O(gen[3204]),
			.E(gen[3206]),

			.SO(gen[3299]),
			.S(gen[3300]),
			.SE(gen[3301]),

			.SELF(gen[3205]),
			.cell_state(gen[3205])
		); 

/******************* CELL 3206 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3206 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3110]),
			.N(gen[3111]),
			.NE(gen[3112]),

			.O(gen[3205]),
			.E(gen[3207]),

			.SO(gen[3300]),
			.S(gen[3301]),
			.SE(gen[3302]),

			.SELF(gen[3206]),
			.cell_state(gen[3206])
		); 

/******************* CELL 3207 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3207 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3111]),
			.N(gen[3112]),
			.NE(gen[3113]),

			.O(gen[3206]),
			.E(gen[3208]),

			.SO(gen[3301]),
			.S(gen[3302]),
			.SE(gen[3303]),

			.SELF(gen[3207]),
			.cell_state(gen[3207])
		); 

/******************* CELL 3208 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3208 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3112]),
			.N(gen[3113]),
			.NE(gen[3114]),

			.O(gen[3207]),
			.E(gen[3209]),

			.SO(gen[3302]),
			.S(gen[3303]),
			.SE(gen[3304]),

			.SELF(gen[3208]),
			.cell_state(gen[3208])
		); 

/******************* CELL 3209 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3209 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3113]),
			.N(gen[3114]),
			.NE(gen[3115]),

			.O(gen[3208]),
			.E(gen[3210]),

			.SO(gen[3303]),
			.S(gen[3304]),
			.SE(gen[3305]),

			.SELF(gen[3209]),
			.cell_state(gen[3209])
		); 

/******************* CELL 3210 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3210 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3114]),
			.N(gen[3115]),
			.NE(gen[3116]),

			.O(gen[3209]),
			.E(gen[3211]),

			.SO(gen[3304]),
			.S(gen[3305]),
			.SE(gen[3306]),

			.SELF(gen[3210]),
			.cell_state(gen[3210])
		); 

/******************* CELL 3211 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3211 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3115]),
			.N(gen[3116]),
			.NE(gen[3117]),

			.O(gen[3210]),
			.E(gen[3212]),

			.SO(gen[3305]),
			.S(gen[3306]),
			.SE(gen[3307]),

			.SELF(gen[3211]),
			.cell_state(gen[3211])
		); 

/******************* CELL 3212 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3212 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3116]),
			.N(gen[3117]),
			.NE(gen[3118]),

			.O(gen[3211]),
			.E(gen[3213]),

			.SO(gen[3306]),
			.S(gen[3307]),
			.SE(gen[3308]),

			.SELF(gen[3212]),
			.cell_state(gen[3212])
		); 

/******************* CELL 3213 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3213 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3117]),
			.N(gen[3118]),
			.NE(gen[3119]),

			.O(gen[3212]),
			.E(gen[3214]),

			.SO(gen[3307]),
			.S(gen[3308]),
			.SE(gen[3309]),

			.SELF(gen[3213]),
			.cell_state(gen[3213])
		); 

/******************* CELL 3214 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3214 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3118]),
			.N(gen[3119]),
			.NE(gen[3120]),

			.O(gen[3213]),
			.E(gen[3215]),

			.SO(gen[3308]),
			.S(gen[3309]),
			.SE(gen[3310]),

			.SELF(gen[3214]),
			.cell_state(gen[3214])
		); 

/******************* CELL 3215 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3215 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3119]),
			.N(gen[3120]),
			.NE(gen[3121]),

			.O(gen[3214]),
			.E(gen[3216]),

			.SO(gen[3309]),
			.S(gen[3310]),
			.SE(gen[3311]),

			.SELF(gen[3215]),
			.cell_state(gen[3215])
		); 

/******************* CELL 3216 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3216 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3120]),
			.N(gen[3121]),
			.NE(gen[3122]),

			.O(gen[3215]),
			.E(gen[3217]),

			.SO(gen[3310]),
			.S(gen[3311]),
			.SE(gen[3312]),

			.SELF(gen[3216]),
			.cell_state(gen[3216])
		); 

/******************* CELL 3217 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3217 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3121]),
			.N(gen[3122]),
			.NE(gen[3123]),

			.O(gen[3216]),
			.E(gen[3218]),

			.SO(gen[3311]),
			.S(gen[3312]),
			.SE(gen[3313]),

			.SELF(gen[3217]),
			.cell_state(gen[3217])
		); 

/******************* CELL 3218 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3218 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3122]),
			.N(gen[3123]),
			.NE(gen[3124]),

			.O(gen[3217]),
			.E(gen[3219]),

			.SO(gen[3312]),
			.S(gen[3313]),
			.SE(gen[3314]),

			.SELF(gen[3218]),
			.cell_state(gen[3218])
		); 

/******************* CELL 3219 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3219 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3123]),
			.N(gen[3124]),
			.NE(gen[3125]),

			.O(gen[3218]),
			.E(gen[3220]),

			.SO(gen[3313]),
			.S(gen[3314]),
			.SE(gen[3315]),

			.SELF(gen[3219]),
			.cell_state(gen[3219])
		); 

/******************* CELL 3220 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3220 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3124]),
			.N(gen[3125]),
			.NE(gen[3126]),

			.O(gen[3219]),
			.E(gen[3221]),

			.SO(gen[3314]),
			.S(gen[3315]),
			.SE(gen[3316]),

			.SELF(gen[3220]),
			.cell_state(gen[3220])
		); 

/******************* CELL 3221 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3221 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3125]),
			.N(gen[3126]),
			.NE(gen[3127]),

			.O(gen[3220]),
			.E(gen[3222]),

			.SO(gen[3315]),
			.S(gen[3316]),
			.SE(gen[3317]),

			.SELF(gen[3221]),
			.cell_state(gen[3221])
		); 

/******************* CELL 3222 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3222 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3126]),
			.N(gen[3127]),
			.NE(gen[3128]),

			.O(gen[3221]),
			.E(gen[3223]),

			.SO(gen[3316]),
			.S(gen[3317]),
			.SE(gen[3318]),

			.SELF(gen[3222]),
			.cell_state(gen[3222])
		); 

/******************* CELL 3223 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3223 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3127]),
			.N(gen[3128]),
			.NE(gen[3129]),

			.O(gen[3222]),
			.E(gen[3224]),

			.SO(gen[3317]),
			.S(gen[3318]),
			.SE(gen[3319]),

			.SELF(gen[3223]),
			.cell_state(gen[3223])
		); 

/******************* CELL 3224 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3224 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3128]),
			.N(gen[3129]),
			.NE(gen[3130]),

			.O(gen[3223]),
			.E(gen[3225]),

			.SO(gen[3318]),
			.S(gen[3319]),
			.SE(gen[3320]),

			.SELF(gen[3224]),
			.cell_state(gen[3224])
		); 

/******************* CELL 3225 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3225 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3129]),
			.N(gen[3130]),
			.NE(gen[3131]),

			.O(gen[3224]),
			.E(gen[3226]),

			.SO(gen[3319]),
			.S(gen[3320]),
			.SE(gen[3321]),

			.SELF(gen[3225]),
			.cell_state(gen[3225])
		); 

/******************* CELL 3226 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3226 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3130]),
			.N(gen[3131]),
			.NE(gen[3132]),

			.O(gen[3225]),
			.E(gen[3227]),

			.SO(gen[3320]),
			.S(gen[3321]),
			.SE(gen[3322]),

			.SELF(gen[3226]),
			.cell_state(gen[3226])
		); 

/******************* CELL 3227 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3227 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3131]),
			.N(gen[3132]),
			.NE(gen[3133]),

			.O(gen[3226]),
			.E(gen[3228]),

			.SO(gen[3321]),
			.S(gen[3322]),
			.SE(gen[3323]),

			.SELF(gen[3227]),
			.cell_state(gen[3227])
		); 

/******************* CELL 3228 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3228 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3132]),
			.N(gen[3133]),
			.NE(gen[3134]),

			.O(gen[3227]),
			.E(gen[3229]),

			.SO(gen[3322]),
			.S(gen[3323]),
			.SE(gen[3324]),

			.SELF(gen[3228]),
			.cell_state(gen[3228])
		); 

/******************* CELL 3229 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3229 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3133]),
			.N(gen[3134]),
			.NE(gen[3133]),

			.O(gen[3228]),
			.E(gen[3228]),

			.SO(gen[3323]),
			.S(gen[3324]),
			.SE(gen[3323]),

			.SELF(gen[3229]),
			.cell_state(gen[3229])
		); 

/******************* CELL 3230 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3230 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3136]),
			.N(gen[3135]),
			.NE(gen[3136]),

			.O(gen[3231]),
			.E(gen[3231]),

			.SO(gen[3326]),
			.S(gen[3325]),
			.SE(gen[3326]),

			.SELF(gen[3230]),
			.cell_state(gen[3230])
		); 

/******************* CELL 3231 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3231 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3135]),
			.N(gen[3136]),
			.NE(gen[3137]),

			.O(gen[3230]),
			.E(gen[3232]),

			.SO(gen[3325]),
			.S(gen[3326]),
			.SE(gen[3327]),

			.SELF(gen[3231]),
			.cell_state(gen[3231])
		); 

/******************* CELL 3232 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3232 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3136]),
			.N(gen[3137]),
			.NE(gen[3138]),

			.O(gen[3231]),
			.E(gen[3233]),

			.SO(gen[3326]),
			.S(gen[3327]),
			.SE(gen[3328]),

			.SELF(gen[3232]),
			.cell_state(gen[3232])
		); 

/******************* CELL 3233 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3233 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3137]),
			.N(gen[3138]),
			.NE(gen[3139]),

			.O(gen[3232]),
			.E(gen[3234]),

			.SO(gen[3327]),
			.S(gen[3328]),
			.SE(gen[3329]),

			.SELF(gen[3233]),
			.cell_state(gen[3233])
		); 

/******************* CELL 3234 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3234 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3138]),
			.N(gen[3139]),
			.NE(gen[3140]),

			.O(gen[3233]),
			.E(gen[3235]),

			.SO(gen[3328]),
			.S(gen[3329]),
			.SE(gen[3330]),

			.SELF(gen[3234]),
			.cell_state(gen[3234])
		); 

/******************* CELL 3235 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3235 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3139]),
			.N(gen[3140]),
			.NE(gen[3141]),

			.O(gen[3234]),
			.E(gen[3236]),

			.SO(gen[3329]),
			.S(gen[3330]),
			.SE(gen[3331]),

			.SELF(gen[3235]),
			.cell_state(gen[3235])
		); 

/******************* CELL 3236 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3236 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3140]),
			.N(gen[3141]),
			.NE(gen[3142]),

			.O(gen[3235]),
			.E(gen[3237]),

			.SO(gen[3330]),
			.S(gen[3331]),
			.SE(gen[3332]),

			.SELF(gen[3236]),
			.cell_state(gen[3236])
		); 

/******************* CELL 3237 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3237 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3141]),
			.N(gen[3142]),
			.NE(gen[3143]),

			.O(gen[3236]),
			.E(gen[3238]),

			.SO(gen[3331]),
			.S(gen[3332]),
			.SE(gen[3333]),

			.SELF(gen[3237]),
			.cell_state(gen[3237])
		); 

/******************* CELL 3238 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3238 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3142]),
			.N(gen[3143]),
			.NE(gen[3144]),

			.O(gen[3237]),
			.E(gen[3239]),

			.SO(gen[3332]),
			.S(gen[3333]),
			.SE(gen[3334]),

			.SELF(gen[3238]),
			.cell_state(gen[3238])
		); 

/******************* CELL 3239 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3239 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3143]),
			.N(gen[3144]),
			.NE(gen[3145]),

			.O(gen[3238]),
			.E(gen[3240]),

			.SO(gen[3333]),
			.S(gen[3334]),
			.SE(gen[3335]),

			.SELF(gen[3239]),
			.cell_state(gen[3239])
		); 

/******************* CELL 3240 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3240 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3144]),
			.N(gen[3145]),
			.NE(gen[3146]),

			.O(gen[3239]),
			.E(gen[3241]),

			.SO(gen[3334]),
			.S(gen[3335]),
			.SE(gen[3336]),

			.SELF(gen[3240]),
			.cell_state(gen[3240])
		); 

/******************* CELL 3241 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3241 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3145]),
			.N(gen[3146]),
			.NE(gen[3147]),

			.O(gen[3240]),
			.E(gen[3242]),

			.SO(gen[3335]),
			.S(gen[3336]),
			.SE(gen[3337]),

			.SELF(gen[3241]),
			.cell_state(gen[3241])
		); 

/******************* CELL 3242 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3242 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3146]),
			.N(gen[3147]),
			.NE(gen[3148]),

			.O(gen[3241]),
			.E(gen[3243]),

			.SO(gen[3336]),
			.S(gen[3337]),
			.SE(gen[3338]),

			.SELF(gen[3242]),
			.cell_state(gen[3242])
		); 

/******************* CELL 3243 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3243 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3147]),
			.N(gen[3148]),
			.NE(gen[3149]),

			.O(gen[3242]),
			.E(gen[3244]),

			.SO(gen[3337]),
			.S(gen[3338]),
			.SE(gen[3339]),

			.SELF(gen[3243]),
			.cell_state(gen[3243])
		); 

/******************* CELL 3244 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3244 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3148]),
			.N(gen[3149]),
			.NE(gen[3150]),

			.O(gen[3243]),
			.E(gen[3245]),

			.SO(gen[3338]),
			.S(gen[3339]),
			.SE(gen[3340]),

			.SELF(gen[3244]),
			.cell_state(gen[3244])
		); 

/******************* CELL 3245 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3245 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3149]),
			.N(gen[3150]),
			.NE(gen[3151]),

			.O(gen[3244]),
			.E(gen[3246]),

			.SO(gen[3339]),
			.S(gen[3340]),
			.SE(gen[3341]),

			.SELF(gen[3245]),
			.cell_state(gen[3245])
		); 

/******************* CELL 3246 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3246 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3150]),
			.N(gen[3151]),
			.NE(gen[3152]),

			.O(gen[3245]),
			.E(gen[3247]),

			.SO(gen[3340]),
			.S(gen[3341]),
			.SE(gen[3342]),

			.SELF(gen[3246]),
			.cell_state(gen[3246])
		); 

/******************* CELL 3247 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3247 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3151]),
			.N(gen[3152]),
			.NE(gen[3153]),

			.O(gen[3246]),
			.E(gen[3248]),

			.SO(gen[3341]),
			.S(gen[3342]),
			.SE(gen[3343]),

			.SELF(gen[3247]),
			.cell_state(gen[3247])
		); 

/******************* CELL 3248 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3248 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3152]),
			.N(gen[3153]),
			.NE(gen[3154]),

			.O(gen[3247]),
			.E(gen[3249]),

			.SO(gen[3342]),
			.S(gen[3343]),
			.SE(gen[3344]),

			.SELF(gen[3248]),
			.cell_state(gen[3248])
		); 

/******************* CELL 3249 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3249 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3153]),
			.N(gen[3154]),
			.NE(gen[3155]),

			.O(gen[3248]),
			.E(gen[3250]),

			.SO(gen[3343]),
			.S(gen[3344]),
			.SE(gen[3345]),

			.SELF(gen[3249]),
			.cell_state(gen[3249])
		); 

/******************* CELL 3250 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3250 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3154]),
			.N(gen[3155]),
			.NE(gen[3156]),

			.O(gen[3249]),
			.E(gen[3251]),

			.SO(gen[3344]),
			.S(gen[3345]),
			.SE(gen[3346]),

			.SELF(gen[3250]),
			.cell_state(gen[3250])
		); 

/******************* CELL 3251 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3251 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3155]),
			.N(gen[3156]),
			.NE(gen[3157]),

			.O(gen[3250]),
			.E(gen[3252]),

			.SO(gen[3345]),
			.S(gen[3346]),
			.SE(gen[3347]),

			.SELF(gen[3251]),
			.cell_state(gen[3251])
		); 

/******************* CELL 3252 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3252 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3156]),
			.N(gen[3157]),
			.NE(gen[3158]),

			.O(gen[3251]),
			.E(gen[3253]),

			.SO(gen[3346]),
			.S(gen[3347]),
			.SE(gen[3348]),

			.SELF(gen[3252]),
			.cell_state(gen[3252])
		); 

/******************* CELL 3253 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3253 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3157]),
			.N(gen[3158]),
			.NE(gen[3159]),

			.O(gen[3252]),
			.E(gen[3254]),

			.SO(gen[3347]),
			.S(gen[3348]),
			.SE(gen[3349]),

			.SELF(gen[3253]),
			.cell_state(gen[3253])
		); 

/******************* CELL 3254 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3254 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3158]),
			.N(gen[3159]),
			.NE(gen[3160]),

			.O(gen[3253]),
			.E(gen[3255]),

			.SO(gen[3348]),
			.S(gen[3349]),
			.SE(gen[3350]),

			.SELF(gen[3254]),
			.cell_state(gen[3254])
		); 

/******************* CELL 3255 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3255 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3159]),
			.N(gen[3160]),
			.NE(gen[3161]),

			.O(gen[3254]),
			.E(gen[3256]),

			.SO(gen[3349]),
			.S(gen[3350]),
			.SE(gen[3351]),

			.SELF(gen[3255]),
			.cell_state(gen[3255])
		); 

/******************* CELL 3256 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3256 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3160]),
			.N(gen[3161]),
			.NE(gen[3162]),

			.O(gen[3255]),
			.E(gen[3257]),

			.SO(gen[3350]),
			.S(gen[3351]),
			.SE(gen[3352]),

			.SELF(gen[3256]),
			.cell_state(gen[3256])
		); 

/******************* CELL 3257 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3257 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3161]),
			.N(gen[3162]),
			.NE(gen[3163]),

			.O(gen[3256]),
			.E(gen[3258]),

			.SO(gen[3351]),
			.S(gen[3352]),
			.SE(gen[3353]),

			.SELF(gen[3257]),
			.cell_state(gen[3257])
		); 

/******************* CELL 3258 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3258 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3162]),
			.N(gen[3163]),
			.NE(gen[3164]),

			.O(gen[3257]),
			.E(gen[3259]),

			.SO(gen[3352]),
			.S(gen[3353]),
			.SE(gen[3354]),

			.SELF(gen[3258]),
			.cell_state(gen[3258])
		); 

/******************* CELL 3259 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3259 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3163]),
			.N(gen[3164]),
			.NE(gen[3165]),

			.O(gen[3258]),
			.E(gen[3260]),

			.SO(gen[3353]),
			.S(gen[3354]),
			.SE(gen[3355]),

			.SELF(gen[3259]),
			.cell_state(gen[3259])
		); 

/******************* CELL 3260 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3260 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3164]),
			.N(gen[3165]),
			.NE(gen[3166]),

			.O(gen[3259]),
			.E(gen[3261]),

			.SO(gen[3354]),
			.S(gen[3355]),
			.SE(gen[3356]),

			.SELF(gen[3260]),
			.cell_state(gen[3260])
		); 

/******************* CELL 3261 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3261 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3165]),
			.N(gen[3166]),
			.NE(gen[3167]),

			.O(gen[3260]),
			.E(gen[3262]),

			.SO(gen[3355]),
			.S(gen[3356]),
			.SE(gen[3357]),

			.SELF(gen[3261]),
			.cell_state(gen[3261])
		); 

/******************* CELL 3262 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3262 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3166]),
			.N(gen[3167]),
			.NE(gen[3168]),

			.O(gen[3261]),
			.E(gen[3263]),

			.SO(gen[3356]),
			.S(gen[3357]),
			.SE(gen[3358]),

			.SELF(gen[3262]),
			.cell_state(gen[3262])
		); 

/******************* CELL 3263 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3263 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3167]),
			.N(gen[3168]),
			.NE(gen[3169]),

			.O(gen[3262]),
			.E(gen[3264]),

			.SO(gen[3357]),
			.S(gen[3358]),
			.SE(gen[3359]),

			.SELF(gen[3263]),
			.cell_state(gen[3263])
		); 

/******************* CELL 3264 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3264 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3168]),
			.N(gen[3169]),
			.NE(gen[3170]),

			.O(gen[3263]),
			.E(gen[3265]),

			.SO(gen[3358]),
			.S(gen[3359]),
			.SE(gen[3360]),

			.SELF(gen[3264]),
			.cell_state(gen[3264])
		); 

/******************* CELL 3265 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3265 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3169]),
			.N(gen[3170]),
			.NE(gen[3171]),

			.O(gen[3264]),
			.E(gen[3266]),

			.SO(gen[3359]),
			.S(gen[3360]),
			.SE(gen[3361]),

			.SELF(gen[3265]),
			.cell_state(gen[3265])
		); 

/******************* CELL 3266 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3266 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3170]),
			.N(gen[3171]),
			.NE(gen[3172]),

			.O(gen[3265]),
			.E(gen[3267]),

			.SO(gen[3360]),
			.S(gen[3361]),
			.SE(gen[3362]),

			.SELF(gen[3266]),
			.cell_state(gen[3266])
		); 

/******************* CELL 3267 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3267 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3171]),
			.N(gen[3172]),
			.NE(gen[3173]),

			.O(gen[3266]),
			.E(gen[3268]),

			.SO(gen[3361]),
			.S(gen[3362]),
			.SE(gen[3363]),

			.SELF(gen[3267]),
			.cell_state(gen[3267])
		); 

/******************* CELL 3268 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3268 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3172]),
			.N(gen[3173]),
			.NE(gen[3174]),

			.O(gen[3267]),
			.E(gen[3269]),

			.SO(gen[3362]),
			.S(gen[3363]),
			.SE(gen[3364]),

			.SELF(gen[3268]),
			.cell_state(gen[3268])
		); 

/******************* CELL 3269 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3269 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3173]),
			.N(gen[3174]),
			.NE(gen[3175]),

			.O(gen[3268]),
			.E(gen[3270]),

			.SO(gen[3363]),
			.S(gen[3364]),
			.SE(gen[3365]),

			.SELF(gen[3269]),
			.cell_state(gen[3269])
		); 

/******************* CELL 3270 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3270 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3174]),
			.N(gen[3175]),
			.NE(gen[3176]),

			.O(gen[3269]),
			.E(gen[3271]),

			.SO(gen[3364]),
			.S(gen[3365]),
			.SE(gen[3366]),

			.SELF(gen[3270]),
			.cell_state(gen[3270])
		); 

/******************* CELL 3271 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3271 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3175]),
			.N(gen[3176]),
			.NE(gen[3177]),

			.O(gen[3270]),
			.E(gen[3272]),

			.SO(gen[3365]),
			.S(gen[3366]),
			.SE(gen[3367]),

			.SELF(gen[3271]),
			.cell_state(gen[3271])
		); 

/******************* CELL 3272 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3272 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3176]),
			.N(gen[3177]),
			.NE(gen[3178]),

			.O(gen[3271]),
			.E(gen[3273]),

			.SO(gen[3366]),
			.S(gen[3367]),
			.SE(gen[3368]),

			.SELF(gen[3272]),
			.cell_state(gen[3272])
		); 

/******************* CELL 3273 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3273 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3177]),
			.N(gen[3178]),
			.NE(gen[3179]),

			.O(gen[3272]),
			.E(gen[3274]),

			.SO(gen[3367]),
			.S(gen[3368]),
			.SE(gen[3369]),

			.SELF(gen[3273]),
			.cell_state(gen[3273])
		); 

/******************* CELL 3274 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3274 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3178]),
			.N(gen[3179]),
			.NE(gen[3180]),

			.O(gen[3273]),
			.E(gen[3275]),

			.SO(gen[3368]),
			.S(gen[3369]),
			.SE(gen[3370]),

			.SELF(gen[3274]),
			.cell_state(gen[3274])
		); 

/******************* CELL 3275 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3275 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3179]),
			.N(gen[3180]),
			.NE(gen[3181]),

			.O(gen[3274]),
			.E(gen[3276]),

			.SO(gen[3369]),
			.S(gen[3370]),
			.SE(gen[3371]),

			.SELF(gen[3275]),
			.cell_state(gen[3275])
		); 

/******************* CELL 3276 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3276 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3180]),
			.N(gen[3181]),
			.NE(gen[3182]),

			.O(gen[3275]),
			.E(gen[3277]),

			.SO(gen[3370]),
			.S(gen[3371]),
			.SE(gen[3372]),

			.SELF(gen[3276]),
			.cell_state(gen[3276])
		); 

/******************* CELL 3277 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3277 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3181]),
			.N(gen[3182]),
			.NE(gen[3183]),

			.O(gen[3276]),
			.E(gen[3278]),

			.SO(gen[3371]),
			.S(gen[3372]),
			.SE(gen[3373]),

			.SELF(gen[3277]),
			.cell_state(gen[3277])
		); 

/******************* CELL 3278 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3278 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3182]),
			.N(gen[3183]),
			.NE(gen[3184]),

			.O(gen[3277]),
			.E(gen[3279]),

			.SO(gen[3372]),
			.S(gen[3373]),
			.SE(gen[3374]),

			.SELF(gen[3278]),
			.cell_state(gen[3278])
		); 

/******************* CELL 3279 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3279 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3183]),
			.N(gen[3184]),
			.NE(gen[3185]),

			.O(gen[3278]),
			.E(gen[3280]),

			.SO(gen[3373]),
			.S(gen[3374]),
			.SE(gen[3375]),

			.SELF(gen[3279]),
			.cell_state(gen[3279])
		); 

/******************* CELL 3280 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3280 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3184]),
			.N(gen[3185]),
			.NE(gen[3186]),

			.O(gen[3279]),
			.E(gen[3281]),

			.SO(gen[3374]),
			.S(gen[3375]),
			.SE(gen[3376]),

			.SELF(gen[3280]),
			.cell_state(gen[3280])
		); 

/******************* CELL 3281 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3281 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3185]),
			.N(gen[3186]),
			.NE(gen[3187]),

			.O(gen[3280]),
			.E(gen[3282]),

			.SO(gen[3375]),
			.S(gen[3376]),
			.SE(gen[3377]),

			.SELF(gen[3281]),
			.cell_state(gen[3281])
		); 

/******************* CELL 3282 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3282 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3186]),
			.N(gen[3187]),
			.NE(gen[3188]),

			.O(gen[3281]),
			.E(gen[3283]),

			.SO(gen[3376]),
			.S(gen[3377]),
			.SE(gen[3378]),

			.SELF(gen[3282]),
			.cell_state(gen[3282])
		); 

/******************* CELL 3283 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3283 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3187]),
			.N(gen[3188]),
			.NE(gen[3189]),

			.O(gen[3282]),
			.E(gen[3284]),

			.SO(gen[3377]),
			.S(gen[3378]),
			.SE(gen[3379]),

			.SELF(gen[3283]),
			.cell_state(gen[3283])
		); 

/******************* CELL 3284 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3284 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3188]),
			.N(gen[3189]),
			.NE(gen[3190]),

			.O(gen[3283]),
			.E(gen[3285]),

			.SO(gen[3378]),
			.S(gen[3379]),
			.SE(gen[3380]),

			.SELF(gen[3284]),
			.cell_state(gen[3284])
		); 

/******************* CELL 3285 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3285 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3189]),
			.N(gen[3190]),
			.NE(gen[3191]),

			.O(gen[3284]),
			.E(gen[3286]),

			.SO(gen[3379]),
			.S(gen[3380]),
			.SE(gen[3381]),

			.SELF(gen[3285]),
			.cell_state(gen[3285])
		); 

/******************* CELL 3286 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3286 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3190]),
			.N(gen[3191]),
			.NE(gen[3192]),

			.O(gen[3285]),
			.E(gen[3287]),

			.SO(gen[3380]),
			.S(gen[3381]),
			.SE(gen[3382]),

			.SELF(gen[3286]),
			.cell_state(gen[3286])
		); 

/******************* CELL 3287 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3287 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3191]),
			.N(gen[3192]),
			.NE(gen[3193]),

			.O(gen[3286]),
			.E(gen[3288]),

			.SO(gen[3381]),
			.S(gen[3382]),
			.SE(gen[3383]),

			.SELF(gen[3287]),
			.cell_state(gen[3287])
		); 

/******************* CELL 3288 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3288 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3192]),
			.N(gen[3193]),
			.NE(gen[3194]),

			.O(gen[3287]),
			.E(gen[3289]),

			.SO(gen[3382]),
			.S(gen[3383]),
			.SE(gen[3384]),

			.SELF(gen[3288]),
			.cell_state(gen[3288])
		); 

/******************* CELL 3289 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3289 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3193]),
			.N(gen[3194]),
			.NE(gen[3195]),

			.O(gen[3288]),
			.E(gen[3290]),

			.SO(gen[3383]),
			.S(gen[3384]),
			.SE(gen[3385]),

			.SELF(gen[3289]),
			.cell_state(gen[3289])
		); 

/******************* CELL 3290 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3290 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3194]),
			.N(gen[3195]),
			.NE(gen[3196]),

			.O(gen[3289]),
			.E(gen[3291]),

			.SO(gen[3384]),
			.S(gen[3385]),
			.SE(gen[3386]),

			.SELF(gen[3290]),
			.cell_state(gen[3290])
		); 

/******************* CELL 3291 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3291 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3195]),
			.N(gen[3196]),
			.NE(gen[3197]),

			.O(gen[3290]),
			.E(gen[3292]),

			.SO(gen[3385]),
			.S(gen[3386]),
			.SE(gen[3387]),

			.SELF(gen[3291]),
			.cell_state(gen[3291])
		); 

/******************* CELL 3292 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3292 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3196]),
			.N(gen[3197]),
			.NE(gen[3198]),

			.O(gen[3291]),
			.E(gen[3293]),

			.SO(gen[3386]),
			.S(gen[3387]),
			.SE(gen[3388]),

			.SELF(gen[3292]),
			.cell_state(gen[3292])
		); 

/******************* CELL 3293 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3293 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3197]),
			.N(gen[3198]),
			.NE(gen[3199]),

			.O(gen[3292]),
			.E(gen[3294]),

			.SO(gen[3387]),
			.S(gen[3388]),
			.SE(gen[3389]),

			.SELF(gen[3293]),
			.cell_state(gen[3293])
		); 

/******************* CELL 3294 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3294 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3198]),
			.N(gen[3199]),
			.NE(gen[3200]),

			.O(gen[3293]),
			.E(gen[3295]),

			.SO(gen[3388]),
			.S(gen[3389]),
			.SE(gen[3390]),

			.SELF(gen[3294]),
			.cell_state(gen[3294])
		); 

/******************* CELL 3295 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3295 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3199]),
			.N(gen[3200]),
			.NE(gen[3201]),

			.O(gen[3294]),
			.E(gen[3296]),

			.SO(gen[3389]),
			.S(gen[3390]),
			.SE(gen[3391]),

			.SELF(gen[3295]),
			.cell_state(gen[3295])
		); 

/******************* CELL 3296 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3296 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3200]),
			.N(gen[3201]),
			.NE(gen[3202]),

			.O(gen[3295]),
			.E(gen[3297]),

			.SO(gen[3390]),
			.S(gen[3391]),
			.SE(gen[3392]),

			.SELF(gen[3296]),
			.cell_state(gen[3296])
		); 

/******************* CELL 3297 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3297 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3201]),
			.N(gen[3202]),
			.NE(gen[3203]),

			.O(gen[3296]),
			.E(gen[3298]),

			.SO(gen[3391]),
			.S(gen[3392]),
			.SE(gen[3393]),

			.SELF(gen[3297]),
			.cell_state(gen[3297])
		); 

/******************* CELL 3298 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3298 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3202]),
			.N(gen[3203]),
			.NE(gen[3204]),

			.O(gen[3297]),
			.E(gen[3299]),

			.SO(gen[3392]),
			.S(gen[3393]),
			.SE(gen[3394]),

			.SELF(gen[3298]),
			.cell_state(gen[3298])
		); 

/******************* CELL 3299 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3299 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3203]),
			.N(gen[3204]),
			.NE(gen[3205]),

			.O(gen[3298]),
			.E(gen[3300]),

			.SO(gen[3393]),
			.S(gen[3394]),
			.SE(gen[3395]),

			.SELF(gen[3299]),
			.cell_state(gen[3299])
		); 

/******************* CELL 3300 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3300 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3204]),
			.N(gen[3205]),
			.NE(gen[3206]),

			.O(gen[3299]),
			.E(gen[3301]),

			.SO(gen[3394]),
			.S(gen[3395]),
			.SE(gen[3396]),

			.SELF(gen[3300]),
			.cell_state(gen[3300])
		); 

/******************* CELL 3301 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3301 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3205]),
			.N(gen[3206]),
			.NE(gen[3207]),

			.O(gen[3300]),
			.E(gen[3302]),

			.SO(gen[3395]),
			.S(gen[3396]),
			.SE(gen[3397]),

			.SELF(gen[3301]),
			.cell_state(gen[3301])
		); 

/******************* CELL 3302 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3302 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3206]),
			.N(gen[3207]),
			.NE(gen[3208]),

			.O(gen[3301]),
			.E(gen[3303]),

			.SO(gen[3396]),
			.S(gen[3397]),
			.SE(gen[3398]),

			.SELF(gen[3302]),
			.cell_state(gen[3302])
		); 

/******************* CELL 3303 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3303 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3207]),
			.N(gen[3208]),
			.NE(gen[3209]),

			.O(gen[3302]),
			.E(gen[3304]),

			.SO(gen[3397]),
			.S(gen[3398]),
			.SE(gen[3399]),

			.SELF(gen[3303]),
			.cell_state(gen[3303])
		); 

/******************* CELL 3304 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3304 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3208]),
			.N(gen[3209]),
			.NE(gen[3210]),

			.O(gen[3303]),
			.E(gen[3305]),

			.SO(gen[3398]),
			.S(gen[3399]),
			.SE(gen[3400]),

			.SELF(gen[3304]),
			.cell_state(gen[3304])
		); 

/******************* CELL 3305 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3305 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3209]),
			.N(gen[3210]),
			.NE(gen[3211]),

			.O(gen[3304]),
			.E(gen[3306]),

			.SO(gen[3399]),
			.S(gen[3400]),
			.SE(gen[3401]),

			.SELF(gen[3305]),
			.cell_state(gen[3305])
		); 

/******************* CELL 3306 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3306 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3210]),
			.N(gen[3211]),
			.NE(gen[3212]),

			.O(gen[3305]),
			.E(gen[3307]),

			.SO(gen[3400]),
			.S(gen[3401]),
			.SE(gen[3402]),

			.SELF(gen[3306]),
			.cell_state(gen[3306])
		); 

/******************* CELL 3307 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3307 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3211]),
			.N(gen[3212]),
			.NE(gen[3213]),

			.O(gen[3306]),
			.E(gen[3308]),

			.SO(gen[3401]),
			.S(gen[3402]),
			.SE(gen[3403]),

			.SELF(gen[3307]),
			.cell_state(gen[3307])
		); 

/******************* CELL 3308 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3308 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3212]),
			.N(gen[3213]),
			.NE(gen[3214]),

			.O(gen[3307]),
			.E(gen[3309]),

			.SO(gen[3402]),
			.S(gen[3403]),
			.SE(gen[3404]),

			.SELF(gen[3308]),
			.cell_state(gen[3308])
		); 

/******************* CELL 3309 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3309 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3213]),
			.N(gen[3214]),
			.NE(gen[3215]),

			.O(gen[3308]),
			.E(gen[3310]),

			.SO(gen[3403]),
			.S(gen[3404]),
			.SE(gen[3405]),

			.SELF(gen[3309]),
			.cell_state(gen[3309])
		); 

/******************* CELL 3310 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3310 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3214]),
			.N(gen[3215]),
			.NE(gen[3216]),

			.O(gen[3309]),
			.E(gen[3311]),

			.SO(gen[3404]),
			.S(gen[3405]),
			.SE(gen[3406]),

			.SELF(gen[3310]),
			.cell_state(gen[3310])
		); 

/******************* CELL 3311 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3311 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3215]),
			.N(gen[3216]),
			.NE(gen[3217]),

			.O(gen[3310]),
			.E(gen[3312]),

			.SO(gen[3405]),
			.S(gen[3406]),
			.SE(gen[3407]),

			.SELF(gen[3311]),
			.cell_state(gen[3311])
		); 

/******************* CELL 3312 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3312 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3216]),
			.N(gen[3217]),
			.NE(gen[3218]),

			.O(gen[3311]),
			.E(gen[3313]),

			.SO(gen[3406]),
			.S(gen[3407]),
			.SE(gen[3408]),

			.SELF(gen[3312]),
			.cell_state(gen[3312])
		); 

/******************* CELL 3313 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3313 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3217]),
			.N(gen[3218]),
			.NE(gen[3219]),

			.O(gen[3312]),
			.E(gen[3314]),

			.SO(gen[3407]),
			.S(gen[3408]),
			.SE(gen[3409]),

			.SELF(gen[3313]),
			.cell_state(gen[3313])
		); 

/******************* CELL 3314 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3314 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3218]),
			.N(gen[3219]),
			.NE(gen[3220]),

			.O(gen[3313]),
			.E(gen[3315]),

			.SO(gen[3408]),
			.S(gen[3409]),
			.SE(gen[3410]),

			.SELF(gen[3314]),
			.cell_state(gen[3314])
		); 

/******************* CELL 3315 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3315 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3219]),
			.N(gen[3220]),
			.NE(gen[3221]),

			.O(gen[3314]),
			.E(gen[3316]),

			.SO(gen[3409]),
			.S(gen[3410]),
			.SE(gen[3411]),

			.SELF(gen[3315]),
			.cell_state(gen[3315])
		); 

/******************* CELL 3316 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3316 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3220]),
			.N(gen[3221]),
			.NE(gen[3222]),

			.O(gen[3315]),
			.E(gen[3317]),

			.SO(gen[3410]),
			.S(gen[3411]),
			.SE(gen[3412]),

			.SELF(gen[3316]),
			.cell_state(gen[3316])
		); 

/******************* CELL 3317 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3317 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3221]),
			.N(gen[3222]),
			.NE(gen[3223]),

			.O(gen[3316]),
			.E(gen[3318]),

			.SO(gen[3411]),
			.S(gen[3412]),
			.SE(gen[3413]),

			.SELF(gen[3317]),
			.cell_state(gen[3317])
		); 

/******************* CELL 3318 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3318 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3222]),
			.N(gen[3223]),
			.NE(gen[3224]),

			.O(gen[3317]),
			.E(gen[3319]),

			.SO(gen[3412]),
			.S(gen[3413]),
			.SE(gen[3414]),

			.SELF(gen[3318]),
			.cell_state(gen[3318])
		); 

/******************* CELL 3319 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3319 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3223]),
			.N(gen[3224]),
			.NE(gen[3225]),

			.O(gen[3318]),
			.E(gen[3320]),

			.SO(gen[3413]),
			.S(gen[3414]),
			.SE(gen[3415]),

			.SELF(gen[3319]),
			.cell_state(gen[3319])
		); 

/******************* CELL 3320 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3320 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3224]),
			.N(gen[3225]),
			.NE(gen[3226]),

			.O(gen[3319]),
			.E(gen[3321]),

			.SO(gen[3414]),
			.S(gen[3415]),
			.SE(gen[3416]),

			.SELF(gen[3320]),
			.cell_state(gen[3320])
		); 

/******************* CELL 3321 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3321 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3225]),
			.N(gen[3226]),
			.NE(gen[3227]),

			.O(gen[3320]),
			.E(gen[3322]),

			.SO(gen[3415]),
			.S(gen[3416]),
			.SE(gen[3417]),

			.SELF(gen[3321]),
			.cell_state(gen[3321])
		); 

/******************* CELL 3322 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3322 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3226]),
			.N(gen[3227]),
			.NE(gen[3228]),

			.O(gen[3321]),
			.E(gen[3323]),

			.SO(gen[3416]),
			.S(gen[3417]),
			.SE(gen[3418]),

			.SELF(gen[3322]),
			.cell_state(gen[3322])
		); 

/******************* CELL 3323 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3323 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3227]),
			.N(gen[3228]),
			.NE(gen[3229]),

			.O(gen[3322]),
			.E(gen[3324]),

			.SO(gen[3417]),
			.S(gen[3418]),
			.SE(gen[3419]),

			.SELF(gen[3323]),
			.cell_state(gen[3323])
		); 

/******************* CELL 3324 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3324 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3228]),
			.N(gen[3229]),
			.NE(gen[3228]),

			.O(gen[3323]),
			.E(gen[3323]),

			.SO(gen[3418]),
			.S(gen[3419]),
			.SE(gen[3418]),

			.SELF(gen[3324]),
			.cell_state(gen[3324])
		); 

/******************* CELL 3325 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3325 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3231]),
			.N(gen[3230]),
			.NE(gen[3231]),

			.O(gen[3326]),
			.E(gen[3326]),

			.SO(gen[3421]),
			.S(gen[3420]),
			.SE(gen[3421]),

			.SELF(gen[3325]),
			.cell_state(gen[3325])
		); 

/******************* CELL 3326 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3326 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3230]),
			.N(gen[3231]),
			.NE(gen[3232]),

			.O(gen[3325]),
			.E(gen[3327]),

			.SO(gen[3420]),
			.S(gen[3421]),
			.SE(gen[3422]),

			.SELF(gen[3326]),
			.cell_state(gen[3326])
		); 

/******************* CELL 3327 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3327 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3231]),
			.N(gen[3232]),
			.NE(gen[3233]),

			.O(gen[3326]),
			.E(gen[3328]),

			.SO(gen[3421]),
			.S(gen[3422]),
			.SE(gen[3423]),

			.SELF(gen[3327]),
			.cell_state(gen[3327])
		); 

/******************* CELL 3328 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3328 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3232]),
			.N(gen[3233]),
			.NE(gen[3234]),

			.O(gen[3327]),
			.E(gen[3329]),

			.SO(gen[3422]),
			.S(gen[3423]),
			.SE(gen[3424]),

			.SELF(gen[3328]),
			.cell_state(gen[3328])
		); 

/******************* CELL 3329 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3329 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3233]),
			.N(gen[3234]),
			.NE(gen[3235]),

			.O(gen[3328]),
			.E(gen[3330]),

			.SO(gen[3423]),
			.S(gen[3424]),
			.SE(gen[3425]),

			.SELF(gen[3329]),
			.cell_state(gen[3329])
		); 

/******************* CELL 3330 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3330 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3234]),
			.N(gen[3235]),
			.NE(gen[3236]),

			.O(gen[3329]),
			.E(gen[3331]),

			.SO(gen[3424]),
			.S(gen[3425]),
			.SE(gen[3426]),

			.SELF(gen[3330]),
			.cell_state(gen[3330])
		); 

/******************* CELL 3331 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3331 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3235]),
			.N(gen[3236]),
			.NE(gen[3237]),

			.O(gen[3330]),
			.E(gen[3332]),

			.SO(gen[3425]),
			.S(gen[3426]),
			.SE(gen[3427]),

			.SELF(gen[3331]),
			.cell_state(gen[3331])
		); 

/******************* CELL 3332 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3332 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3236]),
			.N(gen[3237]),
			.NE(gen[3238]),

			.O(gen[3331]),
			.E(gen[3333]),

			.SO(gen[3426]),
			.S(gen[3427]),
			.SE(gen[3428]),

			.SELF(gen[3332]),
			.cell_state(gen[3332])
		); 

/******************* CELL 3333 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3333 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3237]),
			.N(gen[3238]),
			.NE(gen[3239]),

			.O(gen[3332]),
			.E(gen[3334]),

			.SO(gen[3427]),
			.S(gen[3428]),
			.SE(gen[3429]),

			.SELF(gen[3333]),
			.cell_state(gen[3333])
		); 

/******************* CELL 3334 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3334 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3238]),
			.N(gen[3239]),
			.NE(gen[3240]),

			.O(gen[3333]),
			.E(gen[3335]),

			.SO(gen[3428]),
			.S(gen[3429]),
			.SE(gen[3430]),

			.SELF(gen[3334]),
			.cell_state(gen[3334])
		); 

/******************* CELL 3335 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3335 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3239]),
			.N(gen[3240]),
			.NE(gen[3241]),

			.O(gen[3334]),
			.E(gen[3336]),

			.SO(gen[3429]),
			.S(gen[3430]),
			.SE(gen[3431]),

			.SELF(gen[3335]),
			.cell_state(gen[3335])
		); 

/******************* CELL 3336 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3336 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3240]),
			.N(gen[3241]),
			.NE(gen[3242]),

			.O(gen[3335]),
			.E(gen[3337]),

			.SO(gen[3430]),
			.S(gen[3431]),
			.SE(gen[3432]),

			.SELF(gen[3336]),
			.cell_state(gen[3336])
		); 

/******************* CELL 3337 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3337 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3241]),
			.N(gen[3242]),
			.NE(gen[3243]),

			.O(gen[3336]),
			.E(gen[3338]),

			.SO(gen[3431]),
			.S(gen[3432]),
			.SE(gen[3433]),

			.SELF(gen[3337]),
			.cell_state(gen[3337])
		); 

/******************* CELL 3338 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3338 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3242]),
			.N(gen[3243]),
			.NE(gen[3244]),

			.O(gen[3337]),
			.E(gen[3339]),

			.SO(gen[3432]),
			.S(gen[3433]),
			.SE(gen[3434]),

			.SELF(gen[3338]),
			.cell_state(gen[3338])
		); 

/******************* CELL 3339 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3339 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3243]),
			.N(gen[3244]),
			.NE(gen[3245]),

			.O(gen[3338]),
			.E(gen[3340]),

			.SO(gen[3433]),
			.S(gen[3434]),
			.SE(gen[3435]),

			.SELF(gen[3339]),
			.cell_state(gen[3339])
		); 

/******************* CELL 3340 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3340 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3244]),
			.N(gen[3245]),
			.NE(gen[3246]),

			.O(gen[3339]),
			.E(gen[3341]),

			.SO(gen[3434]),
			.S(gen[3435]),
			.SE(gen[3436]),

			.SELF(gen[3340]),
			.cell_state(gen[3340])
		); 

/******************* CELL 3341 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3341 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3245]),
			.N(gen[3246]),
			.NE(gen[3247]),

			.O(gen[3340]),
			.E(gen[3342]),

			.SO(gen[3435]),
			.S(gen[3436]),
			.SE(gen[3437]),

			.SELF(gen[3341]),
			.cell_state(gen[3341])
		); 

/******************* CELL 3342 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3342 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3246]),
			.N(gen[3247]),
			.NE(gen[3248]),

			.O(gen[3341]),
			.E(gen[3343]),

			.SO(gen[3436]),
			.S(gen[3437]),
			.SE(gen[3438]),

			.SELF(gen[3342]),
			.cell_state(gen[3342])
		); 

/******************* CELL 3343 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3343 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3247]),
			.N(gen[3248]),
			.NE(gen[3249]),

			.O(gen[3342]),
			.E(gen[3344]),

			.SO(gen[3437]),
			.S(gen[3438]),
			.SE(gen[3439]),

			.SELF(gen[3343]),
			.cell_state(gen[3343])
		); 

/******************* CELL 3344 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3344 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3248]),
			.N(gen[3249]),
			.NE(gen[3250]),

			.O(gen[3343]),
			.E(gen[3345]),

			.SO(gen[3438]),
			.S(gen[3439]),
			.SE(gen[3440]),

			.SELF(gen[3344]),
			.cell_state(gen[3344])
		); 

/******************* CELL 3345 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3345 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3249]),
			.N(gen[3250]),
			.NE(gen[3251]),

			.O(gen[3344]),
			.E(gen[3346]),

			.SO(gen[3439]),
			.S(gen[3440]),
			.SE(gen[3441]),

			.SELF(gen[3345]),
			.cell_state(gen[3345])
		); 

/******************* CELL 3346 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3346 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3250]),
			.N(gen[3251]),
			.NE(gen[3252]),

			.O(gen[3345]),
			.E(gen[3347]),

			.SO(gen[3440]),
			.S(gen[3441]),
			.SE(gen[3442]),

			.SELF(gen[3346]),
			.cell_state(gen[3346])
		); 

/******************* CELL 3347 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3347 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3251]),
			.N(gen[3252]),
			.NE(gen[3253]),

			.O(gen[3346]),
			.E(gen[3348]),

			.SO(gen[3441]),
			.S(gen[3442]),
			.SE(gen[3443]),

			.SELF(gen[3347]),
			.cell_state(gen[3347])
		); 

/******************* CELL 3348 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3348 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3252]),
			.N(gen[3253]),
			.NE(gen[3254]),

			.O(gen[3347]),
			.E(gen[3349]),

			.SO(gen[3442]),
			.S(gen[3443]),
			.SE(gen[3444]),

			.SELF(gen[3348]),
			.cell_state(gen[3348])
		); 

/******************* CELL 3349 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3349 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3253]),
			.N(gen[3254]),
			.NE(gen[3255]),

			.O(gen[3348]),
			.E(gen[3350]),

			.SO(gen[3443]),
			.S(gen[3444]),
			.SE(gen[3445]),

			.SELF(gen[3349]),
			.cell_state(gen[3349])
		); 

/******************* CELL 3350 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3350 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3254]),
			.N(gen[3255]),
			.NE(gen[3256]),

			.O(gen[3349]),
			.E(gen[3351]),

			.SO(gen[3444]),
			.S(gen[3445]),
			.SE(gen[3446]),

			.SELF(gen[3350]),
			.cell_state(gen[3350])
		); 

/******************* CELL 3351 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3351 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3255]),
			.N(gen[3256]),
			.NE(gen[3257]),

			.O(gen[3350]),
			.E(gen[3352]),

			.SO(gen[3445]),
			.S(gen[3446]),
			.SE(gen[3447]),

			.SELF(gen[3351]),
			.cell_state(gen[3351])
		); 

/******************* CELL 3352 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3352 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3256]),
			.N(gen[3257]),
			.NE(gen[3258]),

			.O(gen[3351]),
			.E(gen[3353]),

			.SO(gen[3446]),
			.S(gen[3447]),
			.SE(gen[3448]),

			.SELF(gen[3352]),
			.cell_state(gen[3352])
		); 

/******************* CELL 3353 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3353 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3257]),
			.N(gen[3258]),
			.NE(gen[3259]),

			.O(gen[3352]),
			.E(gen[3354]),

			.SO(gen[3447]),
			.S(gen[3448]),
			.SE(gen[3449]),

			.SELF(gen[3353]),
			.cell_state(gen[3353])
		); 

/******************* CELL 3354 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3354 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3258]),
			.N(gen[3259]),
			.NE(gen[3260]),

			.O(gen[3353]),
			.E(gen[3355]),

			.SO(gen[3448]),
			.S(gen[3449]),
			.SE(gen[3450]),

			.SELF(gen[3354]),
			.cell_state(gen[3354])
		); 

/******************* CELL 3355 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3355 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3259]),
			.N(gen[3260]),
			.NE(gen[3261]),

			.O(gen[3354]),
			.E(gen[3356]),

			.SO(gen[3449]),
			.S(gen[3450]),
			.SE(gen[3451]),

			.SELF(gen[3355]),
			.cell_state(gen[3355])
		); 

/******************* CELL 3356 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3356 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3260]),
			.N(gen[3261]),
			.NE(gen[3262]),

			.O(gen[3355]),
			.E(gen[3357]),

			.SO(gen[3450]),
			.S(gen[3451]),
			.SE(gen[3452]),

			.SELF(gen[3356]),
			.cell_state(gen[3356])
		); 

/******************* CELL 3357 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3357 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3261]),
			.N(gen[3262]),
			.NE(gen[3263]),

			.O(gen[3356]),
			.E(gen[3358]),

			.SO(gen[3451]),
			.S(gen[3452]),
			.SE(gen[3453]),

			.SELF(gen[3357]),
			.cell_state(gen[3357])
		); 

/******************* CELL 3358 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3358 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3262]),
			.N(gen[3263]),
			.NE(gen[3264]),

			.O(gen[3357]),
			.E(gen[3359]),

			.SO(gen[3452]),
			.S(gen[3453]),
			.SE(gen[3454]),

			.SELF(gen[3358]),
			.cell_state(gen[3358])
		); 

/******************* CELL 3359 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3359 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3263]),
			.N(gen[3264]),
			.NE(gen[3265]),

			.O(gen[3358]),
			.E(gen[3360]),

			.SO(gen[3453]),
			.S(gen[3454]),
			.SE(gen[3455]),

			.SELF(gen[3359]),
			.cell_state(gen[3359])
		); 

/******************* CELL 3360 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3360 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3264]),
			.N(gen[3265]),
			.NE(gen[3266]),

			.O(gen[3359]),
			.E(gen[3361]),

			.SO(gen[3454]),
			.S(gen[3455]),
			.SE(gen[3456]),

			.SELF(gen[3360]),
			.cell_state(gen[3360])
		); 

/******************* CELL 3361 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3361 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3265]),
			.N(gen[3266]),
			.NE(gen[3267]),

			.O(gen[3360]),
			.E(gen[3362]),

			.SO(gen[3455]),
			.S(gen[3456]),
			.SE(gen[3457]),

			.SELF(gen[3361]),
			.cell_state(gen[3361])
		); 

/******************* CELL 3362 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3362 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3266]),
			.N(gen[3267]),
			.NE(gen[3268]),

			.O(gen[3361]),
			.E(gen[3363]),

			.SO(gen[3456]),
			.S(gen[3457]),
			.SE(gen[3458]),

			.SELF(gen[3362]),
			.cell_state(gen[3362])
		); 

/******************* CELL 3363 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3363 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3267]),
			.N(gen[3268]),
			.NE(gen[3269]),

			.O(gen[3362]),
			.E(gen[3364]),

			.SO(gen[3457]),
			.S(gen[3458]),
			.SE(gen[3459]),

			.SELF(gen[3363]),
			.cell_state(gen[3363])
		); 

/******************* CELL 3364 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3364 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3268]),
			.N(gen[3269]),
			.NE(gen[3270]),

			.O(gen[3363]),
			.E(gen[3365]),

			.SO(gen[3458]),
			.S(gen[3459]),
			.SE(gen[3460]),

			.SELF(gen[3364]),
			.cell_state(gen[3364])
		); 

/******************* CELL 3365 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3365 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3269]),
			.N(gen[3270]),
			.NE(gen[3271]),

			.O(gen[3364]),
			.E(gen[3366]),

			.SO(gen[3459]),
			.S(gen[3460]),
			.SE(gen[3461]),

			.SELF(gen[3365]),
			.cell_state(gen[3365])
		); 

/******************* CELL 3366 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3366 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3270]),
			.N(gen[3271]),
			.NE(gen[3272]),

			.O(gen[3365]),
			.E(gen[3367]),

			.SO(gen[3460]),
			.S(gen[3461]),
			.SE(gen[3462]),

			.SELF(gen[3366]),
			.cell_state(gen[3366])
		); 

/******************* CELL 3367 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3367 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3271]),
			.N(gen[3272]),
			.NE(gen[3273]),

			.O(gen[3366]),
			.E(gen[3368]),

			.SO(gen[3461]),
			.S(gen[3462]),
			.SE(gen[3463]),

			.SELF(gen[3367]),
			.cell_state(gen[3367])
		); 

/******************* CELL 3368 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3368 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3272]),
			.N(gen[3273]),
			.NE(gen[3274]),

			.O(gen[3367]),
			.E(gen[3369]),

			.SO(gen[3462]),
			.S(gen[3463]),
			.SE(gen[3464]),

			.SELF(gen[3368]),
			.cell_state(gen[3368])
		); 

/******************* CELL 3369 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3369 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3273]),
			.N(gen[3274]),
			.NE(gen[3275]),

			.O(gen[3368]),
			.E(gen[3370]),

			.SO(gen[3463]),
			.S(gen[3464]),
			.SE(gen[3465]),

			.SELF(gen[3369]),
			.cell_state(gen[3369])
		); 

/******************* CELL 3370 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3370 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3274]),
			.N(gen[3275]),
			.NE(gen[3276]),

			.O(gen[3369]),
			.E(gen[3371]),

			.SO(gen[3464]),
			.S(gen[3465]),
			.SE(gen[3466]),

			.SELF(gen[3370]),
			.cell_state(gen[3370])
		); 

/******************* CELL 3371 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3371 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3275]),
			.N(gen[3276]),
			.NE(gen[3277]),

			.O(gen[3370]),
			.E(gen[3372]),

			.SO(gen[3465]),
			.S(gen[3466]),
			.SE(gen[3467]),

			.SELF(gen[3371]),
			.cell_state(gen[3371])
		); 

/******************* CELL 3372 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3372 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3276]),
			.N(gen[3277]),
			.NE(gen[3278]),

			.O(gen[3371]),
			.E(gen[3373]),

			.SO(gen[3466]),
			.S(gen[3467]),
			.SE(gen[3468]),

			.SELF(gen[3372]),
			.cell_state(gen[3372])
		); 

/******************* CELL 3373 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3373 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3277]),
			.N(gen[3278]),
			.NE(gen[3279]),

			.O(gen[3372]),
			.E(gen[3374]),

			.SO(gen[3467]),
			.S(gen[3468]),
			.SE(gen[3469]),

			.SELF(gen[3373]),
			.cell_state(gen[3373])
		); 

/******************* CELL 3374 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3374 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3278]),
			.N(gen[3279]),
			.NE(gen[3280]),

			.O(gen[3373]),
			.E(gen[3375]),

			.SO(gen[3468]),
			.S(gen[3469]),
			.SE(gen[3470]),

			.SELF(gen[3374]),
			.cell_state(gen[3374])
		); 

/******************* CELL 3375 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3375 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3279]),
			.N(gen[3280]),
			.NE(gen[3281]),

			.O(gen[3374]),
			.E(gen[3376]),

			.SO(gen[3469]),
			.S(gen[3470]),
			.SE(gen[3471]),

			.SELF(gen[3375]),
			.cell_state(gen[3375])
		); 

/******************* CELL 3376 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3376 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3280]),
			.N(gen[3281]),
			.NE(gen[3282]),

			.O(gen[3375]),
			.E(gen[3377]),

			.SO(gen[3470]),
			.S(gen[3471]),
			.SE(gen[3472]),

			.SELF(gen[3376]),
			.cell_state(gen[3376])
		); 

/******************* CELL 3377 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3377 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3281]),
			.N(gen[3282]),
			.NE(gen[3283]),

			.O(gen[3376]),
			.E(gen[3378]),

			.SO(gen[3471]),
			.S(gen[3472]),
			.SE(gen[3473]),

			.SELF(gen[3377]),
			.cell_state(gen[3377])
		); 

/******************* CELL 3378 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3378 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3282]),
			.N(gen[3283]),
			.NE(gen[3284]),

			.O(gen[3377]),
			.E(gen[3379]),

			.SO(gen[3472]),
			.S(gen[3473]),
			.SE(gen[3474]),

			.SELF(gen[3378]),
			.cell_state(gen[3378])
		); 

/******************* CELL 3379 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3379 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3283]),
			.N(gen[3284]),
			.NE(gen[3285]),

			.O(gen[3378]),
			.E(gen[3380]),

			.SO(gen[3473]),
			.S(gen[3474]),
			.SE(gen[3475]),

			.SELF(gen[3379]),
			.cell_state(gen[3379])
		); 

/******************* CELL 3380 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3380 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3284]),
			.N(gen[3285]),
			.NE(gen[3286]),

			.O(gen[3379]),
			.E(gen[3381]),

			.SO(gen[3474]),
			.S(gen[3475]),
			.SE(gen[3476]),

			.SELF(gen[3380]),
			.cell_state(gen[3380])
		); 

/******************* CELL 3381 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3381 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3285]),
			.N(gen[3286]),
			.NE(gen[3287]),

			.O(gen[3380]),
			.E(gen[3382]),

			.SO(gen[3475]),
			.S(gen[3476]),
			.SE(gen[3477]),

			.SELF(gen[3381]),
			.cell_state(gen[3381])
		); 

/******************* CELL 3382 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3382 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3286]),
			.N(gen[3287]),
			.NE(gen[3288]),

			.O(gen[3381]),
			.E(gen[3383]),

			.SO(gen[3476]),
			.S(gen[3477]),
			.SE(gen[3478]),

			.SELF(gen[3382]),
			.cell_state(gen[3382])
		); 

/******************* CELL 3383 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3383 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3287]),
			.N(gen[3288]),
			.NE(gen[3289]),

			.O(gen[3382]),
			.E(gen[3384]),

			.SO(gen[3477]),
			.S(gen[3478]),
			.SE(gen[3479]),

			.SELF(gen[3383]),
			.cell_state(gen[3383])
		); 

/******************* CELL 3384 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3384 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3288]),
			.N(gen[3289]),
			.NE(gen[3290]),

			.O(gen[3383]),
			.E(gen[3385]),

			.SO(gen[3478]),
			.S(gen[3479]),
			.SE(gen[3480]),

			.SELF(gen[3384]),
			.cell_state(gen[3384])
		); 

/******************* CELL 3385 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3385 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3289]),
			.N(gen[3290]),
			.NE(gen[3291]),

			.O(gen[3384]),
			.E(gen[3386]),

			.SO(gen[3479]),
			.S(gen[3480]),
			.SE(gen[3481]),

			.SELF(gen[3385]),
			.cell_state(gen[3385])
		); 

/******************* CELL 3386 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3386 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3290]),
			.N(gen[3291]),
			.NE(gen[3292]),

			.O(gen[3385]),
			.E(gen[3387]),

			.SO(gen[3480]),
			.S(gen[3481]),
			.SE(gen[3482]),

			.SELF(gen[3386]),
			.cell_state(gen[3386])
		); 

/******************* CELL 3387 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3387 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3291]),
			.N(gen[3292]),
			.NE(gen[3293]),

			.O(gen[3386]),
			.E(gen[3388]),

			.SO(gen[3481]),
			.S(gen[3482]),
			.SE(gen[3483]),

			.SELF(gen[3387]),
			.cell_state(gen[3387])
		); 

/******************* CELL 3388 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3388 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3292]),
			.N(gen[3293]),
			.NE(gen[3294]),

			.O(gen[3387]),
			.E(gen[3389]),

			.SO(gen[3482]),
			.S(gen[3483]),
			.SE(gen[3484]),

			.SELF(gen[3388]),
			.cell_state(gen[3388])
		); 

/******************* CELL 3389 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3389 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3293]),
			.N(gen[3294]),
			.NE(gen[3295]),

			.O(gen[3388]),
			.E(gen[3390]),

			.SO(gen[3483]),
			.S(gen[3484]),
			.SE(gen[3485]),

			.SELF(gen[3389]),
			.cell_state(gen[3389])
		); 

/******************* CELL 3390 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3390 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3294]),
			.N(gen[3295]),
			.NE(gen[3296]),

			.O(gen[3389]),
			.E(gen[3391]),

			.SO(gen[3484]),
			.S(gen[3485]),
			.SE(gen[3486]),

			.SELF(gen[3390]),
			.cell_state(gen[3390])
		); 

/******************* CELL 3391 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3391 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3295]),
			.N(gen[3296]),
			.NE(gen[3297]),

			.O(gen[3390]),
			.E(gen[3392]),

			.SO(gen[3485]),
			.S(gen[3486]),
			.SE(gen[3487]),

			.SELF(gen[3391]),
			.cell_state(gen[3391])
		); 

/******************* CELL 3392 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3392 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3296]),
			.N(gen[3297]),
			.NE(gen[3298]),

			.O(gen[3391]),
			.E(gen[3393]),

			.SO(gen[3486]),
			.S(gen[3487]),
			.SE(gen[3488]),

			.SELF(gen[3392]),
			.cell_state(gen[3392])
		); 

/******************* CELL 3393 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3393 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3297]),
			.N(gen[3298]),
			.NE(gen[3299]),

			.O(gen[3392]),
			.E(gen[3394]),

			.SO(gen[3487]),
			.S(gen[3488]),
			.SE(gen[3489]),

			.SELF(gen[3393]),
			.cell_state(gen[3393])
		); 

/******************* CELL 3394 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3394 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3298]),
			.N(gen[3299]),
			.NE(gen[3300]),

			.O(gen[3393]),
			.E(gen[3395]),

			.SO(gen[3488]),
			.S(gen[3489]),
			.SE(gen[3490]),

			.SELF(gen[3394]),
			.cell_state(gen[3394])
		); 

/******************* CELL 3395 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3395 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3299]),
			.N(gen[3300]),
			.NE(gen[3301]),

			.O(gen[3394]),
			.E(gen[3396]),

			.SO(gen[3489]),
			.S(gen[3490]),
			.SE(gen[3491]),

			.SELF(gen[3395]),
			.cell_state(gen[3395])
		); 

/******************* CELL 3396 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3396 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3300]),
			.N(gen[3301]),
			.NE(gen[3302]),

			.O(gen[3395]),
			.E(gen[3397]),

			.SO(gen[3490]),
			.S(gen[3491]),
			.SE(gen[3492]),

			.SELF(gen[3396]),
			.cell_state(gen[3396])
		); 

/******************* CELL 3397 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3397 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3301]),
			.N(gen[3302]),
			.NE(gen[3303]),

			.O(gen[3396]),
			.E(gen[3398]),

			.SO(gen[3491]),
			.S(gen[3492]),
			.SE(gen[3493]),

			.SELF(gen[3397]),
			.cell_state(gen[3397])
		); 

/******************* CELL 3398 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3398 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3302]),
			.N(gen[3303]),
			.NE(gen[3304]),

			.O(gen[3397]),
			.E(gen[3399]),

			.SO(gen[3492]),
			.S(gen[3493]),
			.SE(gen[3494]),

			.SELF(gen[3398]),
			.cell_state(gen[3398])
		); 

/******************* CELL 3399 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3399 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3303]),
			.N(gen[3304]),
			.NE(gen[3305]),

			.O(gen[3398]),
			.E(gen[3400]),

			.SO(gen[3493]),
			.S(gen[3494]),
			.SE(gen[3495]),

			.SELF(gen[3399]),
			.cell_state(gen[3399])
		); 

/******************* CELL 3400 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3400 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3304]),
			.N(gen[3305]),
			.NE(gen[3306]),

			.O(gen[3399]),
			.E(gen[3401]),

			.SO(gen[3494]),
			.S(gen[3495]),
			.SE(gen[3496]),

			.SELF(gen[3400]),
			.cell_state(gen[3400])
		); 

/******************* CELL 3401 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3401 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3305]),
			.N(gen[3306]),
			.NE(gen[3307]),

			.O(gen[3400]),
			.E(gen[3402]),

			.SO(gen[3495]),
			.S(gen[3496]),
			.SE(gen[3497]),

			.SELF(gen[3401]),
			.cell_state(gen[3401])
		); 

/******************* CELL 3402 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3402 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3306]),
			.N(gen[3307]),
			.NE(gen[3308]),

			.O(gen[3401]),
			.E(gen[3403]),

			.SO(gen[3496]),
			.S(gen[3497]),
			.SE(gen[3498]),

			.SELF(gen[3402]),
			.cell_state(gen[3402])
		); 

/******************* CELL 3403 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3403 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3307]),
			.N(gen[3308]),
			.NE(gen[3309]),

			.O(gen[3402]),
			.E(gen[3404]),

			.SO(gen[3497]),
			.S(gen[3498]),
			.SE(gen[3499]),

			.SELF(gen[3403]),
			.cell_state(gen[3403])
		); 

/******************* CELL 3404 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3404 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3308]),
			.N(gen[3309]),
			.NE(gen[3310]),

			.O(gen[3403]),
			.E(gen[3405]),

			.SO(gen[3498]),
			.S(gen[3499]),
			.SE(gen[3500]),

			.SELF(gen[3404]),
			.cell_state(gen[3404])
		); 

/******************* CELL 3405 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3405 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3309]),
			.N(gen[3310]),
			.NE(gen[3311]),

			.O(gen[3404]),
			.E(gen[3406]),

			.SO(gen[3499]),
			.S(gen[3500]),
			.SE(gen[3501]),

			.SELF(gen[3405]),
			.cell_state(gen[3405])
		); 

/******************* CELL 3406 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3406 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3310]),
			.N(gen[3311]),
			.NE(gen[3312]),

			.O(gen[3405]),
			.E(gen[3407]),

			.SO(gen[3500]),
			.S(gen[3501]),
			.SE(gen[3502]),

			.SELF(gen[3406]),
			.cell_state(gen[3406])
		); 

/******************* CELL 3407 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3407 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3311]),
			.N(gen[3312]),
			.NE(gen[3313]),

			.O(gen[3406]),
			.E(gen[3408]),

			.SO(gen[3501]),
			.S(gen[3502]),
			.SE(gen[3503]),

			.SELF(gen[3407]),
			.cell_state(gen[3407])
		); 

/******************* CELL 3408 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3408 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3312]),
			.N(gen[3313]),
			.NE(gen[3314]),

			.O(gen[3407]),
			.E(gen[3409]),

			.SO(gen[3502]),
			.S(gen[3503]),
			.SE(gen[3504]),

			.SELF(gen[3408]),
			.cell_state(gen[3408])
		); 

/******************* CELL 3409 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3409 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3313]),
			.N(gen[3314]),
			.NE(gen[3315]),

			.O(gen[3408]),
			.E(gen[3410]),

			.SO(gen[3503]),
			.S(gen[3504]),
			.SE(gen[3505]),

			.SELF(gen[3409]),
			.cell_state(gen[3409])
		); 

/******************* CELL 3410 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3410 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3314]),
			.N(gen[3315]),
			.NE(gen[3316]),

			.O(gen[3409]),
			.E(gen[3411]),

			.SO(gen[3504]),
			.S(gen[3505]),
			.SE(gen[3506]),

			.SELF(gen[3410]),
			.cell_state(gen[3410])
		); 

/******************* CELL 3411 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3411 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3315]),
			.N(gen[3316]),
			.NE(gen[3317]),

			.O(gen[3410]),
			.E(gen[3412]),

			.SO(gen[3505]),
			.S(gen[3506]),
			.SE(gen[3507]),

			.SELF(gen[3411]),
			.cell_state(gen[3411])
		); 

/******************* CELL 3412 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3412 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3316]),
			.N(gen[3317]),
			.NE(gen[3318]),

			.O(gen[3411]),
			.E(gen[3413]),

			.SO(gen[3506]),
			.S(gen[3507]),
			.SE(gen[3508]),

			.SELF(gen[3412]),
			.cell_state(gen[3412])
		); 

/******************* CELL 3413 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3413 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3317]),
			.N(gen[3318]),
			.NE(gen[3319]),

			.O(gen[3412]),
			.E(gen[3414]),

			.SO(gen[3507]),
			.S(gen[3508]),
			.SE(gen[3509]),

			.SELF(gen[3413]),
			.cell_state(gen[3413])
		); 

/******************* CELL 3414 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3414 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3318]),
			.N(gen[3319]),
			.NE(gen[3320]),

			.O(gen[3413]),
			.E(gen[3415]),

			.SO(gen[3508]),
			.S(gen[3509]),
			.SE(gen[3510]),

			.SELF(gen[3414]),
			.cell_state(gen[3414])
		); 

/******************* CELL 3415 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3415 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3319]),
			.N(gen[3320]),
			.NE(gen[3321]),

			.O(gen[3414]),
			.E(gen[3416]),

			.SO(gen[3509]),
			.S(gen[3510]),
			.SE(gen[3511]),

			.SELF(gen[3415]),
			.cell_state(gen[3415])
		); 

/******************* CELL 3416 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3416 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3320]),
			.N(gen[3321]),
			.NE(gen[3322]),

			.O(gen[3415]),
			.E(gen[3417]),

			.SO(gen[3510]),
			.S(gen[3511]),
			.SE(gen[3512]),

			.SELF(gen[3416]),
			.cell_state(gen[3416])
		); 

/******************* CELL 3417 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3417 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3321]),
			.N(gen[3322]),
			.NE(gen[3323]),

			.O(gen[3416]),
			.E(gen[3418]),

			.SO(gen[3511]),
			.S(gen[3512]),
			.SE(gen[3513]),

			.SELF(gen[3417]),
			.cell_state(gen[3417])
		); 

/******************* CELL 3418 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3418 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3322]),
			.N(gen[3323]),
			.NE(gen[3324]),

			.O(gen[3417]),
			.E(gen[3419]),

			.SO(gen[3512]),
			.S(gen[3513]),
			.SE(gen[3514]),

			.SELF(gen[3418]),
			.cell_state(gen[3418])
		); 

/******************* CELL 3419 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3419 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3323]),
			.N(gen[3324]),
			.NE(gen[3323]),

			.O(gen[3418]),
			.E(gen[3418]),

			.SO(gen[3513]),
			.S(gen[3514]),
			.SE(gen[3513]),

			.SELF(gen[3419]),
			.cell_state(gen[3419])
		); 

/******************* CELL 3420 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3420 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3326]),
			.N(gen[3325]),
			.NE(gen[3326]),

			.O(gen[3421]),
			.E(gen[3421]),

			.SO(gen[3516]),
			.S(gen[3515]),
			.SE(gen[3516]),

			.SELF(gen[3420]),
			.cell_state(gen[3420])
		); 

/******************* CELL 3421 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3421 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3325]),
			.N(gen[3326]),
			.NE(gen[3327]),

			.O(gen[3420]),
			.E(gen[3422]),

			.SO(gen[3515]),
			.S(gen[3516]),
			.SE(gen[3517]),

			.SELF(gen[3421]),
			.cell_state(gen[3421])
		); 

/******************* CELL 3422 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3422 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3326]),
			.N(gen[3327]),
			.NE(gen[3328]),

			.O(gen[3421]),
			.E(gen[3423]),

			.SO(gen[3516]),
			.S(gen[3517]),
			.SE(gen[3518]),

			.SELF(gen[3422]),
			.cell_state(gen[3422])
		); 

/******************* CELL 3423 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3423 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3327]),
			.N(gen[3328]),
			.NE(gen[3329]),

			.O(gen[3422]),
			.E(gen[3424]),

			.SO(gen[3517]),
			.S(gen[3518]),
			.SE(gen[3519]),

			.SELF(gen[3423]),
			.cell_state(gen[3423])
		); 

/******************* CELL 3424 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3424 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3328]),
			.N(gen[3329]),
			.NE(gen[3330]),

			.O(gen[3423]),
			.E(gen[3425]),

			.SO(gen[3518]),
			.S(gen[3519]),
			.SE(gen[3520]),

			.SELF(gen[3424]),
			.cell_state(gen[3424])
		); 

/******************* CELL 3425 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3425 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3329]),
			.N(gen[3330]),
			.NE(gen[3331]),

			.O(gen[3424]),
			.E(gen[3426]),

			.SO(gen[3519]),
			.S(gen[3520]),
			.SE(gen[3521]),

			.SELF(gen[3425]),
			.cell_state(gen[3425])
		); 

/******************* CELL 3426 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3426 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3330]),
			.N(gen[3331]),
			.NE(gen[3332]),

			.O(gen[3425]),
			.E(gen[3427]),

			.SO(gen[3520]),
			.S(gen[3521]),
			.SE(gen[3522]),

			.SELF(gen[3426]),
			.cell_state(gen[3426])
		); 

/******************* CELL 3427 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3427 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3331]),
			.N(gen[3332]),
			.NE(gen[3333]),

			.O(gen[3426]),
			.E(gen[3428]),

			.SO(gen[3521]),
			.S(gen[3522]),
			.SE(gen[3523]),

			.SELF(gen[3427]),
			.cell_state(gen[3427])
		); 

/******************* CELL 3428 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3428 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3332]),
			.N(gen[3333]),
			.NE(gen[3334]),

			.O(gen[3427]),
			.E(gen[3429]),

			.SO(gen[3522]),
			.S(gen[3523]),
			.SE(gen[3524]),

			.SELF(gen[3428]),
			.cell_state(gen[3428])
		); 

/******************* CELL 3429 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3429 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3333]),
			.N(gen[3334]),
			.NE(gen[3335]),

			.O(gen[3428]),
			.E(gen[3430]),

			.SO(gen[3523]),
			.S(gen[3524]),
			.SE(gen[3525]),

			.SELF(gen[3429]),
			.cell_state(gen[3429])
		); 

/******************* CELL 3430 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3430 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3334]),
			.N(gen[3335]),
			.NE(gen[3336]),

			.O(gen[3429]),
			.E(gen[3431]),

			.SO(gen[3524]),
			.S(gen[3525]),
			.SE(gen[3526]),

			.SELF(gen[3430]),
			.cell_state(gen[3430])
		); 

/******************* CELL 3431 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3431 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3335]),
			.N(gen[3336]),
			.NE(gen[3337]),

			.O(gen[3430]),
			.E(gen[3432]),

			.SO(gen[3525]),
			.S(gen[3526]),
			.SE(gen[3527]),

			.SELF(gen[3431]),
			.cell_state(gen[3431])
		); 

/******************* CELL 3432 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3432 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3336]),
			.N(gen[3337]),
			.NE(gen[3338]),

			.O(gen[3431]),
			.E(gen[3433]),

			.SO(gen[3526]),
			.S(gen[3527]),
			.SE(gen[3528]),

			.SELF(gen[3432]),
			.cell_state(gen[3432])
		); 

/******************* CELL 3433 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3433 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3337]),
			.N(gen[3338]),
			.NE(gen[3339]),

			.O(gen[3432]),
			.E(gen[3434]),

			.SO(gen[3527]),
			.S(gen[3528]),
			.SE(gen[3529]),

			.SELF(gen[3433]),
			.cell_state(gen[3433])
		); 

/******************* CELL 3434 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3434 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3338]),
			.N(gen[3339]),
			.NE(gen[3340]),

			.O(gen[3433]),
			.E(gen[3435]),

			.SO(gen[3528]),
			.S(gen[3529]),
			.SE(gen[3530]),

			.SELF(gen[3434]),
			.cell_state(gen[3434])
		); 

/******************* CELL 3435 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3435 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3339]),
			.N(gen[3340]),
			.NE(gen[3341]),

			.O(gen[3434]),
			.E(gen[3436]),

			.SO(gen[3529]),
			.S(gen[3530]),
			.SE(gen[3531]),

			.SELF(gen[3435]),
			.cell_state(gen[3435])
		); 

/******************* CELL 3436 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3436 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3340]),
			.N(gen[3341]),
			.NE(gen[3342]),

			.O(gen[3435]),
			.E(gen[3437]),

			.SO(gen[3530]),
			.S(gen[3531]),
			.SE(gen[3532]),

			.SELF(gen[3436]),
			.cell_state(gen[3436])
		); 

/******************* CELL 3437 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3437 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3341]),
			.N(gen[3342]),
			.NE(gen[3343]),

			.O(gen[3436]),
			.E(gen[3438]),

			.SO(gen[3531]),
			.S(gen[3532]),
			.SE(gen[3533]),

			.SELF(gen[3437]),
			.cell_state(gen[3437])
		); 

/******************* CELL 3438 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3438 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3342]),
			.N(gen[3343]),
			.NE(gen[3344]),

			.O(gen[3437]),
			.E(gen[3439]),

			.SO(gen[3532]),
			.S(gen[3533]),
			.SE(gen[3534]),

			.SELF(gen[3438]),
			.cell_state(gen[3438])
		); 

/******************* CELL 3439 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3439 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3343]),
			.N(gen[3344]),
			.NE(gen[3345]),

			.O(gen[3438]),
			.E(gen[3440]),

			.SO(gen[3533]),
			.S(gen[3534]),
			.SE(gen[3535]),

			.SELF(gen[3439]),
			.cell_state(gen[3439])
		); 

/******************* CELL 3440 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3440 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3344]),
			.N(gen[3345]),
			.NE(gen[3346]),

			.O(gen[3439]),
			.E(gen[3441]),

			.SO(gen[3534]),
			.S(gen[3535]),
			.SE(gen[3536]),

			.SELF(gen[3440]),
			.cell_state(gen[3440])
		); 

/******************* CELL 3441 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3441 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3345]),
			.N(gen[3346]),
			.NE(gen[3347]),

			.O(gen[3440]),
			.E(gen[3442]),

			.SO(gen[3535]),
			.S(gen[3536]),
			.SE(gen[3537]),

			.SELF(gen[3441]),
			.cell_state(gen[3441])
		); 

/******************* CELL 3442 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3442 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3346]),
			.N(gen[3347]),
			.NE(gen[3348]),

			.O(gen[3441]),
			.E(gen[3443]),

			.SO(gen[3536]),
			.S(gen[3537]),
			.SE(gen[3538]),

			.SELF(gen[3442]),
			.cell_state(gen[3442])
		); 

/******************* CELL 3443 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3443 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3347]),
			.N(gen[3348]),
			.NE(gen[3349]),

			.O(gen[3442]),
			.E(gen[3444]),

			.SO(gen[3537]),
			.S(gen[3538]),
			.SE(gen[3539]),

			.SELF(gen[3443]),
			.cell_state(gen[3443])
		); 

/******************* CELL 3444 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3444 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3348]),
			.N(gen[3349]),
			.NE(gen[3350]),

			.O(gen[3443]),
			.E(gen[3445]),

			.SO(gen[3538]),
			.S(gen[3539]),
			.SE(gen[3540]),

			.SELF(gen[3444]),
			.cell_state(gen[3444])
		); 

/******************* CELL 3445 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3445 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3349]),
			.N(gen[3350]),
			.NE(gen[3351]),

			.O(gen[3444]),
			.E(gen[3446]),

			.SO(gen[3539]),
			.S(gen[3540]),
			.SE(gen[3541]),

			.SELF(gen[3445]),
			.cell_state(gen[3445])
		); 

/******************* CELL 3446 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3446 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3350]),
			.N(gen[3351]),
			.NE(gen[3352]),

			.O(gen[3445]),
			.E(gen[3447]),

			.SO(gen[3540]),
			.S(gen[3541]),
			.SE(gen[3542]),

			.SELF(gen[3446]),
			.cell_state(gen[3446])
		); 

/******************* CELL 3447 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3447 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3351]),
			.N(gen[3352]),
			.NE(gen[3353]),

			.O(gen[3446]),
			.E(gen[3448]),

			.SO(gen[3541]),
			.S(gen[3542]),
			.SE(gen[3543]),

			.SELF(gen[3447]),
			.cell_state(gen[3447])
		); 

/******************* CELL 3448 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3448 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3352]),
			.N(gen[3353]),
			.NE(gen[3354]),

			.O(gen[3447]),
			.E(gen[3449]),

			.SO(gen[3542]),
			.S(gen[3543]),
			.SE(gen[3544]),

			.SELF(gen[3448]),
			.cell_state(gen[3448])
		); 

/******************* CELL 3449 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3449 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3353]),
			.N(gen[3354]),
			.NE(gen[3355]),

			.O(gen[3448]),
			.E(gen[3450]),

			.SO(gen[3543]),
			.S(gen[3544]),
			.SE(gen[3545]),

			.SELF(gen[3449]),
			.cell_state(gen[3449])
		); 

/******************* CELL 3450 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3450 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3354]),
			.N(gen[3355]),
			.NE(gen[3356]),

			.O(gen[3449]),
			.E(gen[3451]),

			.SO(gen[3544]),
			.S(gen[3545]),
			.SE(gen[3546]),

			.SELF(gen[3450]),
			.cell_state(gen[3450])
		); 

/******************* CELL 3451 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3451 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3355]),
			.N(gen[3356]),
			.NE(gen[3357]),

			.O(gen[3450]),
			.E(gen[3452]),

			.SO(gen[3545]),
			.S(gen[3546]),
			.SE(gen[3547]),

			.SELF(gen[3451]),
			.cell_state(gen[3451])
		); 

/******************* CELL 3452 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3452 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3356]),
			.N(gen[3357]),
			.NE(gen[3358]),

			.O(gen[3451]),
			.E(gen[3453]),

			.SO(gen[3546]),
			.S(gen[3547]),
			.SE(gen[3548]),

			.SELF(gen[3452]),
			.cell_state(gen[3452])
		); 

/******************* CELL 3453 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3453 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3357]),
			.N(gen[3358]),
			.NE(gen[3359]),

			.O(gen[3452]),
			.E(gen[3454]),

			.SO(gen[3547]),
			.S(gen[3548]),
			.SE(gen[3549]),

			.SELF(gen[3453]),
			.cell_state(gen[3453])
		); 

/******************* CELL 3454 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3454 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3358]),
			.N(gen[3359]),
			.NE(gen[3360]),

			.O(gen[3453]),
			.E(gen[3455]),

			.SO(gen[3548]),
			.S(gen[3549]),
			.SE(gen[3550]),

			.SELF(gen[3454]),
			.cell_state(gen[3454])
		); 

/******************* CELL 3455 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3455 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3359]),
			.N(gen[3360]),
			.NE(gen[3361]),

			.O(gen[3454]),
			.E(gen[3456]),

			.SO(gen[3549]),
			.S(gen[3550]),
			.SE(gen[3551]),

			.SELF(gen[3455]),
			.cell_state(gen[3455])
		); 

/******************* CELL 3456 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3456 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3360]),
			.N(gen[3361]),
			.NE(gen[3362]),

			.O(gen[3455]),
			.E(gen[3457]),

			.SO(gen[3550]),
			.S(gen[3551]),
			.SE(gen[3552]),

			.SELF(gen[3456]),
			.cell_state(gen[3456])
		); 

/******************* CELL 3457 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3457 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3361]),
			.N(gen[3362]),
			.NE(gen[3363]),

			.O(gen[3456]),
			.E(gen[3458]),

			.SO(gen[3551]),
			.S(gen[3552]),
			.SE(gen[3553]),

			.SELF(gen[3457]),
			.cell_state(gen[3457])
		); 

/******************* CELL 3458 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3458 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3362]),
			.N(gen[3363]),
			.NE(gen[3364]),

			.O(gen[3457]),
			.E(gen[3459]),

			.SO(gen[3552]),
			.S(gen[3553]),
			.SE(gen[3554]),

			.SELF(gen[3458]),
			.cell_state(gen[3458])
		); 

/******************* CELL 3459 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3459 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3363]),
			.N(gen[3364]),
			.NE(gen[3365]),

			.O(gen[3458]),
			.E(gen[3460]),

			.SO(gen[3553]),
			.S(gen[3554]),
			.SE(gen[3555]),

			.SELF(gen[3459]),
			.cell_state(gen[3459])
		); 

/******************* CELL 3460 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3460 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3364]),
			.N(gen[3365]),
			.NE(gen[3366]),

			.O(gen[3459]),
			.E(gen[3461]),

			.SO(gen[3554]),
			.S(gen[3555]),
			.SE(gen[3556]),

			.SELF(gen[3460]),
			.cell_state(gen[3460])
		); 

/******************* CELL 3461 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3461 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3365]),
			.N(gen[3366]),
			.NE(gen[3367]),

			.O(gen[3460]),
			.E(gen[3462]),

			.SO(gen[3555]),
			.S(gen[3556]),
			.SE(gen[3557]),

			.SELF(gen[3461]),
			.cell_state(gen[3461])
		); 

/******************* CELL 3462 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3462 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3366]),
			.N(gen[3367]),
			.NE(gen[3368]),

			.O(gen[3461]),
			.E(gen[3463]),

			.SO(gen[3556]),
			.S(gen[3557]),
			.SE(gen[3558]),

			.SELF(gen[3462]),
			.cell_state(gen[3462])
		); 

/******************* CELL 3463 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3463 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3367]),
			.N(gen[3368]),
			.NE(gen[3369]),

			.O(gen[3462]),
			.E(gen[3464]),

			.SO(gen[3557]),
			.S(gen[3558]),
			.SE(gen[3559]),

			.SELF(gen[3463]),
			.cell_state(gen[3463])
		); 

/******************* CELL 3464 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3464 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3368]),
			.N(gen[3369]),
			.NE(gen[3370]),

			.O(gen[3463]),
			.E(gen[3465]),

			.SO(gen[3558]),
			.S(gen[3559]),
			.SE(gen[3560]),

			.SELF(gen[3464]),
			.cell_state(gen[3464])
		); 

/******************* CELL 3465 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3465 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3369]),
			.N(gen[3370]),
			.NE(gen[3371]),

			.O(gen[3464]),
			.E(gen[3466]),

			.SO(gen[3559]),
			.S(gen[3560]),
			.SE(gen[3561]),

			.SELF(gen[3465]),
			.cell_state(gen[3465])
		); 

/******************* CELL 3466 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3466 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3370]),
			.N(gen[3371]),
			.NE(gen[3372]),

			.O(gen[3465]),
			.E(gen[3467]),

			.SO(gen[3560]),
			.S(gen[3561]),
			.SE(gen[3562]),

			.SELF(gen[3466]),
			.cell_state(gen[3466])
		); 

/******************* CELL 3467 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3467 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3371]),
			.N(gen[3372]),
			.NE(gen[3373]),

			.O(gen[3466]),
			.E(gen[3468]),

			.SO(gen[3561]),
			.S(gen[3562]),
			.SE(gen[3563]),

			.SELF(gen[3467]),
			.cell_state(gen[3467])
		); 

/******************* CELL 3468 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3468 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3372]),
			.N(gen[3373]),
			.NE(gen[3374]),

			.O(gen[3467]),
			.E(gen[3469]),

			.SO(gen[3562]),
			.S(gen[3563]),
			.SE(gen[3564]),

			.SELF(gen[3468]),
			.cell_state(gen[3468])
		); 

/******************* CELL 3469 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3469 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3373]),
			.N(gen[3374]),
			.NE(gen[3375]),

			.O(gen[3468]),
			.E(gen[3470]),

			.SO(gen[3563]),
			.S(gen[3564]),
			.SE(gen[3565]),

			.SELF(gen[3469]),
			.cell_state(gen[3469])
		); 

/******************* CELL 3470 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3470 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3374]),
			.N(gen[3375]),
			.NE(gen[3376]),

			.O(gen[3469]),
			.E(gen[3471]),

			.SO(gen[3564]),
			.S(gen[3565]),
			.SE(gen[3566]),

			.SELF(gen[3470]),
			.cell_state(gen[3470])
		); 

/******************* CELL 3471 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3471 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3375]),
			.N(gen[3376]),
			.NE(gen[3377]),

			.O(gen[3470]),
			.E(gen[3472]),

			.SO(gen[3565]),
			.S(gen[3566]),
			.SE(gen[3567]),

			.SELF(gen[3471]),
			.cell_state(gen[3471])
		); 

/******************* CELL 3472 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3472 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3376]),
			.N(gen[3377]),
			.NE(gen[3378]),

			.O(gen[3471]),
			.E(gen[3473]),

			.SO(gen[3566]),
			.S(gen[3567]),
			.SE(gen[3568]),

			.SELF(gen[3472]),
			.cell_state(gen[3472])
		); 

/******************* CELL 3473 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3473 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3377]),
			.N(gen[3378]),
			.NE(gen[3379]),

			.O(gen[3472]),
			.E(gen[3474]),

			.SO(gen[3567]),
			.S(gen[3568]),
			.SE(gen[3569]),

			.SELF(gen[3473]),
			.cell_state(gen[3473])
		); 

/******************* CELL 3474 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3474 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3378]),
			.N(gen[3379]),
			.NE(gen[3380]),

			.O(gen[3473]),
			.E(gen[3475]),

			.SO(gen[3568]),
			.S(gen[3569]),
			.SE(gen[3570]),

			.SELF(gen[3474]),
			.cell_state(gen[3474])
		); 

/******************* CELL 3475 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3475 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3379]),
			.N(gen[3380]),
			.NE(gen[3381]),

			.O(gen[3474]),
			.E(gen[3476]),

			.SO(gen[3569]),
			.S(gen[3570]),
			.SE(gen[3571]),

			.SELF(gen[3475]),
			.cell_state(gen[3475])
		); 

/******************* CELL 3476 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3476 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3380]),
			.N(gen[3381]),
			.NE(gen[3382]),

			.O(gen[3475]),
			.E(gen[3477]),

			.SO(gen[3570]),
			.S(gen[3571]),
			.SE(gen[3572]),

			.SELF(gen[3476]),
			.cell_state(gen[3476])
		); 

/******************* CELL 3477 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3477 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3381]),
			.N(gen[3382]),
			.NE(gen[3383]),

			.O(gen[3476]),
			.E(gen[3478]),

			.SO(gen[3571]),
			.S(gen[3572]),
			.SE(gen[3573]),

			.SELF(gen[3477]),
			.cell_state(gen[3477])
		); 

/******************* CELL 3478 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3478 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3382]),
			.N(gen[3383]),
			.NE(gen[3384]),

			.O(gen[3477]),
			.E(gen[3479]),

			.SO(gen[3572]),
			.S(gen[3573]),
			.SE(gen[3574]),

			.SELF(gen[3478]),
			.cell_state(gen[3478])
		); 

/******************* CELL 3479 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3479 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3383]),
			.N(gen[3384]),
			.NE(gen[3385]),

			.O(gen[3478]),
			.E(gen[3480]),

			.SO(gen[3573]),
			.S(gen[3574]),
			.SE(gen[3575]),

			.SELF(gen[3479]),
			.cell_state(gen[3479])
		); 

/******************* CELL 3480 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3480 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3384]),
			.N(gen[3385]),
			.NE(gen[3386]),

			.O(gen[3479]),
			.E(gen[3481]),

			.SO(gen[3574]),
			.S(gen[3575]),
			.SE(gen[3576]),

			.SELF(gen[3480]),
			.cell_state(gen[3480])
		); 

/******************* CELL 3481 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3481 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3385]),
			.N(gen[3386]),
			.NE(gen[3387]),

			.O(gen[3480]),
			.E(gen[3482]),

			.SO(gen[3575]),
			.S(gen[3576]),
			.SE(gen[3577]),

			.SELF(gen[3481]),
			.cell_state(gen[3481])
		); 

/******************* CELL 3482 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3482 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3386]),
			.N(gen[3387]),
			.NE(gen[3388]),

			.O(gen[3481]),
			.E(gen[3483]),

			.SO(gen[3576]),
			.S(gen[3577]),
			.SE(gen[3578]),

			.SELF(gen[3482]),
			.cell_state(gen[3482])
		); 

/******************* CELL 3483 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3483 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3387]),
			.N(gen[3388]),
			.NE(gen[3389]),

			.O(gen[3482]),
			.E(gen[3484]),

			.SO(gen[3577]),
			.S(gen[3578]),
			.SE(gen[3579]),

			.SELF(gen[3483]),
			.cell_state(gen[3483])
		); 

/******************* CELL 3484 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3484 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3388]),
			.N(gen[3389]),
			.NE(gen[3390]),

			.O(gen[3483]),
			.E(gen[3485]),

			.SO(gen[3578]),
			.S(gen[3579]),
			.SE(gen[3580]),

			.SELF(gen[3484]),
			.cell_state(gen[3484])
		); 

/******************* CELL 3485 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3485 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3389]),
			.N(gen[3390]),
			.NE(gen[3391]),

			.O(gen[3484]),
			.E(gen[3486]),

			.SO(gen[3579]),
			.S(gen[3580]),
			.SE(gen[3581]),

			.SELF(gen[3485]),
			.cell_state(gen[3485])
		); 

/******************* CELL 3486 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3486 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3390]),
			.N(gen[3391]),
			.NE(gen[3392]),

			.O(gen[3485]),
			.E(gen[3487]),

			.SO(gen[3580]),
			.S(gen[3581]),
			.SE(gen[3582]),

			.SELF(gen[3486]),
			.cell_state(gen[3486])
		); 

/******************* CELL 3487 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3487 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3391]),
			.N(gen[3392]),
			.NE(gen[3393]),

			.O(gen[3486]),
			.E(gen[3488]),

			.SO(gen[3581]),
			.S(gen[3582]),
			.SE(gen[3583]),

			.SELF(gen[3487]),
			.cell_state(gen[3487])
		); 

/******************* CELL 3488 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3488 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3392]),
			.N(gen[3393]),
			.NE(gen[3394]),

			.O(gen[3487]),
			.E(gen[3489]),

			.SO(gen[3582]),
			.S(gen[3583]),
			.SE(gen[3584]),

			.SELF(gen[3488]),
			.cell_state(gen[3488])
		); 

/******************* CELL 3489 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3489 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3393]),
			.N(gen[3394]),
			.NE(gen[3395]),

			.O(gen[3488]),
			.E(gen[3490]),

			.SO(gen[3583]),
			.S(gen[3584]),
			.SE(gen[3585]),

			.SELF(gen[3489]),
			.cell_state(gen[3489])
		); 

/******************* CELL 3490 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3490 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3394]),
			.N(gen[3395]),
			.NE(gen[3396]),

			.O(gen[3489]),
			.E(gen[3491]),

			.SO(gen[3584]),
			.S(gen[3585]),
			.SE(gen[3586]),

			.SELF(gen[3490]),
			.cell_state(gen[3490])
		); 

/******************* CELL 3491 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3491 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3395]),
			.N(gen[3396]),
			.NE(gen[3397]),

			.O(gen[3490]),
			.E(gen[3492]),

			.SO(gen[3585]),
			.S(gen[3586]),
			.SE(gen[3587]),

			.SELF(gen[3491]),
			.cell_state(gen[3491])
		); 

/******************* CELL 3492 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3492 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3396]),
			.N(gen[3397]),
			.NE(gen[3398]),

			.O(gen[3491]),
			.E(gen[3493]),

			.SO(gen[3586]),
			.S(gen[3587]),
			.SE(gen[3588]),

			.SELF(gen[3492]),
			.cell_state(gen[3492])
		); 

/******************* CELL 3493 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3493 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3397]),
			.N(gen[3398]),
			.NE(gen[3399]),

			.O(gen[3492]),
			.E(gen[3494]),

			.SO(gen[3587]),
			.S(gen[3588]),
			.SE(gen[3589]),

			.SELF(gen[3493]),
			.cell_state(gen[3493])
		); 

/******************* CELL 3494 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3494 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3398]),
			.N(gen[3399]),
			.NE(gen[3400]),

			.O(gen[3493]),
			.E(gen[3495]),

			.SO(gen[3588]),
			.S(gen[3589]),
			.SE(gen[3590]),

			.SELF(gen[3494]),
			.cell_state(gen[3494])
		); 

/******************* CELL 3495 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3495 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3399]),
			.N(gen[3400]),
			.NE(gen[3401]),

			.O(gen[3494]),
			.E(gen[3496]),

			.SO(gen[3589]),
			.S(gen[3590]),
			.SE(gen[3591]),

			.SELF(gen[3495]),
			.cell_state(gen[3495])
		); 

/******************* CELL 3496 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3496 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3400]),
			.N(gen[3401]),
			.NE(gen[3402]),

			.O(gen[3495]),
			.E(gen[3497]),

			.SO(gen[3590]),
			.S(gen[3591]),
			.SE(gen[3592]),

			.SELF(gen[3496]),
			.cell_state(gen[3496])
		); 

/******************* CELL 3497 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3497 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3401]),
			.N(gen[3402]),
			.NE(gen[3403]),

			.O(gen[3496]),
			.E(gen[3498]),

			.SO(gen[3591]),
			.S(gen[3592]),
			.SE(gen[3593]),

			.SELF(gen[3497]),
			.cell_state(gen[3497])
		); 

/******************* CELL 3498 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3498 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3402]),
			.N(gen[3403]),
			.NE(gen[3404]),

			.O(gen[3497]),
			.E(gen[3499]),

			.SO(gen[3592]),
			.S(gen[3593]),
			.SE(gen[3594]),

			.SELF(gen[3498]),
			.cell_state(gen[3498])
		); 

/******************* CELL 3499 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3499 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3403]),
			.N(gen[3404]),
			.NE(gen[3405]),

			.O(gen[3498]),
			.E(gen[3500]),

			.SO(gen[3593]),
			.S(gen[3594]),
			.SE(gen[3595]),

			.SELF(gen[3499]),
			.cell_state(gen[3499])
		); 

/******************* CELL 3500 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3500 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3404]),
			.N(gen[3405]),
			.NE(gen[3406]),

			.O(gen[3499]),
			.E(gen[3501]),

			.SO(gen[3594]),
			.S(gen[3595]),
			.SE(gen[3596]),

			.SELF(gen[3500]),
			.cell_state(gen[3500])
		); 

/******************* CELL 3501 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3501 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3405]),
			.N(gen[3406]),
			.NE(gen[3407]),

			.O(gen[3500]),
			.E(gen[3502]),

			.SO(gen[3595]),
			.S(gen[3596]),
			.SE(gen[3597]),

			.SELF(gen[3501]),
			.cell_state(gen[3501])
		); 

/******************* CELL 3502 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3502 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3406]),
			.N(gen[3407]),
			.NE(gen[3408]),

			.O(gen[3501]),
			.E(gen[3503]),

			.SO(gen[3596]),
			.S(gen[3597]),
			.SE(gen[3598]),

			.SELF(gen[3502]),
			.cell_state(gen[3502])
		); 

/******************* CELL 3503 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3503 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3407]),
			.N(gen[3408]),
			.NE(gen[3409]),

			.O(gen[3502]),
			.E(gen[3504]),

			.SO(gen[3597]),
			.S(gen[3598]),
			.SE(gen[3599]),

			.SELF(gen[3503]),
			.cell_state(gen[3503])
		); 

/******************* CELL 3504 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3504 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3408]),
			.N(gen[3409]),
			.NE(gen[3410]),

			.O(gen[3503]),
			.E(gen[3505]),

			.SO(gen[3598]),
			.S(gen[3599]),
			.SE(gen[3600]),

			.SELF(gen[3504]),
			.cell_state(gen[3504])
		); 

/******************* CELL 3505 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3505 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3409]),
			.N(gen[3410]),
			.NE(gen[3411]),

			.O(gen[3504]),
			.E(gen[3506]),

			.SO(gen[3599]),
			.S(gen[3600]),
			.SE(gen[3601]),

			.SELF(gen[3505]),
			.cell_state(gen[3505])
		); 

/******************* CELL 3506 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3506 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3410]),
			.N(gen[3411]),
			.NE(gen[3412]),

			.O(gen[3505]),
			.E(gen[3507]),

			.SO(gen[3600]),
			.S(gen[3601]),
			.SE(gen[3602]),

			.SELF(gen[3506]),
			.cell_state(gen[3506])
		); 

/******************* CELL 3507 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3507 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3411]),
			.N(gen[3412]),
			.NE(gen[3413]),

			.O(gen[3506]),
			.E(gen[3508]),

			.SO(gen[3601]),
			.S(gen[3602]),
			.SE(gen[3603]),

			.SELF(gen[3507]),
			.cell_state(gen[3507])
		); 

/******************* CELL 3508 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3508 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3412]),
			.N(gen[3413]),
			.NE(gen[3414]),

			.O(gen[3507]),
			.E(gen[3509]),

			.SO(gen[3602]),
			.S(gen[3603]),
			.SE(gen[3604]),

			.SELF(gen[3508]),
			.cell_state(gen[3508])
		); 

/******************* CELL 3509 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3509 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3413]),
			.N(gen[3414]),
			.NE(gen[3415]),

			.O(gen[3508]),
			.E(gen[3510]),

			.SO(gen[3603]),
			.S(gen[3604]),
			.SE(gen[3605]),

			.SELF(gen[3509]),
			.cell_state(gen[3509])
		); 

/******************* CELL 3510 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3510 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3414]),
			.N(gen[3415]),
			.NE(gen[3416]),

			.O(gen[3509]),
			.E(gen[3511]),

			.SO(gen[3604]),
			.S(gen[3605]),
			.SE(gen[3606]),

			.SELF(gen[3510]),
			.cell_state(gen[3510])
		); 

/******************* CELL 3511 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3511 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3415]),
			.N(gen[3416]),
			.NE(gen[3417]),

			.O(gen[3510]),
			.E(gen[3512]),

			.SO(gen[3605]),
			.S(gen[3606]),
			.SE(gen[3607]),

			.SELF(gen[3511]),
			.cell_state(gen[3511])
		); 

/******************* CELL 3512 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3512 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3416]),
			.N(gen[3417]),
			.NE(gen[3418]),

			.O(gen[3511]),
			.E(gen[3513]),

			.SO(gen[3606]),
			.S(gen[3607]),
			.SE(gen[3608]),

			.SELF(gen[3512]),
			.cell_state(gen[3512])
		); 

/******************* CELL 3513 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3513 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3417]),
			.N(gen[3418]),
			.NE(gen[3419]),

			.O(gen[3512]),
			.E(gen[3514]),

			.SO(gen[3607]),
			.S(gen[3608]),
			.SE(gen[3609]),

			.SELF(gen[3513]),
			.cell_state(gen[3513])
		); 

/******************* CELL 3514 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3514 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3418]),
			.N(gen[3419]),
			.NE(gen[3418]),

			.O(gen[3513]),
			.E(gen[3513]),

			.SO(gen[3608]),
			.S(gen[3609]),
			.SE(gen[3608]),

			.SELF(gen[3514]),
			.cell_state(gen[3514])
		); 

/******************* CELL 3515 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3515 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3421]),
			.N(gen[3420]),
			.NE(gen[3421]),

			.O(gen[3516]),
			.E(gen[3516]),

			.SO(gen[3611]),
			.S(gen[3610]),
			.SE(gen[3611]),

			.SELF(gen[3515]),
			.cell_state(gen[3515])
		); 

/******************* CELL 3516 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3516 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3420]),
			.N(gen[3421]),
			.NE(gen[3422]),

			.O(gen[3515]),
			.E(gen[3517]),

			.SO(gen[3610]),
			.S(gen[3611]),
			.SE(gen[3612]),

			.SELF(gen[3516]),
			.cell_state(gen[3516])
		); 

/******************* CELL 3517 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3517 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3421]),
			.N(gen[3422]),
			.NE(gen[3423]),

			.O(gen[3516]),
			.E(gen[3518]),

			.SO(gen[3611]),
			.S(gen[3612]),
			.SE(gen[3613]),

			.SELF(gen[3517]),
			.cell_state(gen[3517])
		); 

/******************* CELL 3518 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3518 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3422]),
			.N(gen[3423]),
			.NE(gen[3424]),

			.O(gen[3517]),
			.E(gen[3519]),

			.SO(gen[3612]),
			.S(gen[3613]),
			.SE(gen[3614]),

			.SELF(gen[3518]),
			.cell_state(gen[3518])
		); 

/******************* CELL 3519 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3519 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3423]),
			.N(gen[3424]),
			.NE(gen[3425]),

			.O(gen[3518]),
			.E(gen[3520]),

			.SO(gen[3613]),
			.S(gen[3614]),
			.SE(gen[3615]),

			.SELF(gen[3519]),
			.cell_state(gen[3519])
		); 

/******************* CELL 3520 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3520 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3424]),
			.N(gen[3425]),
			.NE(gen[3426]),

			.O(gen[3519]),
			.E(gen[3521]),

			.SO(gen[3614]),
			.S(gen[3615]),
			.SE(gen[3616]),

			.SELF(gen[3520]),
			.cell_state(gen[3520])
		); 

/******************* CELL 3521 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3521 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3425]),
			.N(gen[3426]),
			.NE(gen[3427]),

			.O(gen[3520]),
			.E(gen[3522]),

			.SO(gen[3615]),
			.S(gen[3616]),
			.SE(gen[3617]),

			.SELF(gen[3521]),
			.cell_state(gen[3521])
		); 

/******************* CELL 3522 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3522 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3426]),
			.N(gen[3427]),
			.NE(gen[3428]),

			.O(gen[3521]),
			.E(gen[3523]),

			.SO(gen[3616]),
			.S(gen[3617]),
			.SE(gen[3618]),

			.SELF(gen[3522]),
			.cell_state(gen[3522])
		); 

/******************* CELL 3523 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3523 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3427]),
			.N(gen[3428]),
			.NE(gen[3429]),

			.O(gen[3522]),
			.E(gen[3524]),

			.SO(gen[3617]),
			.S(gen[3618]),
			.SE(gen[3619]),

			.SELF(gen[3523]),
			.cell_state(gen[3523])
		); 

/******************* CELL 3524 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3524 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3428]),
			.N(gen[3429]),
			.NE(gen[3430]),

			.O(gen[3523]),
			.E(gen[3525]),

			.SO(gen[3618]),
			.S(gen[3619]),
			.SE(gen[3620]),

			.SELF(gen[3524]),
			.cell_state(gen[3524])
		); 

/******************* CELL 3525 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3525 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3429]),
			.N(gen[3430]),
			.NE(gen[3431]),

			.O(gen[3524]),
			.E(gen[3526]),

			.SO(gen[3619]),
			.S(gen[3620]),
			.SE(gen[3621]),

			.SELF(gen[3525]),
			.cell_state(gen[3525])
		); 

/******************* CELL 3526 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3526 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3430]),
			.N(gen[3431]),
			.NE(gen[3432]),

			.O(gen[3525]),
			.E(gen[3527]),

			.SO(gen[3620]),
			.S(gen[3621]),
			.SE(gen[3622]),

			.SELF(gen[3526]),
			.cell_state(gen[3526])
		); 

/******************* CELL 3527 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3527 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3431]),
			.N(gen[3432]),
			.NE(gen[3433]),

			.O(gen[3526]),
			.E(gen[3528]),

			.SO(gen[3621]),
			.S(gen[3622]),
			.SE(gen[3623]),

			.SELF(gen[3527]),
			.cell_state(gen[3527])
		); 

/******************* CELL 3528 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3528 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3432]),
			.N(gen[3433]),
			.NE(gen[3434]),

			.O(gen[3527]),
			.E(gen[3529]),

			.SO(gen[3622]),
			.S(gen[3623]),
			.SE(gen[3624]),

			.SELF(gen[3528]),
			.cell_state(gen[3528])
		); 

/******************* CELL 3529 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3529 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3433]),
			.N(gen[3434]),
			.NE(gen[3435]),

			.O(gen[3528]),
			.E(gen[3530]),

			.SO(gen[3623]),
			.S(gen[3624]),
			.SE(gen[3625]),

			.SELF(gen[3529]),
			.cell_state(gen[3529])
		); 

/******************* CELL 3530 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3530 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3434]),
			.N(gen[3435]),
			.NE(gen[3436]),

			.O(gen[3529]),
			.E(gen[3531]),

			.SO(gen[3624]),
			.S(gen[3625]),
			.SE(gen[3626]),

			.SELF(gen[3530]),
			.cell_state(gen[3530])
		); 

/******************* CELL 3531 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3531 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3435]),
			.N(gen[3436]),
			.NE(gen[3437]),

			.O(gen[3530]),
			.E(gen[3532]),

			.SO(gen[3625]),
			.S(gen[3626]),
			.SE(gen[3627]),

			.SELF(gen[3531]),
			.cell_state(gen[3531])
		); 

/******************* CELL 3532 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3532 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3436]),
			.N(gen[3437]),
			.NE(gen[3438]),

			.O(gen[3531]),
			.E(gen[3533]),

			.SO(gen[3626]),
			.S(gen[3627]),
			.SE(gen[3628]),

			.SELF(gen[3532]),
			.cell_state(gen[3532])
		); 

/******************* CELL 3533 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3533 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3437]),
			.N(gen[3438]),
			.NE(gen[3439]),

			.O(gen[3532]),
			.E(gen[3534]),

			.SO(gen[3627]),
			.S(gen[3628]),
			.SE(gen[3629]),

			.SELF(gen[3533]),
			.cell_state(gen[3533])
		); 

/******************* CELL 3534 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3534 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3438]),
			.N(gen[3439]),
			.NE(gen[3440]),

			.O(gen[3533]),
			.E(gen[3535]),

			.SO(gen[3628]),
			.S(gen[3629]),
			.SE(gen[3630]),

			.SELF(gen[3534]),
			.cell_state(gen[3534])
		); 

/******************* CELL 3535 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3535 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3439]),
			.N(gen[3440]),
			.NE(gen[3441]),

			.O(gen[3534]),
			.E(gen[3536]),

			.SO(gen[3629]),
			.S(gen[3630]),
			.SE(gen[3631]),

			.SELF(gen[3535]),
			.cell_state(gen[3535])
		); 

/******************* CELL 3536 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3536 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3440]),
			.N(gen[3441]),
			.NE(gen[3442]),

			.O(gen[3535]),
			.E(gen[3537]),

			.SO(gen[3630]),
			.S(gen[3631]),
			.SE(gen[3632]),

			.SELF(gen[3536]),
			.cell_state(gen[3536])
		); 

/******************* CELL 3537 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3537 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3441]),
			.N(gen[3442]),
			.NE(gen[3443]),

			.O(gen[3536]),
			.E(gen[3538]),

			.SO(gen[3631]),
			.S(gen[3632]),
			.SE(gen[3633]),

			.SELF(gen[3537]),
			.cell_state(gen[3537])
		); 

/******************* CELL 3538 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3538 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3442]),
			.N(gen[3443]),
			.NE(gen[3444]),

			.O(gen[3537]),
			.E(gen[3539]),

			.SO(gen[3632]),
			.S(gen[3633]),
			.SE(gen[3634]),

			.SELF(gen[3538]),
			.cell_state(gen[3538])
		); 

/******************* CELL 3539 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3539 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3443]),
			.N(gen[3444]),
			.NE(gen[3445]),

			.O(gen[3538]),
			.E(gen[3540]),

			.SO(gen[3633]),
			.S(gen[3634]),
			.SE(gen[3635]),

			.SELF(gen[3539]),
			.cell_state(gen[3539])
		); 

/******************* CELL 3540 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3540 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3444]),
			.N(gen[3445]),
			.NE(gen[3446]),

			.O(gen[3539]),
			.E(gen[3541]),

			.SO(gen[3634]),
			.S(gen[3635]),
			.SE(gen[3636]),

			.SELF(gen[3540]),
			.cell_state(gen[3540])
		); 

/******************* CELL 3541 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3541 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3445]),
			.N(gen[3446]),
			.NE(gen[3447]),

			.O(gen[3540]),
			.E(gen[3542]),

			.SO(gen[3635]),
			.S(gen[3636]),
			.SE(gen[3637]),

			.SELF(gen[3541]),
			.cell_state(gen[3541])
		); 

/******************* CELL 3542 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3542 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3446]),
			.N(gen[3447]),
			.NE(gen[3448]),

			.O(gen[3541]),
			.E(gen[3543]),

			.SO(gen[3636]),
			.S(gen[3637]),
			.SE(gen[3638]),

			.SELF(gen[3542]),
			.cell_state(gen[3542])
		); 

/******************* CELL 3543 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3543 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3447]),
			.N(gen[3448]),
			.NE(gen[3449]),

			.O(gen[3542]),
			.E(gen[3544]),

			.SO(gen[3637]),
			.S(gen[3638]),
			.SE(gen[3639]),

			.SELF(gen[3543]),
			.cell_state(gen[3543])
		); 

/******************* CELL 3544 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3544 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3448]),
			.N(gen[3449]),
			.NE(gen[3450]),

			.O(gen[3543]),
			.E(gen[3545]),

			.SO(gen[3638]),
			.S(gen[3639]),
			.SE(gen[3640]),

			.SELF(gen[3544]),
			.cell_state(gen[3544])
		); 

/******************* CELL 3545 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3545 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3449]),
			.N(gen[3450]),
			.NE(gen[3451]),

			.O(gen[3544]),
			.E(gen[3546]),

			.SO(gen[3639]),
			.S(gen[3640]),
			.SE(gen[3641]),

			.SELF(gen[3545]),
			.cell_state(gen[3545])
		); 

/******************* CELL 3546 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3546 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3450]),
			.N(gen[3451]),
			.NE(gen[3452]),

			.O(gen[3545]),
			.E(gen[3547]),

			.SO(gen[3640]),
			.S(gen[3641]),
			.SE(gen[3642]),

			.SELF(gen[3546]),
			.cell_state(gen[3546])
		); 

/******************* CELL 3547 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3547 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3451]),
			.N(gen[3452]),
			.NE(gen[3453]),

			.O(gen[3546]),
			.E(gen[3548]),

			.SO(gen[3641]),
			.S(gen[3642]),
			.SE(gen[3643]),

			.SELF(gen[3547]),
			.cell_state(gen[3547])
		); 

/******************* CELL 3548 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3548 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3452]),
			.N(gen[3453]),
			.NE(gen[3454]),

			.O(gen[3547]),
			.E(gen[3549]),

			.SO(gen[3642]),
			.S(gen[3643]),
			.SE(gen[3644]),

			.SELF(gen[3548]),
			.cell_state(gen[3548])
		); 

/******************* CELL 3549 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3549 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3453]),
			.N(gen[3454]),
			.NE(gen[3455]),

			.O(gen[3548]),
			.E(gen[3550]),

			.SO(gen[3643]),
			.S(gen[3644]),
			.SE(gen[3645]),

			.SELF(gen[3549]),
			.cell_state(gen[3549])
		); 

/******************* CELL 3550 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3550 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3454]),
			.N(gen[3455]),
			.NE(gen[3456]),

			.O(gen[3549]),
			.E(gen[3551]),

			.SO(gen[3644]),
			.S(gen[3645]),
			.SE(gen[3646]),

			.SELF(gen[3550]),
			.cell_state(gen[3550])
		); 

/******************* CELL 3551 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3551 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3455]),
			.N(gen[3456]),
			.NE(gen[3457]),

			.O(gen[3550]),
			.E(gen[3552]),

			.SO(gen[3645]),
			.S(gen[3646]),
			.SE(gen[3647]),

			.SELF(gen[3551]),
			.cell_state(gen[3551])
		); 

/******************* CELL 3552 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3552 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3456]),
			.N(gen[3457]),
			.NE(gen[3458]),

			.O(gen[3551]),
			.E(gen[3553]),

			.SO(gen[3646]),
			.S(gen[3647]),
			.SE(gen[3648]),

			.SELF(gen[3552]),
			.cell_state(gen[3552])
		); 

/******************* CELL 3553 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3553 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3457]),
			.N(gen[3458]),
			.NE(gen[3459]),

			.O(gen[3552]),
			.E(gen[3554]),

			.SO(gen[3647]),
			.S(gen[3648]),
			.SE(gen[3649]),

			.SELF(gen[3553]),
			.cell_state(gen[3553])
		); 

/******************* CELL 3554 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3554 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3458]),
			.N(gen[3459]),
			.NE(gen[3460]),

			.O(gen[3553]),
			.E(gen[3555]),

			.SO(gen[3648]),
			.S(gen[3649]),
			.SE(gen[3650]),

			.SELF(gen[3554]),
			.cell_state(gen[3554])
		); 

/******************* CELL 3555 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3555 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3459]),
			.N(gen[3460]),
			.NE(gen[3461]),

			.O(gen[3554]),
			.E(gen[3556]),

			.SO(gen[3649]),
			.S(gen[3650]),
			.SE(gen[3651]),

			.SELF(gen[3555]),
			.cell_state(gen[3555])
		); 

/******************* CELL 3556 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3556 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3460]),
			.N(gen[3461]),
			.NE(gen[3462]),

			.O(gen[3555]),
			.E(gen[3557]),

			.SO(gen[3650]),
			.S(gen[3651]),
			.SE(gen[3652]),

			.SELF(gen[3556]),
			.cell_state(gen[3556])
		); 

/******************* CELL 3557 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3557 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3461]),
			.N(gen[3462]),
			.NE(gen[3463]),

			.O(gen[3556]),
			.E(gen[3558]),

			.SO(gen[3651]),
			.S(gen[3652]),
			.SE(gen[3653]),

			.SELF(gen[3557]),
			.cell_state(gen[3557])
		); 

/******************* CELL 3558 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3558 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3462]),
			.N(gen[3463]),
			.NE(gen[3464]),

			.O(gen[3557]),
			.E(gen[3559]),

			.SO(gen[3652]),
			.S(gen[3653]),
			.SE(gen[3654]),

			.SELF(gen[3558]),
			.cell_state(gen[3558])
		); 

/******************* CELL 3559 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3559 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3463]),
			.N(gen[3464]),
			.NE(gen[3465]),

			.O(gen[3558]),
			.E(gen[3560]),

			.SO(gen[3653]),
			.S(gen[3654]),
			.SE(gen[3655]),

			.SELF(gen[3559]),
			.cell_state(gen[3559])
		); 

/******************* CELL 3560 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3560 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3464]),
			.N(gen[3465]),
			.NE(gen[3466]),

			.O(gen[3559]),
			.E(gen[3561]),

			.SO(gen[3654]),
			.S(gen[3655]),
			.SE(gen[3656]),

			.SELF(gen[3560]),
			.cell_state(gen[3560])
		); 

/******************* CELL 3561 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3561 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3465]),
			.N(gen[3466]),
			.NE(gen[3467]),

			.O(gen[3560]),
			.E(gen[3562]),

			.SO(gen[3655]),
			.S(gen[3656]),
			.SE(gen[3657]),

			.SELF(gen[3561]),
			.cell_state(gen[3561])
		); 

/******************* CELL 3562 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3562 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3466]),
			.N(gen[3467]),
			.NE(gen[3468]),

			.O(gen[3561]),
			.E(gen[3563]),

			.SO(gen[3656]),
			.S(gen[3657]),
			.SE(gen[3658]),

			.SELF(gen[3562]),
			.cell_state(gen[3562])
		); 

/******************* CELL 3563 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3563 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3467]),
			.N(gen[3468]),
			.NE(gen[3469]),

			.O(gen[3562]),
			.E(gen[3564]),

			.SO(gen[3657]),
			.S(gen[3658]),
			.SE(gen[3659]),

			.SELF(gen[3563]),
			.cell_state(gen[3563])
		); 

/******************* CELL 3564 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3564 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3468]),
			.N(gen[3469]),
			.NE(gen[3470]),

			.O(gen[3563]),
			.E(gen[3565]),

			.SO(gen[3658]),
			.S(gen[3659]),
			.SE(gen[3660]),

			.SELF(gen[3564]),
			.cell_state(gen[3564])
		); 

/******************* CELL 3565 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3565 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3469]),
			.N(gen[3470]),
			.NE(gen[3471]),

			.O(gen[3564]),
			.E(gen[3566]),

			.SO(gen[3659]),
			.S(gen[3660]),
			.SE(gen[3661]),

			.SELF(gen[3565]),
			.cell_state(gen[3565])
		); 

/******************* CELL 3566 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3566 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3470]),
			.N(gen[3471]),
			.NE(gen[3472]),

			.O(gen[3565]),
			.E(gen[3567]),

			.SO(gen[3660]),
			.S(gen[3661]),
			.SE(gen[3662]),

			.SELF(gen[3566]),
			.cell_state(gen[3566])
		); 

/******************* CELL 3567 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3567 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3471]),
			.N(gen[3472]),
			.NE(gen[3473]),

			.O(gen[3566]),
			.E(gen[3568]),

			.SO(gen[3661]),
			.S(gen[3662]),
			.SE(gen[3663]),

			.SELF(gen[3567]),
			.cell_state(gen[3567])
		); 

/******************* CELL 3568 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3568 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3472]),
			.N(gen[3473]),
			.NE(gen[3474]),

			.O(gen[3567]),
			.E(gen[3569]),

			.SO(gen[3662]),
			.S(gen[3663]),
			.SE(gen[3664]),

			.SELF(gen[3568]),
			.cell_state(gen[3568])
		); 

/******************* CELL 3569 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3569 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3473]),
			.N(gen[3474]),
			.NE(gen[3475]),

			.O(gen[3568]),
			.E(gen[3570]),

			.SO(gen[3663]),
			.S(gen[3664]),
			.SE(gen[3665]),

			.SELF(gen[3569]),
			.cell_state(gen[3569])
		); 

/******************* CELL 3570 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3570 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3474]),
			.N(gen[3475]),
			.NE(gen[3476]),

			.O(gen[3569]),
			.E(gen[3571]),

			.SO(gen[3664]),
			.S(gen[3665]),
			.SE(gen[3666]),

			.SELF(gen[3570]),
			.cell_state(gen[3570])
		); 

/******************* CELL 3571 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3571 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3475]),
			.N(gen[3476]),
			.NE(gen[3477]),

			.O(gen[3570]),
			.E(gen[3572]),

			.SO(gen[3665]),
			.S(gen[3666]),
			.SE(gen[3667]),

			.SELF(gen[3571]),
			.cell_state(gen[3571])
		); 

/******************* CELL 3572 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3572 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3476]),
			.N(gen[3477]),
			.NE(gen[3478]),

			.O(gen[3571]),
			.E(gen[3573]),

			.SO(gen[3666]),
			.S(gen[3667]),
			.SE(gen[3668]),

			.SELF(gen[3572]),
			.cell_state(gen[3572])
		); 

/******************* CELL 3573 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3573 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3477]),
			.N(gen[3478]),
			.NE(gen[3479]),

			.O(gen[3572]),
			.E(gen[3574]),

			.SO(gen[3667]),
			.S(gen[3668]),
			.SE(gen[3669]),

			.SELF(gen[3573]),
			.cell_state(gen[3573])
		); 

/******************* CELL 3574 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3574 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3478]),
			.N(gen[3479]),
			.NE(gen[3480]),

			.O(gen[3573]),
			.E(gen[3575]),

			.SO(gen[3668]),
			.S(gen[3669]),
			.SE(gen[3670]),

			.SELF(gen[3574]),
			.cell_state(gen[3574])
		); 

/******************* CELL 3575 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3575 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3479]),
			.N(gen[3480]),
			.NE(gen[3481]),

			.O(gen[3574]),
			.E(gen[3576]),

			.SO(gen[3669]),
			.S(gen[3670]),
			.SE(gen[3671]),

			.SELF(gen[3575]),
			.cell_state(gen[3575])
		); 

/******************* CELL 3576 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3576 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3480]),
			.N(gen[3481]),
			.NE(gen[3482]),

			.O(gen[3575]),
			.E(gen[3577]),

			.SO(gen[3670]),
			.S(gen[3671]),
			.SE(gen[3672]),

			.SELF(gen[3576]),
			.cell_state(gen[3576])
		); 

/******************* CELL 3577 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3577 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3481]),
			.N(gen[3482]),
			.NE(gen[3483]),

			.O(gen[3576]),
			.E(gen[3578]),

			.SO(gen[3671]),
			.S(gen[3672]),
			.SE(gen[3673]),

			.SELF(gen[3577]),
			.cell_state(gen[3577])
		); 

/******************* CELL 3578 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3578 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3482]),
			.N(gen[3483]),
			.NE(gen[3484]),

			.O(gen[3577]),
			.E(gen[3579]),

			.SO(gen[3672]),
			.S(gen[3673]),
			.SE(gen[3674]),

			.SELF(gen[3578]),
			.cell_state(gen[3578])
		); 

/******************* CELL 3579 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3579 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3483]),
			.N(gen[3484]),
			.NE(gen[3485]),

			.O(gen[3578]),
			.E(gen[3580]),

			.SO(gen[3673]),
			.S(gen[3674]),
			.SE(gen[3675]),

			.SELF(gen[3579]),
			.cell_state(gen[3579])
		); 

/******************* CELL 3580 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3580 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3484]),
			.N(gen[3485]),
			.NE(gen[3486]),

			.O(gen[3579]),
			.E(gen[3581]),

			.SO(gen[3674]),
			.S(gen[3675]),
			.SE(gen[3676]),

			.SELF(gen[3580]),
			.cell_state(gen[3580])
		); 

/******************* CELL 3581 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3581 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3485]),
			.N(gen[3486]),
			.NE(gen[3487]),

			.O(gen[3580]),
			.E(gen[3582]),

			.SO(gen[3675]),
			.S(gen[3676]),
			.SE(gen[3677]),

			.SELF(gen[3581]),
			.cell_state(gen[3581])
		); 

/******************* CELL 3582 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3582 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3486]),
			.N(gen[3487]),
			.NE(gen[3488]),

			.O(gen[3581]),
			.E(gen[3583]),

			.SO(gen[3676]),
			.S(gen[3677]),
			.SE(gen[3678]),

			.SELF(gen[3582]),
			.cell_state(gen[3582])
		); 

/******************* CELL 3583 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3583 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3487]),
			.N(gen[3488]),
			.NE(gen[3489]),

			.O(gen[3582]),
			.E(gen[3584]),

			.SO(gen[3677]),
			.S(gen[3678]),
			.SE(gen[3679]),

			.SELF(gen[3583]),
			.cell_state(gen[3583])
		); 

/******************* CELL 3584 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3584 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3488]),
			.N(gen[3489]),
			.NE(gen[3490]),

			.O(gen[3583]),
			.E(gen[3585]),

			.SO(gen[3678]),
			.S(gen[3679]),
			.SE(gen[3680]),

			.SELF(gen[3584]),
			.cell_state(gen[3584])
		); 

/******************* CELL 3585 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3585 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3489]),
			.N(gen[3490]),
			.NE(gen[3491]),

			.O(gen[3584]),
			.E(gen[3586]),

			.SO(gen[3679]),
			.S(gen[3680]),
			.SE(gen[3681]),

			.SELF(gen[3585]),
			.cell_state(gen[3585])
		); 

/******************* CELL 3586 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3586 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3490]),
			.N(gen[3491]),
			.NE(gen[3492]),

			.O(gen[3585]),
			.E(gen[3587]),

			.SO(gen[3680]),
			.S(gen[3681]),
			.SE(gen[3682]),

			.SELF(gen[3586]),
			.cell_state(gen[3586])
		); 

/******************* CELL 3587 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3587 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3491]),
			.N(gen[3492]),
			.NE(gen[3493]),

			.O(gen[3586]),
			.E(gen[3588]),

			.SO(gen[3681]),
			.S(gen[3682]),
			.SE(gen[3683]),

			.SELF(gen[3587]),
			.cell_state(gen[3587])
		); 

/******************* CELL 3588 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3588 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3492]),
			.N(gen[3493]),
			.NE(gen[3494]),

			.O(gen[3587]),
			.E(gen[3589]),

			.SO(gen[3682]),
			.S(gen[3683]),
			.SE(gen[3684]),

			.SELF(gen[3588]),
			.cell_state(gen[3588])
		); 

/******************* CELL 3589 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3589 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3493]),
			.N(gen[3494]),
			.NE(gen[3495]),

			.O(gen[3588]),
			.E(gen[3590]),

			.SO(gen[3683]),
			.S(gen[3684]),
			.SE(gen[3685]),

			.SELF(gen[3589]),
			.cell_state(gen[3589])
		); 

/******************* CELL 3590 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3590 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3494]),
			.N(gen[3495]),
			.NE(gen[3496]),

			.O(gen[3589]),
			.E(gen[3591]),

			.SO(gen[3684]),
			.S(gen[3685]),
			.SE(gen[3686]),

			.SELF(gen[3590]),
			.cell_state(gen[3590])
		); 

/******************* CELL 3591 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3591 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3495]),
			.N(gen[3496]),
			.NE(gen[3497]),

			.O(gen[3590]),
			.E(gen[3592]),

			.SO(gen[3685]),
			.S(gen[3686]),
			.SE(gen[3687]),

			.SELF(gen[3591]),
			.cell_state(gen[3591])
		); 

/******************* CELL 3592 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3592 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3496]),
			.N(gen[3497]),
			.NE(gen[3498]),

			.O(gen[3591]),
			.E(gen[3593]),

			.SO(gen[3686]),
			.S(gen[3687]),
			.SE(gen[3688]),

			.SELF(gen[3592]),
			.cell_state(gen[3592])
		); 

/******************* CELL 3593 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3593 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3497]),
			.N(gen[3498]),
			.NE(gen[3499]),

			.O(gen[3592]),
			.E(gen[3594]),

			.SO(gen[3687]),
			.S(gen[3688]),
			.SE(gen[3689]),

			.SELF(gen[3593]),
			.cell_state(gen[3593])
		); 

/******************* CELL 3594 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3594 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3498]),
			.N(gen[3499]),
			.NE(gen[3500]),

			.O(gen[3593]),
			.E(gen[3595]),

			.SO(gen[3688]),
			.S(gen[3689]),
			.SE(gen[3690]),

			.SELF(gen[3594]),
			.cell_state(gen[3594])
		); 

/******************* CELL 3595 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3595 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3499]),
			.N(gen[3500]),
			.NE(gen[3501]),

			.O(gen[3594]),
			.E(gen[3596]),

			.SO(gen[3689]),
			.S(gen[3690]),
			.SE(gen[3691]),

			.SELF(gen[3595]),
			.cell_state(gen[3595])
		); 

/******************* CELL 3596 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3596 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3500]),
			.N(gen[3501]),
			.NE(gen[3502]),

			.O(gen[3595]),
			.E(gen[3597]),

			.SO(gen[3690]),
			.S(gen[3691]),
			.SE(gen[3692]),

			.SELF(gen[3596]),
			.cell_state(gen[3596])
		); 

/******************* CELL 3597 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3597 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3501]),
			.N(gen[3502]),
			.NE(gen[3503]),

			.O(gen[3596]),
			.E(gen[3598]),

			.SO(gen[3691]),
			.S(gen[3692]),
			.SE(gen[3693]),

			.SELF(gen[3597]),
			.cell_state(gen[3597])
		); 

/******************* CELL 3598 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3598 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3502]),
			.N(gen[3503]),
			.NE(gen[3504]),

			.O(gen[3597]),
			.E(gen[3599]),

			.SO(gen[3692]),
			.S(gen[3693]),
			.SE(gen[3694]),

			.SELF(gen[3598]),
			.cell_state(gen[3598])
		); 

/******************* CELL 3599 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3599 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3503]),
			.N(gen[3504]),
			.NE(gen[3505]),

			.O(gen[3598]),
			.E(gen[3600]),

			.SO(gen[3693]),
			.S(gen[3694]),
			.SE(gen[3695]),

			.SELF(gen[3599]),
			.cell_state(gen[3599])
		); 

/******************* CELL 3600 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3600 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3504]),
			.N(gen[3505]),
			.NE(gen[3506]),

			.O(gen[3599]),
			.E(gen[3601]),

			.SO(gen[3694]),
			.S(gen[3695]),
			.SE(gen[3696]),

			.SELF(gen[3600]),
			.cell_state(gen[3600])
		); 

/******************* CELL 3601 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3601 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3505]),
			.N(gen[3506]),
			.NE(gen[3507]),

			.O(gen[3600]),
			.E(gen[3602]),

			.SO(gen[3695]),
			.S(gen[3696]),
			.SE(gen[3697]),

			.SELF(gen[3601]),
			.cell_state(gen[3601])
		); 

/******************* CELL 3602 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3602 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3506]),
			.N(gen[3507]),
			.NE(gen[3508]),

			.O(gen[3601]),
			.E(gen[3603]),

			.SO(gen[3696]),
			.S(gen[3697]),
			.SE(gen[3698]),

			.SELF(gen[3602]),
			.cell_state(gen[3602])
		); 

/******************* CELL 3603 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3603 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3507]),
			.N(gen[3508]),
			.NE(gen[3509]),

			.O(gen[3602]),
			.E(gen[3604]),

			.SO(gen[3697]),
			.S(gen[3698]),
			.SE(gen[3699]),

			.SELF(gen[3603]),
			.cell_state(gen[3603])
		); 

/******************* CELL 3604 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3604 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3508]),
			.N(gen[3509]),
			.NE(gen[3510]),

			.O(gen[3603]),
			.E(gen[3605]),

			.SO(gen[3698]),
			.S(gen[3699]),
			.SE(gen[3700]),

			.SELF(gen[3604]),
			.cell_state(gen[3604])
		); 

/******************* CELL 3605 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3605 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3509]),
			.N(gen[3510]),
			.NE(gen[3511]),

			.O(gen[3604]),
			.E(gen[3606]),

			.SO(gen[3699]),
			.S(gen[3700]),
			.SE(gen[3701]),

			.SELF(gen[3605]),
			.cell_state(gen[3605])
		); 

/******************* CELL 3606 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3606 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3510]),
			.N(gen[3511]),
			.NE(gen[3512]),

			.O(gen[3605]),
			.E(gen[3607]),

			.SO(gen[3700]),
			.S(gen[3701]),
			.SE(gen[3702]),

			.SELF(gen[3606]),
			.cell_state(gen[3606])
		); 

/******************* CELL 3607 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3607 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3511]),
			.N(gen[3512]),
			.NE(gen[3513]),

			.O(gen[3606]),
			.E(gen[3608]),

			.SO(gen[3701]),
			.S(gen[3702]),
			.SE(gen[3703]),

			.SELF(gen[3607]),
			.cell_state(gen[3607])
		); 

/******************* CELL 3608 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3608 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3512]),
			.N(gen[3513]),
			.NE(gen[3514]),

			.O(gen[3607]),
			.E(gen[3609]),

			.SO(gen[3702]),
			.S(gen[3703]),
			.SE(gen[3704]),

			.SELF(gen[3608]),
			.cell_state(gen[3608])
		); 

/******************* CELL 3609 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3609 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3513]),
			.N(gen[3514]),
			.NE(gen[3513]),

			.O(gen[3608]),
			.E(gen[3608]),

			.SO(gen[3703]),
			.S(gen[3704]),
			.SE(gen[3703]),

			.SELF(gen[3609]),
			.cell_state(gen[3609])
		); 

/******************* CELL 3610 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3610 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3516]),
			.N(gen[3515]),
			.NE(gen[3516]),

			.O(gen[3611]),
			.E(gen[3611]),

			.SO(gen[3706]),
			.S(gen[3705]),
			.SE(gen[3706]),

			.SELF(gen[3610]),
			.cell_state(gen[3610])
		); 

/******************* CELL 3611 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3611 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3515]),
			.N(gen[3516]),
			.NE(gen[3517]),

			.O(gen[3610]),
			.E(gen[3612]),

			.SO(gen[3705]),
			.S(gen[3706]),
			.SE(gen[3707]),

			.SELF(gen[3611]),
			.cell_state(gen[3611])
		); 

/******************* CELL 3612 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3612 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3516]),
			.N(gen[3517]),
			.NE(gen[3518]),

			.O(gen[3611]),
			.E(gen[3613]),

			.SO(gen[3706]),
			.S(gen[3707]),
			.SE(gen[3708]),

			.SELF(gen[3612]),
			.cell_state(gen[3612])
		); 

/******************* CELL 3613 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3613 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3517]),
			.N(gen[3518]),
			.NE(gen[3519]),

			.O(gen[3612]),
			.E(gen[3614]),

			.SO(gen[3707]),
			.S(gen[3708]),
			.SE(gen[3709]),

			.SELF(gen[3613]),
			.cell_state(gen[3613])
		); 

/******************* CELL 3614 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3614 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3518]),
			.N(gen[3519]),
			.NE(gen[3520]),

			.O(gen[3613]),
			.E(gen[3615]),

			.SO(gen[3708]),
			.S(gen[3709]),
			.SE(gen[3710]),

			.SELF(gen[3614]),
			.cell_state(gen[3614])
		); 

/******************* CELL 3615 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3615 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3519]),
			.N(gen[3520]),
			.NE(gen[3521]),

			.O(gen[3614]),
			.E(gen[3616]),

			.SO(gen[3709]),
			.S(gen[3710]),
			.SE(gen[3711]),

			.SELF(gen[3615]),
			.cell_state(gen[3615])
		); 

/******************* CELL 3616 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3616 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3520]),
			.N(gen[3521]),
			.NE(gen[3522]),

			.O(gen[3615]),
			.E(gen[3617]),

			.SO(gen[3710]),
			.S(gen[3711]),
			.SE(gen[3712]),

			.SELF(gen[3616]),
			.cell_state(gen[3616])
		); 

/******************* CELL 3617 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3617 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3521]),
			.N(gen[3522]),
			.NE(gen[3523]),

			.O(gen[3616]),
			.E(gen[3618]),

			.SO(gen[3711]),
			.S(gen[3712]),
			.SE(gen[3713]),

			.SELF(gen[3617]),
			.cell_state(gen[3617])
		); 

/******************* CELL 3618 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3618 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3522]),
			.N(gen[3523]),
			.NE(gen[3524]),

			.O(gen[3617]),
			.E(gen[3619]),

			.SO(gen[3712]),
			.S(gen[3713]),
			.SE(gen[3714]),

			.SELF(gen[3618]),
			.cell_state(gen[3618])
		); 

/******************* CELL 3619 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3619 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3523]),
			.N(gen[3524]),
			.NE(gen[3525]),

			.O(gen[3618]),
			.E(gen[3620]),

			.SO(gen[3713]),
			.S(gen[3714]),
			.SE(gen[3715]),

			.SELF(gen[3619]),
			.cell_state(gen[3619])
		); 

/******************* CELL 3620 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3620 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3524]),
			.N(gen[3525]),
			.NE(gen[3526]),

			.O(gen[3619]),
			.E(gen[3621]),

			.SO(gen[3714]),
			.S(gen[3715]),
			.SE(gen[3716]),

			.SELF(gen[3620]),
			.cell_state(gen[3620])
		); 

/******************* CELL 3621 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3621 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3525]),
			.N(gen[3526]),
			.NE(gen[3527]),

			.O(gen[3620]),
			.E(gen[3622]),

			.SO(gen[3715]),
			.S(gen[3716]),
			.SE(gen[3717]),

			.SELF(gen[3621]),
			.cell_state(gen[3621])
		); 

/******************* CELL 3622 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3622 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3526]),
			.N(gen[3527]),
			.NE(gen[3528]),

			.O(gen[3621]),
			.E(gen[3623]),

			.SO(gen[3716]),
			.S(gen[3717]),
			.SE(gen[3718]),

			.SELF(gen[3622]),
			.cell_state(gen[3622])
		); 

/******************* CELL 3623 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3623 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3527]),
			.N(gen[3528]),
			.NE(gen[3529]),

			.O(gen[3622]),
			.E(gen[3624]),

			.SO(gen[3717]),
			.S(gen[3718]),
			.SE(gen[3719]),

			.SELF(gen[3623]),
			.cell_state(gen[3623])
		); 

/******************* CELL 3624 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3624 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3528]),
			.N(gen[3529]),
			.NE(gen[3530]),

			.O(gen[3623]),
			.E(gen[3625]),

			.SO(gen[3718]),
			.S(gen[3719]),
			.SE(gen[3720]),

			.SELF(gen[3624]),
			.cell_state(gen[3624])
		); 

/******************* CELL 3625 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3625 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3529]),
			.N(gen[3530]),
			.NE(gen[3531]),

			.O(gen[3624]),
			.E(gen[3626]),

			.SO(gen[3719]),
			.S(gen[3720]),
			.SE(gen[3721]),

			.SELF(gen[3625]),
			.cell_state(gen[3625])
		); 

/******************* CELL 3626 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3626 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3530]),
			.N(gen[3531]),
			.NE(gen[3532]),

			.O(gen[3625]),
			.E(gen[3627]),

			.SO(gen[3720]),
			.S(gen[3721]),
			.SE(gen[3722]),

			.SELF(gen[3626]),
			.cell_state(gen[3626])
		); 

/******************* CELL 3627 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3627 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3531]),
			.N(gen[3532]),
			.NE(gen[3533]),

			.O(gen[3626]),
			.E(gen[3628]),

			.SO(gen[3721]),
			.S(gen[3722]),
			.SE(gen[3723]),

			.SELF(gen[3627]),
			.cell_state(gen[3627])
		); 

/******************* CELL 3628 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3628 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3532]),
			.N(gen[3533]),
			.NE(gen[3534]),

			.O(gen[3627]),
			.E(gen[3629]),

			.SO(gen[3722]),
			.S(gen[3723]),
			.SE(gen[3724]),

			.SELF(gen[3628]),
			.cell_state(gen[3628])
		); 

/******************* CELL 3629 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3629 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3533]),
			.N(gen[3534]),
			.NE(gen[3535]),

			.O(gen[3628]),
			.E(gen[3630]),

			.SO(gen[3723]),
			.S(gen[3724]),
			.SE(gen[3725]),

			.SELF(gen[3629]),
			.cell_state(gen[3629])
		); 

/******************* CELL 3630 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3630 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3534]),
			.N(gen[3535]),
			.NE(gen[3536]),

			.O(gen[3629]),
			.E(gen[3631]),

			.SO(gen[3724]),
			.S(gen[3725]),
			.SE(gen[3726]),

			.SELF(gen[3630]),
			.cell_state(gen[3630])
		); 

/******************* CELL 3631 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3631 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3535]),
			.N(gen[3536]),
			.NE(gen[3537]),

			.O(gen[3630]),
			.E(gen[3632]),

			.SO(gen[3725]),
			.S(gen[3726]),
			.SE(gen[3727]),

			.SELF(gen[3631]),
			.cell_state(gen[3631])
		); 

/******************* CELL 3632 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3632 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3536]),
			.N(gen[3537]),
			.NE(gen[3538]),

			.O(gen[3631]),
			.E(gen[3633]),

			.SO(gen[3726]),
			.S(gen[3727]),
			.SE(gen[3728]),

			.SELF(gen[3632]),
			.cell_state(gen[3632])
		); 

/******************* CELL 3633 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3633 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3537]),
			.N(gen[3538]),
			.NE(gen[3539]),

			.O(gen[3632]),
			.E(gen[3634]),

			.SO(gen[3727]),
			.S(gen[3728]),
			.SE(gen[3729]),

			.SELF(gen[3633]),
			.cell_state(gen[3633])
		); 

/******************* CELL 3634 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3634 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3538]),
			.N(gen[3539]),
			.NE(gen[3540]),

			.O(gen[3633]),
			.E(gen[3635]),

			.SO(gen[3728]),
			.S(gen[3729]),
			.SE(gen[3730]),

			.SELF(gen[3634]),
			.cell_state(gen[3634])
		); 

/******************* CELL 3635 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3635 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3539]),
			.N(gen[3540]),
			.NE(gen[3541]),

			.O(gen[3634]),
			.E(gen[3636]),

			.SO(gen[3729]),
			.S(gen[3730]),
			.SE(gen[3731]),

			.SELF(gen[3635]),
			.cell_state(gen[3635])
		); 

/******************* CELL 3636 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3636 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3540]),
			.N(gen[3541]),
			.NE(gen[3542]),

			.O(gen[3635]),
			.E(gen[3637]),

			.SO(gen[3730]),
			.S(gen[3731]),
			.SE(gen[3732]),

			.SELF(gen[3636]),
			.cell_state(gen[3636])
		); 

/******************* CELL 3637 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3637 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3541]),
			.N(gen[3542]),
			.NE(gen[3543]),

			.O(gen[3636]),
			.E(gen[3638]),

			.SO(gen[3731]),
			.S(gen[3732]),
			.SE(gen[3733]),

			.SELF(gen[3637]),
			.cell_state(gen[3637])
		); 

/******************* CELL 3638 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3638 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3542]),
			.N(gen[3543]),
			.NE(gen[3544]),

			.O(gen[3637]),
			.E(gen[3639]),

			.SO(gen[3732]),
			.S(gen[3733]),
			.SE(gen[3734]),

			.SELF(gen[3638]),
			.cell_state(gen[3638])
		); 

/******************* CELL 3639 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3639 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3543]),
			.N(gen[3544]),
			.NE(gen[3545]),

			.O(gen[3638]),
			.E(gen[3640]),

			.SO(gen[3733]),
			.S(gen[3734]),
			.SE(gen[3735]),

			.SELF(gen[3639]),
			.cell_state(gen[3639])
		); 

/******************* CELL 3640 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3640 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3544]),
			.N(gen[3545]),
			.NE(gen[3546]),

			.O(gen[3639]),
			.E(gen[3641]),

			.SO(gen[3734]),
			.S(gen[3735]),
			.SE(gen[3736]),

			.SELF(gen[3640]),
			.cell_state(gen[3640])
		); 

/******************* CELL 3641 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3641 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3545]),
			.N(gen[3546]),
			.NE(gen[3547]),

			.O(gen[3640]),
			.E(gen[3642]),

			.SO(gen[3735]),
			.S(gen[3736]),
			.SE(gen[3737]),

			.SELF(gen[3641]),
			.cell_state(gen[3641])
		); 

/******************* CELL 3642 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3642 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3546]),
			.N(gen[3547]),
			.NE(gen[3548]),

			.O(gen[3641]),
			.E(gen[3643]),

			.SO(gen[3736]),
			.S(gen[3737]),
			.SE(gen[3738]),

			.SELF(gen[3642]),
			.cell_state(gen[3642])
		); 

/******************* CELL 3643 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3643 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3547]),
			.N(gen[3548]),
			.NE(gen[3549]),

			.O(gen[3642]),
			.E(gen[3644]),

			.SO(gen[3737]),
			.S(gen[3738]),
			.SE(gen[3739]),

			.SELF(gen[3643]),
			.cell_state(gen[3643])
		); 

/******************* CELL 3644 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3644 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3548]),
			.N(gen[3549]),
			.NE(gen[3550]),

			.O(gen[3643]),
			.E(gen[3645]),

			.SO(gen[3738]),
			.S(gen[3739]),
			.SE(gen[3740]),

			.SELF(gen[3644]),
			.cell_state(gen[3644])
		); 

/******************* CELL 3645 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3645 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3549]),
			.N(gen[3550]),
			.NE(gen[3551]),

			.O(gen[3644]),
			.E(gen[3646]),

			.SO(gen[3739]),
			.S(gen[3740]),
			.SE(gen[3741]),

			.SELF(gen[3645]),
			.cell_state(gen[3645])
		); 

/******************* CELL 3646 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3646 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3550]),
			.N(gen[3551]),
			.NE(gen[3552]),

			.O(gen[3645]),
			.E(gen[3647]),

			.SO(gen[3740]),
			.S(gen[3741]),
			.SE(gen[3742]),

			.SELF(gen[3646]),
			.cell_state(gen[3646])
		); 

/******************* CELL 3647 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3647 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3551]),
			.N(gen[3552]),
			.NE(gen[3553]),

			.O(gen[3646]),
			.E(gen[3648]),

			.SO(gen[3741]),
			.S(gen[3742]),
			.SE(gen[3743]),

			.SELF(gen[3647]),
			.cell_state(gen[3647])
		); 

/******************* CELL 3648 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3648 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3552]),
			.N(gen[3553]),
			.NE(gen[3554]),

			.O(gen[3647]),
			.E(gen[3649]),

			.SO(gen[3742]),
			.S(gen[3743]),
			.SE(gen[3744]),

			.SELF(gen[3648]),
			.cell_state(gen[3648])
		); 

/******************* CELL 3649 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3649 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3553]),
			.N(gen[3554]),
			.NE(gen[3555]),

			.O(gen[3648]),
			.E(gen[3650]),

			.SO(gen[3743]),
			.S(gen[3744]),
			.SE(gen[3745]),

			.SELF(gen[3649]),
			.cell_state(gen[3649])
		); 

/******************* CELL 3650 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3650 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3554]),
			.N(gen[3555]),
			.NE(gen[3556]),

			.O(gen[3649]),
			.E(gen[3651]),

			.SO(gen[3744]),
			.S(gen[3745]),
			.SE(gen[3746]),

			.SELF(gen[3650]),
			.cell_state(gen[3650])
		); 

/******************* CELL 3651 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3651 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3555]),
			.N(gen[3556]),
			.NE(gen[3557]),

			.O(gen[3650]),
			.E(gen[3652]),

			.SO(gen[3745]),
			.S(gen[3746]),
			.SE(gen[3747]),

			.SELF(gen[3651]),
			.cell_state(gen[3651])
		); 

/******************* CELL 3652 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3652 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3556]),
			.N(gen[3557]),
			.NE(gen[3558]),

			.O(gen[3651]),
			.E(gen[3653]),

			.SO(gen[3746]),
			.S(gen[3747]),
			.SE(gen[3748]),

			.SELF(gen[3652]),
			.cell_state(gen[3652])
		); 

/******************* CELL 3653 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3653 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3557]),
			.N(gen[3558]),
			.NE(gen[3559]),

			.O(gen[3652]),
			.E(gen[3654]),

			.SO(gen[3747]),
			.S(gen[3748]),
			.SE(gen[3749]),

			.SELF(gen[3653]),
			.cell_state(gen[3653])
		); 

/******************* CELL 3654 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3654 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3558]),
			.N(gen[3559]),
			.NE(gen[3560]),

			.O(gen[3653]),
			.E(gen[3655]),

			.SO(gen[3748]),
			.S(gen[3749]),
			.SE(gen[3750]),

			.SELF(gen[3654]),
			.cell_state(gen[3654])
		); 

/******************* CELL 3655 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3655 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3559]),
			.N(gen[3560]),
			.NE(gen[3561]),

			.O(gen[3654]),
			.E(gen[3656]),

			.SO(gen[3749]),
			.S(gen[3750]),
			.SE(gen[3751]),

			.SELF(gen[3655]),
			.cell_state(gen[3655])
		); 

/******************* CELL 3656 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3656 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3560]),
			.N(gen[3561]),
			.NE(gen[3562]),

			.O(gen[3655]),
			.E(gen[3657]),

			.SO(gen[3750]),
			.S(gen[3751]),
			.SE(gen[3752]),

			.SELF(gen[3656]),
			.cell_state(gen[3656])
		); 

/******************* CELL 3657 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3657 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3561]),
			.N(gen[3562]),
			.NE(gen[3563]),

			.O(gen[3656]),
			.E(gen[3658]),

			.SO(gen[3751]),
			.S(gen[3752]),
			.SE(gen[3753]),

			.SELF(gen[3657]),
			.cell_state(gen[3657])
		); 

/******************* CELL 3658 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3658 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3562]),
			.N(gen[3563]),
			.NE(gen[3564]),

			.O(gen[3657]),
			.E(gen[3659]),

			.SO(gen[3752]),
			.S(gen[3753]),
			.SE(gen[3754]),

			.SELF(gen[3658]),
			.cell_state(gen[3658])
		); 

/******************* CELL 3659 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3659 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3563]),
			.N(gen[3564]),
			.NE(gen[3565]),

			.O(gen[3658]),
			.E(gen[3660]),

			.SO(gen[3753]),
			.S(gen[3754]),
			.SE(gen[3755]),

			.SELF(gen[3659]),
			.cell_state(gen[3659])
		); 

/******************* CELL 3660 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3660 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3564]),
			.N(gen[3565]),
			.NE(gen[3566]),

			.O(gen[3659]),
			.E(gen[3661]),

			.SO(gen[3754]),
			.S(gen[3755]),
			.SE(gen[3756]),

			.SELF(gen[3660]),
			.cell_state(gen[3660])
		); 

/******************* CELL 3661 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3661 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3565]),
			.N(gen[3566]),
			.NE(gen[3567]),

			.O(gen[3660]),
			.E(gen[3662]),

			.SO(gen[3755]),
			.S(gen[3756]),
			.SE(gen[3757]),

			.SELF(gen[3661]),
			.cell_state(gen[3661])
		); 

/******************* CELL 3662 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3662 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3566]),
			.N(gen[3567]),
			.NE(gen[3568]),

			.O(gen[3661]),
			.E(gen[3663]),

			.SO(gen[3756]),
			.S(gen[3757]),
			.SE(gen[3758]),

			.SELF(gen[3662]),
			.cell_state(gen[3662])
		); 

/******************* CELL 3663 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3663 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3567]),
			.N(gen[3568]),
			.NE(gen[3569]),

			.O(gen[3662]),
			.E(gen[3664]),

			.SO(gen[3757]),
			.S(gen[3758]),
			.SE(gen[3759]),

			.SELF(gen[3663]),
			.cell_state(gen[3663])
		); 

/******************* CELL 3664 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3664 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3568]),
			.N(gen[3569]),
			.NE(gen[3570]),

			.O(gen[3663]),
			.E(gen[3665]),

			.SO(gen[3758]),
			.S(gen[3759]),
			.SE(gen[3760]),

			.SELF(gen[3664]),
			.cell_state(gen[3664])
		); 

/******************* CELL 3665 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3665 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3569]),
			.N(gen[3570]),
			.NE(gen[3571]),

			.O(gen[3664]),
			.E(gen[3666]),

			.SO(gen[3759]),
			.S(gen[3760]),
			.SE(gen[3761]),

			.SELF(gen[3665]),
			.cell_state(gen[3665])
		); 

/******************* CELL 3666 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3666 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3570]),
			.N(gen[3571]),
			.NE(gen[3572]),

			.O(gen[3665]),
			.E(gen[3667]),

			.SO(gen[3760]),
			.S(gen[3761]),
			.SE(gen[3762]),

			.SELF(gen[3666]),
			.cell_state(gen[3666])
		); 

/******************* CELL 3667 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3667 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3571]),
			.N(gen[3572]),
			.NE(gen[3573]),

			.O(gen[3666]),
			.E(gen[3668]),

			.SO(gen[3761]),
			.S(gen[3762]),
			.SE(gen[3763]),

			.SELF(gen[3667]),
			.cell_state(gen[3667])
		); 

/******************* CELL 3668 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3668 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3572]),
			.N(gen[3573]),
			.NE(gen[3574]),

			.O(gen[3667]),
			.E(gen[3669]),

			.SO(gen[3762]),
			.S(gen[3763]),
			.SE(gen[3764]),

			.SELF(gen[3668]),
			.cell_state(gen[3668])
		); 

/******************* CELL 3669 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3669 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3573]),
			.N(gen[3574]),
			.NE(gen[3575]),

			.O(gen[3668]),
			.E(gen[3670]),

			.SO(gen[3763]),
			.S(gen[3764]),
			.SE(gen[3765]),

			.SELF(gen[3669]),
			.cell_state(gen[3669])
		); 

/******************* CELL 3670 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3670 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3574]),
			.N(gen[3575]),
			.NE(gen[3576]),

			.O(gen[3669]),
			.E(gen[3671]),

			.SO(gen[3764]),
			.S(gen[3765]),
			.SE(gen[3766]),

			.SELF(gen[3670]),
			.cell_state(gen[3670])
		); 

/******************* CELL 3671 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3671 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3575]),
			.N(gen[3576]),
			.NE(gen[3577]),

			.O(gen[3670]),
			.E(gen[3672]),

			.SO(gen[3765]),
			.S(gen[3766]),
			.SE(gen[3767]),

			.SELF(gen[3671]),
			.cell_state(gen[3671])
		); 

/******************* CELL 3672 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3672 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3576]),
			.N(gen[3577]),
			.NE(gen[3578]),

			.O(gen[3671]),
			.E(gen[3673]),

			.SO(gen[3766]),
			.S(gen[3767]),
			.SE(gen[3768]),

			.SELF(gen[3672]),
			.cell_state(gen[3672])
		); 

/******************* CELL 3673 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3673 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3577]),
			.N(gen[3578]),
			.NE(gen[3579]),

			.O(gen[3672]),
			.E(gen[3674]),

			.SO(gen[3767]),
			.S(gen[3768]),
			.SE(gen[3769]),

			.SELF(gen[3673]),
			.cell_state(gen[3673])
		); 

/******************* CELL 3674 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3674 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3578]),
			.N(gen[3579]),
			.NE(gen[3580]),

			.O(gen[3673]),
			.E(gen[3675]),

			.SO(gen[3768]),
			.S(gen[3769]),
			.SE(gen[3770]),

			.SELF(gen[3674]),
			.cell_state(gen[3674])
		); 

/******************* CELL 3675 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3675 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3579]),
			.N(gen[3580]),
			.NE(gen[3581]),

			.O(gen[3674]),
			.E(gen[3676]),

			.SO(gen[3769]),
			.S(gen[3770]),
			.SE(gen[3771]),

			.SELF(gen[3675]),
			.cell_state(gen[3675])
		); 

/******************* CELL 3676 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3676 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3580]),
			.N(gen[3581]),
			.NE(gen[3582]),

			.O(gen[3675]),
			.E(gen[3677]),

			.SO(gen[3770]),
			.S(gen[3771]),
			.SE(gen[3772]),

			.SELF(gen[3676]),
			.cell_state(gen[3676])
		); 

/******************* CELL 3677 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3677 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3581]),
			.N(gen[3582]),
			.NE(gen[3583]),

			.O(gen[3676]),
			.E(gen[3678]),

			.SO(gen[3771]),
			.S(gen[3772]),
			.SE(gen[3773]),

			.SELF(gen[3677]),
			.cell_state(gen[3677])
		); 

/******************* CELL 3678 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3678 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3582]),
			.N(gen[3583]),
			.NE(gen[3584]),

			.O(gen[3677]),
			.E(gen[3679]),

			.SO(gen[3772]),
			.S(gen[3773]),
			.SE(gen[3774]),

			.SELF(gen[3678]),
			.cell_state(gen[3678])
		); 

/******************* CELL 3679 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3679 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3583]),
			.N(gen[3584]),
			.NE(gen[3585]),

			.O(gen[3678]),
			.E(gen[3680]),

			.SO(gen[3773]),
			.S(gen[3774]),
			.SE(gen[3775]),

			.SELF(gen[3679]),
			.cell_state(gen[3679])
		); 

/******************* CELL 3680 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3680 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3584]),
			.N(gen[3585]),
			.NE(gen[3586]),

			.O(gen[3679]),
			.E(gen[3681]),

			.SO(gen[3774]),
			.S(gen[3775]),
			.SE(gen[3776]),

			.SELF(gen[3680]),
			.cell_state(gen[3680])
		); 

/******************* CELL 3681 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3681 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3585]),
			.N(gen[3586]),
			.NE(gen[3587]),

			.O(gen[3680]),
			.E(gen[3682]),

			.SO(gen[3775]),
			.S(gen[3776]),
			.SE(gen[3777]),

			.SELF(gen[3681]),
			.cell_state(gen[3681])
		); 

/******************* CELL 3682 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3682 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3586]),
			.N(gen[3587]),
			.NE(gen[3588]),

			.O(gen[3681]),
			.E(gen[3683]),

			.SO(gen[3776]),
			.S(gen[3777]),
			.SE(gen[3778]),

			.SELF(gen[3682]),
			.cell_state(gen[3682])
		); 

/******************* CELL 3683 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3683 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3587]),
			.N(gen[3588]),
			.NE(gen[3589]),

			.O(gen[3682]),
			.E(gen[3684]),

			.SO(gen[3777]),
			.S(gen[3778]),
			.SE(gen[3779]),

			.SELF(gen[3683]),
			.cell_state(gen[3683])
		); 

/******************* CELL 3684 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3684 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3588]),
			.N(gen[3589]),
			.NE(gen[3590]),

			.O(gen[3683]),
			.E(gen[3685]),

			.SO(gen[3778]),
			.S(gen[3779]),
			.SE(gen[3780]),

			.SELF(gen[3684]),
			.cell_state(gen[3684])
		); 

/******************* CELL 3685 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3685 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3589]),
			.N(gen[3590]),
			.NE(gen[3591]),

			.O(gen[3684]),
			.E(gen[3686]),

			.SO(gen[3779]),
			.S(gen[3780]),
			.SE(gen[3781]),

			.SELF(gen[3685]),
			.cell_state(gen[3685])
		); 

/******************* CELL 3686 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3686 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3590]),
			.N(gen[3591]),
			.NE(gen[3592]),

			.O(gen[3685]),
			.E(gen[3687]),

			.SO(gen[3780]),
			.S(gen[3781]),
			.SE(gen[3782]),

			.SELF(gen[3686]),
			.cell_state(gen[3686])
		); 

/******************* CELL 3687 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3687 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3591]),
			.N(gen[3592]),
			.NE(gen[3593]),

			.O(gen[3686]),
			.E(gen[3688]),

			.SO(gen[3781]),
			.S(gen[3782]),
			.SE(gen[3783]),

			.SELF(gen[3687]),
			.cell_state(gen[3687])
		); 

/******************* CELL 3688 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3688 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3592]),
			.N(gen[3593]),
			.NE(gen[3594]),

			.O(gen[3687]),
			.E(gen[3689]),

			.SO(gen[3782]),
			.S(gen[3783]),
			.SE(gen[3784]),

			.SELF(gen[3688]),
			.cell_state(gen[3688])
		); 

/******************* CELL 3689 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3689 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3593]),
			.N(gen[3594]),
			.NE(gen[3595]),

			.O(gen[3688]),
			.E(gen[3690]),

			.SO(gen[3783]),
			.S(gen[3784]),
			.SE(gen[3785]),

			.SELF(gen[3689]),
			.cell_state(gen[3689])
		); 

/******************* CELL 3690 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3690 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3594]),
			.N(gen[3595]),
			.NE(gen[3596]),

			.O(gen[3689]),
			.E(gen[3691]),

			.SO(gen[3784]),
			.S(gen[3785]),
			.SE(gen[3786]),

			.SELF(gen[3690]),
			.cell_state(gen[3690])
		); 

/******************* CELL 3691 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3691 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3595]),
			.N(gen[3596]),
			.NE(gen[3597]),

			.O(gen[3690]),
			.E(gen[3692]),

			.SO(gen[3785]),
			.S(gen[3786]),
			.SE(gen[3787]),

			.SELF(gen[3691]),
			.cell_state(gen[3691])
		); 

/******************* CELL 3692 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3692 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3596]),
			.N(gen[3597]),
			.NE(gen[3598]),

			.O(gen[3691]),
			.E(gen[3693]),

			.SO(gen[3786]),
			.S(gen[3787]),
			.SE(gen[3788]),

			.SELF(gen[3692]),
			.cell_state(gen[3692])
		); 

/******************* CELL 3693 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3693 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3597]),
			.N(gen[3598]),
			.NE(gen[3599]),

			.O(gen[3692]),
			.E(gen[3694]),

			.SO(gen[3787]),
			.S(gen[3788]),
			.SE(gen[3789]),

			.SELF(gen[3693]),
			.cell_state(gen[3693])
		); 

/******************* CELL 3694 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3694 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3598]),
			.N(gen[3599]),
			.NE(gen[3600]),

			.O(gen[3693]),
			.E(gen[3695]),

			.SO(gen[3788]),
			.S(gen[3789]),
			.SE(gen[3790]),

			.SELF(gen[3694]),
			.cell_state(gen[3694])
		); 

/******************* CELL 3695 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3695 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3599]),
			.N(gen[3600]),
			.NE(gen[3601]),

			.O(gen[3694]),
			.E(gen[3696]),

			.SO(gen[3789]),
			.S(gen[3790]),
			.SE(gen[3791]),

			.SELF(gen[3695]),
			.cell_state(gen[3695])
		); 

/******************* CELL 3696 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3696 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3600]),
			.N(gen[3601]),
			.NE(gen[3602]),

			.O(gen[3695]),
			.E(gen[3697]),

			.SO(gen[3790]),
			.S(gen[3791]),
			.SE(gen[3792]),

			.SELF(gen[3696]),
			.cell_state(gen[3696])
		); 

/******************* CELL 3697 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3697 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3601]),
			.N(gen[3602]),
			.NE(gen[3603]),

			.O(gen[3696]),
			.E(gen[3698]),

			.SO(gen[3791]),
			.S(gen[3792]),
			.SE(gen[3793]),

			.SELF(gen[3697]),
			.cell_state(gen[3697])
		); 

/******************* CELL 3698 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3698 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3602]),
			.N(gen[3603]),
			.NE(gen[3604]),

			.O(gen[3697]),
			.E(gen[3699]),

			.SO(gen[3792]),
			.S(gen[3793]),
			.SE(gen[3794]),

			.SELF(gen[3698]),
			.cell_state(gen[3698])
		); 

/******************* CELL 3699 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3699 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3603]),
			.N(gen[3604]),
			.NE(gen[3605]),

			.O(gen[3698]),
			.E(gen[3700]),

			.SO(gen[3793]),
			.S(gen[3794]),
			.SE(gen[3795]),

			.SELF(gen[3699]),
			.cell_state(gen[3699])
		); 

/******************* CELL 3700 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3700 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3604]),
			.N(gen[3605]),
			.NE(gen[3606]),

			.O(gen[3699]),
			.E(gen[3701]),

			.SO(gen[3794]),
			.S(gen[3795]),
			.SE(gen[3796]),

			.SELF(gen[3700]),
			.cell_state(gen[3700])
		); 

/******************* CELL 3701 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3701 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3605]),
			.N(gen[3606]),
			.NE(gen[3607]),

			.O(gen[3700]),
			.E(gen[3702]),

			.SO(gen[3795]),
			.S(gen[3796]),
			.SE(gen[3797]),

			.SELF(gen[3701]),
			.cell_state(gen[3701])
		); 

/******************* CELL 3702 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3702 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3606]),
			.N(gen[3607]),
			.NE(gen[3608]),

			.O(gen[3701]),
			.E(gen[3703]),

			.SO(gen[3796]),
			.S(gen[3797]),
			.SE(gen[3798]),

			.SELF(gen[3702]),
			.cell_state(gen[3702])
		); 

/******************* CELL 3703 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3703 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3607]),
			.N(gen[3608]),
			.NE(gen[3609]),

			.O(gen[3702]),
			.E(gen[3704]),

			.SO(gen[3797]),
			.S(gen[3798]),
			.SE(gen[3799]),

			.SELF(gen[3703]),
			.cell_state(gen[3703])
		); 

/******************* CELL 3704 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3704 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3608]),
			.N(gen[3609]),
			.NE(gen[3608]),

			.O(gen[3703]),
			.E(gen[3703]),

			.SO(gen[3798]),
			.S(gen[3799]),
			.SE(gen[3798]),

			.SELF(gen[3704]),
			.cell_state(gen[3704])
		); 

/******************* CELL 3705 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3705 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3611]),
			.N(gen[3610]),
			.NE(gen[3611]),

			.O(gen[3706]),
			.E(gen[3706]),

			.SO(gen[3801]),
			.S(gen[3800]),
			.SE(gen[3801]),

			.SELF(gen[3705]),
			.cell_state(gen[3705])
		); 

/******************* CELL 3706 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3706 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3610]),
			.N(gen[3611]),
			.NE(gen[3612]),

			.O(gen[3705]),
			.E(gen[3707]),

			.SO(gen[3800]),
			.S(gen[3801]),
			.SE(gen[3802]),

			.SELF(gen[3706]),
			.cell_state(gen[3706])
		); 

/******************* CELL 3707 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3707 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3611]),
			.N(gen[3612]),
			.NE(gen[3613]),

			.O(gen[3706]),
			.E(gen[3708]),

			.SO(gen[3801]),
			.S(gen[3802]),
			.SE(gen[3803]),

			.SELF(gen[3707]),
			.cell_state(gen[3707])
		); 

/******************* CELL 3708 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3708 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3612]),
			.N(gen[3613]),
			.NE(gen[3614]),

			.O(gen[3707]),
			.E(gen[3709]),

			.SO(gen[3802]),
			.S(gen[3803]),
			.SE(gen[3804]),

			.SELF(gen[3708]),
			.cell_state(gen[3708])
		); 

/******************* CELL 3709 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3709 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3613]),
			.N(gen[3614]),
			.NE(gen[3615]),

			.O(gen[3708]),
			.E(gen[3710]),

			.SO(gen[3803]),
			.S(gen[3804]),
			.SE(gen[3805]),

			.SELF(gen[3709]),
			.cell_state(gen[3709])
		); 

/******************* CELL 3710 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3710 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3614]),
			.N(gen[3615]),
			.NE(gen[3616]),

			.O(gen[3709]),
			.E(gen[3711]),

			.SO(gen[3804]),
			.S(gen[3805]),
			.SE(gen[3806]),

			.SELF(gen[3710]),
			.cell_state(gen[3710])
		); 

/******************* CELL 3711 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3711 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3615]),
			.N(gen[3616]),
			.NE(gen[3617]),

			.O(gen[3710]),
			.E(gen[3712]),

			.SO(gen[3805]),
			.S(gen[3806]),
			.SE(gen[3807]),

			.SELF(gen[3711]),
			.cell_state(gen[3711])
		); 

/******************* CELL 3712 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3712 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3616]),
			.N(gen[3617]),
			.NE(gen[3618]),

			.O(gen[3711]),
			.E(gen[3713]),

			.SO(gen[3806]),
			.S(gen[3807]),
			.SE(gen[3808]),

			.SELF(gen[3712]),
			.cell_state(gen[3712])
		); 

/******************* CELL 3713 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3713 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3617]),
			.N(gen[3618]),
			.NE(gen[3619]),

			.O(gen[3712]),
			.E(gen[3714]),

			.SO(gen[3807]),
			.S(gen[3808]),
			.SE(gen[3809]),

			.SELF(gen[3713]),
			.cell_state(gen[3713])
		); 

/******************* CELL 3714 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3714 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3618]),
			.N(gen[3619]),
			.NE(gen[3620]),

			.O(gen[3713]),
			.E(gen[3715]),

			.SO(gen[3808]),
			.S(gen[3809]),
			.SE(gen[3810]),

			.SELF(gen[3714]),
			.cell_state(gen[3714])
		); 

/******************* CELL 3715 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3715 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3619]),
			.N(gen[3620]),
			.NE(gen[3621]),

			.O(gen[3714]),
			.E(gen[3716]),

			.SO(gen[3809]),
			.S(gen[3810]),
			.SE(gen[3811]),

			.SELF(gen[3715]),
			.cell_state(gen[3715])
		); 

/******************* CELL 3716 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3716 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3620]),
			.N(gen[3621]),
			.NE(gen[3622]),

			.O(gen[3715]),
			.E(gen[3717]),

			.SO(gen[3810]),
			.S(gen[3811]),
			.SE(gen[3812]),

			.SELF(gen[3716]),
			.cell_state(gen[3716])
		); 

/******************* CELL 3717 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3717 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3621]),
			.N(gen[3622]),
			.NE(gen[3623]),

			.O(gen[3716]),
			.E(gen[3718]),

			.SO(gen[3811]),
			.S(gen[3812]),
			.SE(gen[3813]),

			.SELF(gen[3717]),
			.cell_state(gen[3717])
		); 

/******************* CELL 3718 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3718 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3622]),
			.N(gen[3623]),
			.NE(gen[3624]),

			.O(gen[3717]),
			.E(gen[3719]),

			.SO(gen[3812]),
			.S(gen[3813]),
			.SE(gen[3814]),

			.SELF(gen[3718]),
			.cell_state(gen[3718])
		); 

/******************* CELL 3719 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3719 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3623]),
			.N(gen[3624]),
			.NE(gen[3625]),

			.O(gen[3718]),
			.E(gen[3720]),

			.SO(gen[3813]),
			.S(gen[3814]),
			.SE(gen[3815]),

			.SELF(gen[3719]),
			.cell_state(gen[3719])
		); 

/******************* CELL 3720 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3720 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3624]),
			.N(gen[3625]),
			.NE(gen[3626]),

			.O(gen[3719]),
			.E(gen[3721]),

			.SO(gen[3814]),
			.S(gen[3815]),
			.SE(gen[3816]),

			.SELF(gen[3720]),
			.cell_state(gen[3720])
		); 

/******************* CELL 3721 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3721 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3625]),
			.N(gen[3626]),
			.NE(gen[3627]),

			.O(gen[3720]),
			.E(gen[3722]),

			.SO(gen[3815]),
			.S(gen[3816]),
			.SE(gen[3817]),

			.SELF(gen[3721]),
			.cell_state(gen[3721])
		); 

/******************* CELL 3722 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3722 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3626]),
			.N(gen[3627]),
			.NE(gen[3628]),

			.O(gen[3721]),
			.E(gen[3723]),

			.SO(gen[3816]),
			.S(gen[3817]),
			.SE(gen[3818]),

			.SELF(gen[3722]),
			.cell_state(gen[3722])
		); 

/******************* CELL 3723 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3723 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3627]),
			.N(gen[3628]),
			.NE(gen[3629]),

			.O(gen[3722]),
			.E(gen[3724]),

			.SO(gen[3817]),
			.S(gen[3818]),
			.SE(gen[3819]),

			.SELF(gen[3723]),
			.cell_state(gen[3723])
		); 

/******************* CELL 3724 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3724 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3628]),
			.N(gen[3629]),
			.NE(gen[3630]),

			.O(gen[3723]),
			.E(gen[3725]),

			.SO(gen[3818]),
			.S(gen[3819]),
			.SE(gen[3820]),

			.SELF(gen[3724]),
			.cell_state(gen[3724])
		); 

/******************* CELL 3725 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3725 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3629]),
			.N(gen[3630]),
			.NE(gen[3631]),

			.O(gen[3724]),
			.E(gen[3726]),

			.SO(gen[3819]),
			.S(gen[3820]),
			.SE(gen[3821]),

			.SELF(gen[3725]),
			.cell_state(gen[3725])
		); 

/******************* CELL 3726 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3726 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3630]),
			.N(gen[3631]),
			.NE(gen[3632]),

			.O(gen[3725]),
			.E(gen[3727]),

			.SO(gen[3820]),
			.S(gen[3821]),
			.SE(gen[3822]),

			.SELF(gen[3726]),
			.cell_state(gen[3726])
		); 

/******************* CELL 3727 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3727 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3631]),
			.N(gen[3632]),
			.NE(gen[3633]),

			.O(gen[3726]),
			.E(gen[3728]),

			.SO(gen[3821]),
			.S(gen[3822]),
			.SE(gen[3823]),

			.SELF(gen[3727]),
			.cell_state(gen[3727])
		); 

/******************* CELL 3728 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3728 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3632]),
			.N(gen[3633]),
			.NE(gen[3634]),

			.O(gen[3727]),
			.E(gen[3729]),

			.SO(gen[3822]),
			.S(gen[3823]),
			.SE(gen[3824]),

			.SELF(gen[3728]),
			.cell_state(gen[3728])
		); 

/******************* CELL 3729 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3729 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3633]),
			.N(gen[3634]),
			.NE(gen[3635]),

			.O(gen[3728]),
			.E(gen[3730]),

			.SO(gen[3823]),
			.S(gen[3824]),
			.SE(gen[3825]),

			.SELF(gen[3729]),
			.cell_state(gen[3729])
		); 

/******************* CELL 3730 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3730 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3634]),
			.N(gen[3635]),
			.NE(gen[3636]),

			.O(gen[3729]),
			.E(gen[3731]),

			.SO(gen[3824]),
			.S(gen[3825]),
			.SE(gen[3826]),

			.SELF(gen[3730]),
			.cell_state(gen[3730])
		); 

/******************* CELL 3731 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3731 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3635]),
			.N(gen[3636]),
			.NE(gen[3637]),

			.O(gen[3730]),
			.E(gen[3732]),

			.SO(gen[3825]),
			.S(gen[3826]),
			.SE(gen[3827]),

			.SELF(gen[3731]),
			.cell_state(gen[3731])
		); 

/******************* CELL 3732 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3732 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3636]),
			.N(gen[3637]),
			.NE(gen[3638]),

			.O(gen[3731]),
			.E(gen[3733]),

			.SO(gen[3826]),
			.S(gen[3827]),
			.SE(gen[3828]),

			.SELF(gen[3732]),
			.cell_state(gen[3732])
		); 

/******************* CELL 3733 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3733 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3637]),
			.N(gen[3638]),
			.NE(gen[3639]),

			.O(gen[3732]),
			.E(gen[3734]),

			.SO(gen[3827]),
			.S(gen[3828]),
			.SE(gen[3829]),

			.SELF(gen[3733]),
			.cell_state(gen[3733])
		); 

/******************* CELL 3734 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3734 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3638]),
			.N(gen[3639]),
			.NE(gen[3640]),

			.O(gen[3733]),
			.E(gen[3735]),

			.SO(gen[3828]),
			.S(gen[3829]),
			.SE(gen[3830]),

			.SELF(gen[3734]),
			.cell_state(gen[3734])
		); 

/******************* CELL 3735 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3735 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3639]),
			.N(gen[3640]),
			.NE(gen[3641]),

			.O(gen[3734]),
			.E(gen[3736]),

			.SO(gen[3829]),
			.S(gen[3830]),
			.SE(gen[3831]),

			.SELF(gen[3735]),
			.cell_state(gen[3735])
		); 

/******************* CELL 3736 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3736 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3640]),
			.N(gen[3641]),
			.NE(gen[3642]),

			.O(gen[3735]),
			.E(gen[3737]),

			.SO(gen[3830]),
			.S(gen[3831]),
			.SE(gen[3832]),

			.SELF(gen[3736]),
			.cell_state(gen[3736])
		); 

/******************* CELL 3737 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3737 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3641]),
			.N(gen[3642]),
			.NE(gen[3643]),

			.O(gen[3736]),
			.E(gen[3738]),

			.SO(gen[3831]),
			.S(gen[3832]),
			.SE(gen[3833]),

			.SELF(gen[3737]),
			.cell_state(gen[3737])
		); 

/******************* CELL 3738 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3738 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3642]),
			.N(gen[3643]),
			.NE(gen[3644]),

			.O(gen[3737]),
			.E(gen[3739]),

			.SO(gen[3832]),
			.S(gen[3833]),
			.SE(gen[3834]),

			.SELF(gen[3738]),
			.cell_state(gen[3738])
		); 

/******************* CELL 3739 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3739 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3643]),
			.N(gen[3644]),
			.NE(gen[3645]),

			.O(gen[3738]),
			.E(gen[3740]),

			.SO(gen[3833]),
			.S(gen[3834]),
			.SE(gen[3835]),

			.SELF(gen[3739]),
			.cell_state(gen[3739])
		); 

/******************* CELL 3740 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3740 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3644]),
			.N(gen[3645]),
			.NE(gen[3646]),

			.O(gen[3739]),
			.E(gen[3741]),

			.SO(gen[3834]),
			.S(gen[3835]),
			.SE(gen[3836]),

			.SELF(gen[3740]),
			.cell_state(gen[3740])
		); 

/******************* CELL 3741 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3741 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3645]),
			.N(gen[3646]),
			.NE(gen[3647]),

			.O(gen[3740]),
			.E(gen[3742]),

			.SO(gen[3835]),
			.S(gen[3836]),
			.SE(gen[3837]),

			.SELF(gen[3741]),
			.cell_state(gen[3741])
		); 

/******************* CELL 3742 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3742 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3646]),
			.N(gen[3647]),
			.NE(gen[3648]),

			.O(gen[3741]),
			.E(gen[3743]),

			.SO(gen[3836]),
			.S(gen[3837]),
			.SE(gen[3838]),

			.SELF(gen[3742]),
			.cell_state(gen[3742])
		); 

/******************* CELL 3743 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3743 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3647]),
			.N(gen[3648]),
			.NE(gen[3649]),

			.O(gen[3742]),
			.E(gen[3744]),

			.SO(gen[3837]),
			.S(gen[3838]),
			.SE(gen[3839]),

			.SELF(gen[3743]),
			.cell_state(gen[3743])
		); 

/******************* CELL 3744 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3744 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3648]),
			.N(gen[3649]),
			.NE(gen[3650]),

			.O(gen[3743]),
			.E(gen[3745]),

			.SO(gen[3838]),
			.S(gen[3839]),
			.SE(gen[3840]),

			.SELF(gen[3744]),
			.cell_state(gen[3744])
		); 

/******************* CELL 3745 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3745 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3649]),
			.N(gen[3650]),
			.NE(gen[3651]),

			.O(gen[3744]),
			.E(gen[3746]),

			.SO(gen[3839]),
			.S(gen[3840]),
			.SE(gen[3841]),

			.SELF(gen[3745]),
			.cell_state(gen[3745])
		); 

/******************* CELL 3746 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3746 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3650]),
			.N(gen[3651]),
			.NE(gen[3652]),

			.O(gen[3745]),
			.E(gen[3747]),

			.SO(gen[3840]),
			.S(gen[3841]),
			.SE(gen[3842]),

			.SELF(gen[3746]),
			.cell_state(gen[3746])
		); 

/******************* CELL 3747 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3747 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3651]),
			.N(gen[3652]),
			.NE(gen[3653]),

			.O(gen[3746]),
			.E(gen[3748]),

			.SO(gen[3841]),
			.S(gen[3842]),
			.SE(gen[3843]),

			.SELF(gen[3747]),
			.cell_state(gen[3747])
		); 

/******************* CELL 3748 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3748 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3652]),
			.N(gen[3653]),
			.NE(gen[3654]),

			.O(gen[3747]),
			.E(gen[3749]),

			.SO(gen[3842]),
			.S(gen[3843]),
			.SE(gen[3844]),

			.SELF(gen[3748]),
			.cell_state(gen[3748])
		); 

/******************* CELL 3749 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3749 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3653]),
			.N(gen[3654]),
			.NE(gen[3655]),

			.O(gen[3748]),
			.E(gen[3750]),

			.SO(gen[3843]),
			.S(gen[3844]),
			.SE(gen[3845]),

			.SELF(gen[3749]),
			.cell_state(gen[3749])
		); 

/******************* CELL 3750 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3750 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3654]),
			.N(gen[3655]),
			.NE(gen[3656]),

			.O(gen[3749]),
			.E(gen[3751]),

			.SO(gen[3844]),
			.S(gen[3845]),
			.SE(gen[3846]),

			.SELF(gen[3750]),
			.cell_state(gen[3750])
		); 

/******************* CELL 3751 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3751 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3655]),
			.N(gen[3656]),
			.NE(gen[3657]),

			.O(gen[3750]),
			.E(gen[3752]),

			.SO(gen[3845]),
			.S(gen[3846]),
			.SE(gen[3847]),

			.SELF(gen[3751]),
			.cell_state(gen[3751])
		); 

/******************* CELL 3752 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3752 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3656]),
			.N(gen[3657]),
			.NE(gen[3658]),

			.O(gen[3751]),
			.E(gen[3753]),

			.SO(gen[3846]),
			.S(gen[3847]),
			.SE(gen[3848]),

			.SELF(gen[3752]),
			.cell_state(gen[3752])
		); 

/******************* CELL 3753 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3753 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3657]),
			.N(gen[3658]),
			.NE(gen[3659]),

			.O(gen[3752]),
			.E(gen[3754]),

			.SO(gen[3847]),
			.S(gen[3848]),
			.SE(gen[3849]),

			.SELF(gen[3753]),
			.cell_state(gen[3753])
		); 

/******************* CELL 3754 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3754 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3658]),
			.N(gen[3659]),
			.NE(gen[3660]),

			.O(gen[3753]),
			.E(gen[3755]),

			.SO(gen[3848]),
			.S(gen[3849]),
			.SE(gen[3850]),

			.SELF(gen[3754]),
			.cell_state(gen[3754])
		); 

/******************* CELL 3755 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3755 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3659]),
			.N(gen[3660]),
			.NE(gen[3661]),

			.O(gen[3754]),
			.E(gen[3756]),

			.SO(gen[3849]),
			.S(gen[3850]),
			.SE(gen[3851]),

			.SELF(gen[3755]),
			.cell_state(gen[3755])
		); 

/******************* CELL 3756 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3756 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3660]),
			.N(gen[3661]),
			.NE(gen[3662]),

			.O(gen[3755]),
			.E(gen[3757]),

			.SO(gen[3850]),
			.S(gen[3851]),
			.SE(gen[3852]),

			.SELF(gen[3756]),
			.cell_state(gen[3756])
		); 

/******************* CELL 3757 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3757 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3661]),
			.N(gen[3662]),
			.NE(gen[3663]),

			.O(gen[3756]),
			.E(gen[3758]),

			.SO(gen[3851]),
			.S(gen[3852]),
			.SE(gen[3853]),

			.SELF(gen[3757]),
			.cell_state(gen[3757])
		); 

/******************* CELL 3758 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3758 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3662]),
			.N(gen[3663]),
			.NE(gen[3664]),

			.O(gen[3757]),
			.E(gen[3759]),

			.SO(gen[3852]),
			.S(gen[3853]),
			.SE(gen[3854]),

			.SELF(gen[3758]),
			.cell_state(gen[3758])
		); 

/******************* CELL 3759 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3759 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3663]),
			.N(gen[3664]),
			.NE(gen[3665]),

			.O(gen[3758]),
			.E(gen[3760]),

			.SO(gen[3853]),
			.S(gen[3854]),
			.SE(gen[3855]),

			.SELF(gen[3759]),
			.cell_state(gen[3759])
		); 

/******************* CELL 3760 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3760 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3664]),
			.N(gen[3665]),
			.NE(gen[3666]),

			.O(gen[3759]),
			.E(gen[3761]),

			.SO(gen[3854]),
			.S(gen[3855]),
			.SE(gen[3856]),

			.SELF(gen[3760]),
			.cell_state(gen[3760])
		); 

/******************* CELL 3761 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3761 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3665]),
			.N(gen[3666]),
			.NE(gen[3667]),

			.O(gen[3760]),
			.E(gen[3762]),

			.SO(gen[3855]),
			.S(gen[3856]),
			.SE(gen[3857]),

			.SELF(gen[3761]),
			.cell_state(gen[3761])
		); 

/******************* CELL 3762 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3762 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3666]),
			.N(gen[3667]),
			.NE(gen[3668]),

			.O(gen[3761]),
			.E(gen[3763]),

			.SO(gen[3856]),
			.S(gen[3857]),
			.SE(gen[3858]),

			.SELF(gen[3762]),
			.cell_state(gen[3762])
		); 

/******************* CELL 3763 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3763 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3667]),
			.N(gen[3668]),
			.NE(gen[3669]),

			.O(gen[3762]),
			.E(gen[3764]),

			.SO(gen[3857]),
			.S(gen[3858]),
			.SE(gen[3859]),

			.SELF(gen[3763]),
			.cell_state(gen[3763])
		); 

/******************* CELL 3764 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3764 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3668]),
			.N(gen[3669]),
			.NE(gen[3670]),

			.O(gen[3763]),
			.E(gen[3765]),

			.SO(gen[3858]),
			.S(gen[3859]),
			.SE(gen[3860]),

			.SELF(gen[3764]),
			.cell_state(gen[3764])
		); 

/******************* CELL 3765 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3765 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3669]),
			.N(gen[3670]),
			.NE(gen[3671]),

			.O(gen[3764]),
			.E(gen[3766]),

			.SO(gen[3859]),
			.S(gen[3860]),
			.SE(gen[3861]),

			.SELF(gen[3765]),
			.cell_state(gen[3765])
		); 

/******************* CELL 3766 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3766 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3670]),
			.N(gen[3671]),
			.NE(gen[3672]),

			.O(gen[3765]),
			.E(gen[3767]),

			.SO(gen[3860]),
			.S(gen[3861]),
			.SE(gen[3862]),

			.SELF(gen[3766]),
			.cell_state(gen[3766])
		); 

/******************* CELL 3767 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3767 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3671]),
			.N(gen[3672]),
			.NE(gen[3673]),

			.O(gen[3766]),
			.E(gen[3768]),

			.SO(gen[3861]),
			.S(gen[3862]),
			.SE(gen[3863]),

			.SELF(gen[3767]),
			.cell_state(gen[3767])
		); 

/******************* CELL 3768 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3768 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3672]),
			.N(gen[3673]),
			.NE(gen[3674]),

			.O(gen[3767]),
			.E(gen[3769]),

			.SO(gen[3862]),
			.S(gen[3863]),
			.SE(gen[3864]),

			.SELF(gen[3768]),
			.cell_state(gen[3768])
		); 

/******************* CELL 3769 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3769 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3673]),
			.N(gen[3674]),
			.NE(gen[3675]),

			.O(gen[3768]),
			.E(gen[3770]),

			.SO(gen[3863]),
			.S(gen[3864]),
			.SE(gen[3865]),

			.SELF(gen[3769]),
			.cell_state(gen[3769])
		); 

/******************* CELL 3770 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3770 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3674]),
			.N(gen[3675]),
			.NE(gen[3676]),

			.O(gen[3769]),
			.E(gen[3771]),

			.SO(gen[3864]),
			.S(gen[3865]),
			.SE(gen[3866]),

			.SELF(gen[3770]),
			.cell_state(gen[3770])
		); 

/******************* CELL 3771 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3771 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3675]),
			.N(gen[3676]),
			.NE(gen[3677]),

			.O(gen[3770]),
			.E(gen[3772]),

			.SO(gen[3865]),
			.S(gen[3866]),
			.SE(gen[3867]),

			.SELF(gen[3771]),
			.cell_state(gen[3771])
		); 

/******************* CELL 3772 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3772 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3676]),
			.N(gen[3677]),
			.NE(gen[3678]),

			.O(gen[3771]),
			.E(gen[3773]),

			.SO(gen[3866]),
			.S(gen[3867]),
			.SE(gen[3868]),

			.SELF(gen[3772]),
			.cell_state(gen[3772])
		); 

/******************* CELL 3773 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3773 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3677]),
			.N(gen[3678]),
			.NE(gen[3679]),

			.O(gen[3772]),
			.E(gen[3774]),

			.SO(gen[3867]),
			.S(gen[3868]),
			.SE(gen[3869]),

			.SELF(gen[3773]),
			.cell_state(gen[3773])
		); 

/******************* CELL 3774 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3774 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3678]),
			.N(gen[3679]),
			.NE(gen[3680]),

			.O(gen[3773]),
			.E(gen[3775]),

			.SO(gen[3868]),
			.S(gen[3869]),
			.SE(gen[3870]),

			.SELF(gen[3774]),
			.cell_state(gen[3774])
		); 

/******************* CELL 3775 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3775 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3679]),
			.N(gen[3680]),
			.NE(gen[3681]),

			.O(gen[3774]),
			.E(gen[3776]),

			.SO(gen[3869]),
			.S(gen[3870]),
			.SE(gen[3871]),

			.SELF(gen[3775]),
			.cell_state(gen[3775])
		); 

/******************* CELL 3776 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3776 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3680]),
			.N(gen[3681]),
			.NE(gen[3682]),

			.O(gen[3775]),
			.E(gen[3777]),

			.SO(gen[3870]),
			.S(gen[3871]),
			.SE(gen[3872]),

			.SELF(gen[3776]),
			.cell_state(gen[3776])
		); 

/******************* CELL 3777 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3777 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3681]),
			.N(gen[3682]),
			.NE(gen[3683]),

			.O(gen[3776]),
			.E(gen[3778]),

			.SO(gen[3871]),
			.S(gen[3872]),
			.SE(gen[3873]),

			.SELF(gen[3777]),
			.cell_state(gen[3777])
		); 

/******************* CELL 3778 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3778 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3682]),
			.N(gen[3683]),
			.NE(gen[3684]),

			.O(gen[3777]),
			.E(gen[3779]),

			.SO(gen[3872]),
			.S(gen[3873]),
			.SE(gen[3874]),

			.SELF(gen[3778]),
			.cell_state(gen[3778])
		); 

/******************* CELL 3779 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3779 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3683]),
			.N(gen[3684]),
			.NE(gen[3685]),

			.O(gen[3778]),
			.E(gen[3780]),

			.SO(gen[3873]),
			.S(gen[3874]),
			.SE(gen[3875]),

			.SELF(gen[3779]),
			.cell_state(gen[3779])
		); 

/******************* CELL 3780 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3780 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3684]),
			.N(gen[3685]),
			.NE(gen[3686]),

			.O(gen[3779]),
			.E(gen[3781]),

			.SO(gen[3874]),
			.S(gen[3875]),
			.SE(gen[3876]),

			.SELF(gen[3780]),
			.cell_state(gen[3780])
		); 

/******************* CELL 3781 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3781 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3685]),
			.N(gen[3686]),
			.NE(gen[3687]),

			.O(gen[3780]),
			.E(gen[3782]),

			.SO(gen[3875]),
			.S(gen[3876]),
			.SE(gen[3877]),

			.SELF(gen[3781]),
			.cell_state(gen[3781])
		); 

/******************* CELL 3782 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3782 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3686]),
			.N(gen[3687]),
			.NE(gen[3688]),

			.O(gen[3781]),
			.E(gen[3783]),

			.SO(gen[3876]),
			.S(gen[3877]),
			.SE(gen[3878]),

			.SELF(gen[3782]),
			.cell_state(gen[3782])
		); 

/******************* CELL 3783 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3783 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3687]),
			.N(gen[3688]),
			.NE(gen[3689]),

			.O(gen[3782]),
			.E(gen[3784]),

			.SO(gen[3877]),
			.S(gen[3878]),
			.SE(gen[3879]),

			.SELF(gen[3783]),
			.cell_state(gen[3783])
		); 

/******************* CELL 3784 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3784 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3688]),
			.N(gen[3689]),
			.NE(gen[3690]),

			.O(gen[3783]),
			.E(gen[3785]),

			.SO(gen[3878]),
			.S(gen[3879]),
			.SE(gen[3880]),

			.SELF(gen[3784]),
			.cell_state(gen[3784])
		); 

/******************* CELL 3785 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3785 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3689]),
			.N(gen[3690]),
			.NE(gen[3691]),

			.O(gen[3784]),
			.E(gen[3786]),

			.SO(gen[3879]),
			.S(gen[3880]),
			.SE(gen[3881]),

			.SELF(gen[3785]),
			.cell_state(gen[3785])
		); 

/******************* CELL 3786 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3786 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3690]),
			.N(gen[3691]),
			.NE(gen[3692]),

			.O(gen[3785]),
			.E(gen[3787]),

			.SO(gen[3880]),
			.S(gen[3881]),
			.SE(gen[3882]),

			.SELF(gen[3786]),
			.cell_state(gen[3786])
		); 

/******************* CELL 3787 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3787 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3691]),
			.N(gen[3692]),
			.NE(gen[3693]),

			.O(gen[3786]),
			.E(gen[3788]),

			.SO(gen[3881]),
			.S(gen[3882]),
			.SE(gen[3883]),

			.SELF(gen[3787]),
			.cell_state(gen[3787])
		); 

/******************* CELL 3788 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3788 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3692]),
			.N(gen[3693]),
			.NE(gen[3694]),

			.O(gen[3787]),
			.E(gen[3789]),

			.SO(gen[3882]),
			.S(gen[3883]),
			.SE(gen[3884]),

			.SELF(gen[3788]),
			.cell_state(gen[3788])
		); 

/******************* CELL 3789 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3789 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3693]),
			.N(gen[3694]),
			.NE(gen[3695]),

			.O(gen[3788]),
			.E(gen[3790]),

			.SO(gen[3883]),
			.S(gen[3884]),
			.SE(gen[3885]),

			.SELF(gen[3789]),
			.cell_state(gen[3789])
		); 

/******************* CELL 3790 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3790 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3694]),
			.N(gen[3695]),
			.NE(gen[3696]),

			.O(gen[3789]),
			.E(gen[3791]),

			.SO(gen[3884]),
			.S(gen[3885]),
			.SE(gen[3886]),

			.SELF(gen[3790]),
			.cell_state(gen[3790])
		); 

/******************* CELL 3791 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3791 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3695]),
			.N(gen[3696]),
			.NE(gen[3697]),

			.O(gen[3790]),
			.E(gen[3792]),

			.SO(gen[3885]),
			.S(gen[3886]),
			.SE(gen[3887]),

			.SELF(gen[3791]),
			.cell_state(gen[3791])
		); 

/******************* CELL 3792 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3792 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3696]),
			.N(gen[3697]),
			.NE(gen[3698]),

			.O(gen[3791]),
			.E(gen[3793]),

			.SO(gen[3886]),
			.S(gen[3887]),
			.SE(gen[3888]),

			.SELF(gen[3792]),
			.cell_state(gen[3792])
		); 

/******************* CELL 3793 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3793 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3697]),
			.N(gen[3698]),
			.NE(gen[3699]),

			.O(gen[3792]),
			.E(gen[3794]),

			.SO(gen[3887]),
			.S(gen[3888]),
			.SE(gen[3889]),

			.SELF(gen[3793]),
			.cell_state(gen[3793])
		); 

/******************* CELL 3794 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3794 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3698]),
			.N(gen[3699]),
			.NE(gen[3700]),

			.O(gen[3793]),
			.E(gen[3795]),

			.SO(gen[3888]),
			.S(gen[3889]),
			.SE(gen[3890]),

			.SELF(gen[3794]),
			.cell_state(gen[3794])
		); 

/******************* CELL 3795 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3795 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3699]),
			.N(gen[3700]),
			.NE(gen[3701]),

			.O(gen[3794]),
			.E(gen[3796]),

			.SO(gen[3889]),
			.S(gen[3890]),
			.SE(gen[3891]),

			.SELF(gen[3795]),
			.cell_state(gen[3795])
		); 

/******************* CELL 3796 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3796 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3700]),
			.N(gen[3701]),
			.NE(gen[3702]),

			.O(gen[3795]),
			.E(gen[3797]),

			.SO(gen[3890]),
			.S(gen[3891]),
			.SE(gen[3892]),

			.SELF(gen[3796]),
			.cell_state(gen[3796])
		); 

/******************* CELL 3797 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3797 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3701]),
			.N(gen[3702]),
			.NE(gen[3703]),

			.O(gen[3796]),
			.E(gen[3798]),

			.SO(gen[3891]),
			.S(gen[3892]),
			.SE(gen[3893]),

			.SELF(gen[3797]),
			.cell_state(gen[3797])
		); 

/******************* CELL 3798 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3798 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3702]),
			.N(gen[3703]),
			.NE(gen[3704]),

			.O(gen[3797]),
			.E(gen[3799]),

			.SO(gen[3892]),
			.S(gen[3893]),
			.SE(gen[3894]),

			.SELF(gen[3798]),
			.cell_state(gen[3798])
		); 

/******************* CELL 3799 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3799 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3703]),
			.N(gen[3704]),
			.NE(gen[3703]),

			.O(gen[3798]),
			.E(gen[3798]),

			.SO(gen[3893]),
			.S(gen[3894]),
			.SE(gen[3893]),

			.SELF(gen[3799]),
			.cell_state(gen[3799])
		); 

/******************* CELL 3800 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3800 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3706]),
			.N(gen[3705]),
			.NE(gen[3706]),

			.O(gen[3801]),
			.E(gen[3801]),

			.SO(gen[3896]),
			.S(gen[3895]),
			.SE(gen[3896]),

			.SELF(gen[3800]),
			.cell_state(gen[3800])
		); 

/******************* CELL 3801 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3801 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3705]),
			.N(gen[3706]),
			.NE(gen[3707]),

			.O(gen[3800]),
			.E(gen[3802]),

			.SO(gen[3895]),
			.S(gen[3896]),
			.SE(gen[3897]),

			.SELF(gen[3801]),
			.cell_state(gen[3801])
		); 

/******************* CELL 3802 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3802 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3706]),
			.N(gen[3707]),
			.NE(gen[3708]),

			.O(gen[3801]),
			.E(gen[3803]),

			.SO(gen[3896]),
			.S(gen[3897]),
			.SE(gen[3898]),

			.SELF(gen[3802]),
			.cell_state(gen[3802])
		); 

/******************* CELL 3803 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3803 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3707]),
			.N(gen[3708]),
			.NE(gen[3709]),

			.O(gen[3802]),
			.E(gen[3804]),

			.SO(gen[3897]),
			.S(gen[3898]),
			.SE(gen[3899]),

			.SELF(gen[3803]),
			.cell_state(gen[3803])
		); 

/******************* CELL 3804 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3804 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3708]),
			.N(gen[3709]),
			.NE(gen[3710]),

			.O(gen[3803]),
			.E(gen[3805]),

			.SO(gen[3898]),
			.S(gen[3899]),
			.SE(gen[3900]),

			.SELF(gen[3804]),
			.cell_state(gen[3804])
		); 

/******************* CELL 3805 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3805 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3709]),
			.N(gen[3710]),
			.NE(gen[3711]),

			.O(gen[3804]),
			.E(gen[3806]),

			.SO(gen[3899]),
			.S(gen[3900]),
			.SE(gen[3901]),

			.SELF(gen[3805]),
			.cell_state(gen[3805])
		); 

/******************* CELL 3806 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3806 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3710]),
			.N(gen[3711]),
			.NE(gen[3712]),

			.O(gen[3805]),
			.E(gen[3807]),

			.SO(gen[3900]),
			.S(gen[3901]),
			.SE(gen[3902]),

			.SELF(gen[3806]),
			.cell_state(gen[3806])
		); 

/******************* CELL 3807 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3807 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3711]),
			.N(gen[3712]),
			.NE(gen[3713]),

			.O(gen[3806]),
			.E(gen[3808]),

			.SO(gen[3901]),
			.S(gen[3902]),
			.SE(gen[3903]),

			.SELF(gen[3807]),
			.cell_state(gen[3807])
		); 

/******************* CELL 3808 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3808 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3712]),
			.N(gen[3713]),
			.NE(gen[3714]),

			.O(gen[3807]),
			.E(gen[3809]),

			.SO(gen[3902]),
			.S(gen[3903]),
			.SE(gen[3904]),

			.SELF(gen[3808]),
			.cell_state(gen[3808])
		); 

/******************* CELL 3809 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3809 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3713]),
			.N(gen[3714]),
			.NE(gen[3715]),

			.O(gen[3808]),
			.E(gen[3810]),

			.SO(gen[3903]),
			.S(gen[3904]),
			.SE(gen[3905]),

			.SELF(gen[3809]),
			.cell_state(gen[3809])
		); 

/******************* CELL 3810 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3810 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3714]),
			.N(gen[3715]),
			.NE(gen[3716]),

			.O(gen[3809]),
			.E(gen[3811]),

			.SO(gen[3904]),
			.S(gen[3905]),
			.SE(gen[3906]),

			.SELF(gen[3810]),
			.cell_state(gen[3810])
		); 

/******************* CELL 3811 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3811 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3715]),
			.N(gen[3716]),
			.NE(gen[3717]),

			.O(gen[3810]),
			.E(gen[3812]),

			.SO(gen[3905]),
			.S(gen[3906]),
			.SE(gen[3907]),

			.SELF(gen[3811]),
			.cell_state(gen[3811])
		); 

/******************* CELL 3812 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3812 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3716]),
			.N(gen[3717]),
			.NE(gen[3718]),

			.O(gen[3811]),
			.E(gen[3813]),

			.SO(gen[3906]),
			.S(gen[3907]),
			.SE(gen[3908]),

			.SELF(gen[3812]),
			.cell_state(gen[3812])
		); 

/******************* CELL 3813 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3813 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3717]),
			.N(gen[3718]),
			.NE(gen[3719]),

			.O(gen[3812]),
			.E(gen[3814]),

			.SO(gen[3907]),
			.S(gen[3908]),
			.SE(gen[3909]),

			.SELF(gen[3813]),
			.cell_state(gen[3813])
		); 

/******************* CELL 3814 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3814 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3718]),
			.N(gen[3719]),
			.NE(gen[3720]),

			.O(gen[3813]),
			.E(gen[3815]),

			.SO(gen[3908]),
			.S(gen[3909]),
			.SE(gen[3910]),

			.SELF(gen[3814]),
			.cell_state(gen[3814])
		); 

/******************* CELL 3815 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3815 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3719]),
			.N(gen[3720]),
			.NE(gen[3721]),

			.O(gen[3814]),
			.E(gen[3816]),

			.SO(gen[3909]),
			.S(gen[3910]),
			.SE(gen[3911]),

			.SELF(gen[3815]),
			.cell_state(gen[3815])
		); 

/******************* CELL 3816 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3816 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3720]),
			.N(gen[3721]),
			.NE(gen[3722]),

			.O(gen[3815]),
			.E(gen[3817]),

			.SO(gen[3910]),
			.S(gen[3911]),
			.SE(gen[3912]),

			.SELF(gen[3816]),
			.cell_state(gen[3816])
		); 

/******************* CELL 3817 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3817 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3721]),
			.N(gen[3722]),
			.NE(gen[3723]),

			.O(gen[3816]),
			.E(gen[3818]),

			.SO(gen[3911]),
			.S(gen[3912]),
			.SE(gen[3913]),

			.SELF(gen[3817]),
			.cell_state(gen[3817])
		); 

/******************* CELL 3818 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3818 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3722]),
			.N(gen[3723]),
			.NE(gen[3724]),

			.O(gen[3817]),
			.E(gen[3819]),

			.SO(gen[3912]),
			.S(gen[3913]),
			.SE(gen[3914]),

			.SELF(gen[3818]),
			.cell_state(gen[3818])
		); 

/******************* CELL 3819 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3819 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3723]),
			.N(gen[3724]),
			.NE(gen[3725]),

			.O(gen[3818]),
			.E(gen[3820]),

			.SO(gen[3913]),
			.S(gen[3914]),
			.SE(gen[3915]),

			.SELF(gen[3819]),
			.cell_state(gen[3819])
		); 

/******************* CELL 3820 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3820 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3724]),
			.N(gen[3725]),
			.NE(gen[3726]),

			.O(gen[3819]),
			.E(gen[3821]),

			.SO(gen[3914]),
			.S(gen[3915]),
			.SE(gen[3916]),

			.SELF(gen[3820]),
			.cell_state(gen[3820])
		); 

/******************* CELL 3821 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3821 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3725]),
			.N(gen[3726]),
			.NE(gen[3727]),

			.O(gen[3820]),
			.E(gen[3822]),

			.SO(gen[3915]),
			.S(gen[3916]),
			.SE(gen[3917]),

			.SELF(gen[3821]),
			.cell_state(gen[3821])
		); 

/******************* CELL 3822 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3822 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3726]),
			.N(gen[3727]),
			.NE(gen[3728]),

			.O(gen[3821]),
			.E(gen[3823]),

			.SO(gen[3916]),
			.S(gen[3917]),
			.SE(gen[3918]),

			.SELF(gen[3822]),
			.cell_state(gen[3822])
		); 

/******************* CELL 3823 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3823 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3727]),
			.N(gen[3728]),
			.NE(gen[3729]),

			.O(gen[3822]),
			.E(gen[3824]),

			.SO(gen[3917]),
			.S(gen[3918]),
			.SE(gen[3919]),

			.SELF(gen[3823]),
			.cell_state(gen[3823])
		); 

/******************* CELL 3824 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3824 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3728]),
			.N(gen[3729]),
			.NE(gen[3730]),

			.O(gen[3823]),
			.E(gen[3825]),

			.SO(gen[3918]),
			.S(gen[3919]),
			.SE(gen[3920]),

			.SELF(gen[3824]),
			.cell_state(gen[3824])
		); 

/******************* CELL 3825 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3825 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3729]),
			.N(gen[3730]),
			.NE(gen[3731]),

			.O(gen[3824]),
			.E(gen[3826]),

			.SO(gen[3919]),
			.S(gen[3920]),
			.SE(gen[3921]),

			.SELF(gen[3825]),
			.cell_state(gen[3825])
		); 

/******************* CELL 3826 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3826 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3730]),
			.N(gen[3731]),
			.NE(gen[3732]),

			.O(gen[3825]),
			.E(gen[3827]),

			.SO(gen[3920]),
			.S(gen[3921]),
			.SE(gen[3922]),

			.SELF(gen[3826]),
			.cell_state(gen[3826])
		); 

/******************* CELL 3827 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3827 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3731]),
			.N(gen[3732]),
			.NE(gen[3733]),

			.O(gen[3826]),
			.E(gen[3828]),

			.SO(gen[3921]),
			.S(gen[3922]),
			.SE(gen[3923]),

			.SELF(gen[3827]),
			.cell_state(gen[3827])
		); 

/******************* CELL 3828 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3828 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3732]),
			.N(gen[3733]),
			.NE(gen[3734]),

			.O(gen[3827]),
			.E(gen[3829]),

			.SO(gen[3922]),
			.S(gen[3923]),
			.SE(gen[3924]),

			.SELF(gen[3828]),
			.cell_state(gen[3828])
		); 

/******************* CELL 3829 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3829 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3733]),
			.N(gen[3734]),
			.NE(gen[3735]),

			.O(gen[3828]),
			.E(gen[3830]),

			.SO(gen[3923]),
			.S(gen[3924]),
			.SE(gen[3925]),

			.SELF(gen[3829]),
			.cell_state(gen[3829])
		); 

/******************* CELL 3830 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3830 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3734]),
			.N(gen[3735]),
			.NE(gen[3736]),

			.O(gen[3829]),
			.E(gen[3831]),

			.SO(gen[3924]),
			.S(gen[3925]),
			.SE(gen[3926]),

			.SELF(gen[3830]),
			.cell_state(gen[3830])
		); 

/******************* CELL 3831 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3831 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3735]),
			.N(gen[3736]),
			.NE(gen[3737]),

			.O(gen[3830]),
			.E(gen[3832]),

			.SO(gen[3925]),
			.S(gen[3926]),
			.SE(gen[3927]),

			.SELF(gen[3831]),
			.cell_state(gen[3831])
		); 

/******************* CELL 3832 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3832 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3736]),
			.N(gen[3737]),
			.NE(gen[3738]),

			.O(gen[3831]),
			.E(gen[3833]),

			.SO(gen[3926]),
			.S(gen[3927]),
			.SE(gen[3928]),

			.SELF(gen[3832]),
			.cell_state(gen[3832])
		); 

/******************* CELL 3833 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3833 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3737]),
			.N(gen[3738]),
			.NE(gen[3739]),

			.O(gen[3832]),
			.E(gen[3834]),

			.SO(gen[3927]),
			.S(gen[3928]),
			.SE(gen[3929]),

			.SELF(gen[3833]),
			.cell_state(gen[3833])
		); 

/******************* CELL 3834 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3834 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3738]),
			.N(gen[3739]),
			.NE(gen[3740]),

			.O(gen[3833]),
			.E(gen[3835]),

			.SO(gen[3928]),
			.S(gen[3929]),
			.SE(gen[3930]),

			.SELF(gen[3834]),
			.cell_state(gen[3834])
		); 

/******************* CELL 3835 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3835 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3739]),
			.N(gen[3740]),
			.NE(gen[3741]),

			.O(gen[3834]),
			.E(gen[3836]),

			.SO(gen[3929]),
			.S(gen[3930]),
			.SE(gen[3931]),

			.SELF(gen[3835]),
			.cell_state(gen[3835])
		); 

/******************* CELL 3836 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3836 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3740]),
			.N(gen[3741]),
			.NE(gen[3742]),

			.O(gen[3835]),
			.E(gen[3837]),

			.SO(gen[3930]),
			.S(gen[3931]),
			.SE(gen[3932]),

			.SELF(gen[3836]),
			.cell_state(gen[3836])
		); 

/******************* CELL 3837 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3837 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3741]),
			.N(gen[3742]),
			.NE(gen[3743]),

			.O(gen[3836]),
			.E(gen[3838]),

			.SO(gen[3931]),
			.S(gen[3932]),
			.SE(gen[3933]),

			.SELF(gen[3837]),
			.cell_state(gen[3837])
		); 

/******************* CELL 3838 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3838 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3742]),
			.N(gen[3743]),
			.NE(gen[3744]),

			.O(gen[3837]),
			.E(gen[3839]),

			.SO(gen[3932]),
			.S(gen[3933]),
			.SE(gen[3934]),

			.SELF(gen[3838]),
			.cell_state(gen[3838])
		); 

/******************* CELL 3839 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3839 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3743]),
			.N(gen[3744]),
			.NE(gen[3745]),

			.O(gen[3838]),
			.E(gen[3840]),

			.SO(gen[3933]),
			.S(gen[3934]),
			.SE(gen[3935]),

			.SELF(gen[3839]),
			.cell_state(gen[3839])
		); 

/******************* CELL 3840 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3840 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3744]),
			.N(gen[3745]),
			.NE(gen[3746]),

			.O(gen[3839]),
			.E(gen[3841]),

			.SO(gen[3934]),
			.S(gen[3935]),
			.SE(gen[3936]),

			.SELF(gen[3840]),
			.cell_state(gen[3840])
		); 

/******************* CELL 3841 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3841 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3745]),
			.N(gen[3746]),
			.NE(gen[3747]),

			.O(gen[3840]),
			.E(gen[3842]),

			.SO(gen[3935]),
			.S(gen[3936]),
			.SE(gen[3937]),

			.SELF(gen[3841]),
			.cell_state(gen[3841])
		); 

/******************* CELL 3842 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3842 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3746]),
			.N(gen[3747]),
			.NE(gen[3748]),

			.O(gen[3841]),
			.E(gen[3843]),

			.SO(gen[3936]),
			.S(gen[3937]),
			.SE(gen[3938]),

			.SELF(gen[3842]),
			.cell_state(gen[3842])
		); 

/******************* CELL 3843 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3843 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3747]),
			.N(gen[3748]),
			.NE(gen[3749]),

			.O(gen[3842]),
			.E(gen[3844]),

			.SO(gen[3937]),
			.S(gen[3938]),
			.SE(gen[3939]),

			.SELF(gen[3843]),
			.cell_state(gen[3843])
		); 

/******************* CELL 3844 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3844 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3748]),
			.N(gen[3749]),
			.NE(gen[3750]),

			.O(gen[3843]),
			.E(gen[3845]),

			.SO(gen[3938]),
			.S(gen[3939]),
			.SE(gen[3940]),

			.SELF(gen[3844]),
			.cell_state(gen[3844])
		); 

/******************* CELL 3845 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3845 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3749]),
			.N(gen[3750]),
			.NE(gen[3751]),

			.O(gen[3844]),
			.E(gen[3846]),

			.SO(gen[3939]),
			.S(gen[3940]),
			.SE(gen[3941]),

			.SELF(gen[3845]),
			.cell_state(gen[3845])
		); 

/******************* CELL 3846 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3846 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3750]),
			.N(gen[3751]),
			.NE(gen[3752]),

			.O(gen[3845]),
			.E(gen[3847]),

			.SO(gen[3940]),
			.S(gen[3941]),
			.SE(gen[3942]),

			.SELF(gen[3846]),
			.cell_state(gen[3846])
		); 

/******************* CELL 3847 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3847 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3751]),
			.N(gen[3752]),
			.NE(gen[3753]),

			.O(gen[3846]),
			.E(gen[3848]),

			.SO(gen[3941]),
			.S(gen[3942]),
			.SE(gen[3943]),

			.SELF(gen[3847]),
			.cell_state(gen[3847])
		); 

/******************* CELL 3848 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3848 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3752]),
			.N(gen[3753]),
			.NE(gen[3754]),

			.O(gen[3847]),
			.E(gen[3849]),

			.SO(gen[3942]),
			.S(gen[3943]),
			.SE(gen[3944]),

			.SELF(gen[3848]),
			.cell_state(gen[3848])
		); 

/******************* CELL 3849 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3849 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3753]),
			.N(gen[3754]),
			.NE(gen[3755]),

			.O(gen[3848]),
			.E(gen[3850]),

			.SO(gen[3943]),
			.S(gen[3944]),
			.SE(gen[3945]),

			.SELF(gen[3849]),
			.cell_state(gen[3849])
		); 

/******************* CELL 3850 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3850 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3754]),
			.N(gen[3755]),
			.NE(gen[3756]),

			.O(gen[3849]),
			.E(gen[3851]),

			.SO(gen[3944]),
			.S(gen[3945]),
			.SE(gen[3946]),

			.SELF(gen[3850]),
			.cell_state(gen[3850])
		); 

/******************* CELL 3851 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3851 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3755]),
			.N(gen[3756]),
			.NE(gen[3757]),

			.O(gen[3850]),
			.E(gen[3852]),

			.SO(gen[3945]),
			.S(gen[3946]),
			.SE(gen[3947]),

			.SELF(gen[3851]),
			.cell_state(gen[3851])
		); 

/******************* CELL 3852 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3852 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3756]),
			.N(gen[3757]),
			.NE(gen[3758]),

			.O(gen[3851]),
			.E(gen[3853]),

			.SO(gen[3946]),
			.S(gen[3947]),
			.SE(gen[3948]),

			.SELF(gen[3852]),
			.cell_state(gen[3852])
		); 

/******************* CELL 3853 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3853 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3757]),
			.N(gen[3758]),
			.NE(gen[3759]),

			.O(gen[3852]),
			.E(gen[3854]),

			.SO(gen[3947]),
			.S(gen[3948]),
			.SE(gen[3949]),

			.SELF(gen[3853]),
			.cell_state(gen[3853])
		); 

/******************* CELL 3854 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3854 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3758]),
			.N(gen[3759]),
			.NE(gen[3760]),

			.O(gen[3853]),
			.E(gen[3855]),

			.SO(gen[3948]),
			.S(gen[3949]),
			.SE(gen[3950]),

			.SELF(gen[3854]),
			.cell_state(gen[3854])
		); 

/******************* CELL 3855 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3855 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3759]),
			.N(gen[3760]),
			.NE(gen[3761]),

			.O(gen[3854]),
			.E(gen[3856]),

			.SO(gen[3949]),
			.S(gen[3950]),
			.SE(gen[3951]),

			.SELF(gen[3855]),
			.cell_state(gen[3855])
		); 

/******************* CELL 3856 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3856 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3760]),
			.N(gen[3761]),
			.NE(gen[3762]),

			.O(gen[3855]),
			.E(gen[3857]),

			.SO(gen[3950]),
			.S(gen[3951]),
			.SE(gen[3952]),

			.SELF(gen[3856]),
			.cell_state(gen[3856])
		); 

/******************* CELL 3857 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3857 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3761]),
			.N(gen[3762]),
			.NE(gen[3763]),

			.O(gen[3856]),
			.E(gen[3858]),

			.SO(gen[3951]),
			.S(gen[3952]),
			.SE(gen[3953]),

			.SELF(gen[3857]),
			.cell_state(gen[3857])
		); 

/******************* CELL 3858 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3858 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3762]),
			.N(gen[3763]),
			.NE(gen[3764]),

			.O(gen[3857]),
			.E(gen[3859]),

			.SO(gen[3952]),
			.S(gen[3953]),
			.SE(gen[3954]),

			.SELF(gen[3858]),
			.cell_state(gen[3858])
		); 

/******************* CELL 3859 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3859 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3763]),
			.N(gen[3764]),
			.NE(gen[3765]),

			.O(gen[3858]),
			.E(gen[3860]),

			.SO(gen[3953]),
			.S(gen[3954]),
			.SE(gen[3955]),

			.SELF(gen[3859]),
			.cell_state(gen[3859])
		); 

/******************* CELL 3860 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3860 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3764]),
			.N(gen[3765]),
			.NE(gen[3766]),

			.O(gen[3859]),
			.E(gen[3861]),

			.SO(gen[3954]),
			.S(gen[3955]),
			.SE(gen[3956]),

			.SELF(gen[3860]),
			.cell_state(gen[3860])
		); 

/******************* CELL 3861 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3861 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3765]),
			.N(gen[3766]),
			.NE(gen[3767]),

			.O(gen[3860]),
			.E(gen[3862]),

			.SO(gen[3955]),
			.S(gen[3956]),
			.SE(gen[3957]),

			.SELF(gen[3861]),
			.cell_state(gen[3861])
		); 

/******************* CELL 3862 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3862 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3766]),
			.N(gen[3767]),
			.NE(gen[3768]),

			.O(gen[3861]),
			.E(gen[3863]),

			.SO(gen[3956]),
			.S(gen[3957]),
			.SE(gen[3958]),

			.SELF(gen[3862]),
			.cell_state(gen[3862])
		); 

/******************* CELL 3863 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3863 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3767]),
			.N(gen[3768]),
			.NE(gen[3769]),

			.O(gen[3862]),
			.E(gen[3864]),

			.SO(gen[3957]),
			.S(gen[3958]),
			.SE(gen[3959]),

			.SELF(gen[3863]),
			.cell_state(gen[3863])
		); 

/******************* CELL 3864 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3864 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3768]),
			.N(gen[3769]),
			.NE(gen[3770]),

			.O(gen[3863]),
			.E(gen[3865]),

			.SO(gen[3958]),
			.S(gen[3959]),
			.SE(gen[3960]),

			.SELF(gen[3864]),
			.cell_state(gen[3864])
		); 

/******************* CELL 3865 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3865 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3769]),
			.N(gen[3770]),
			.NE(gen[3771]),

			.O(gen[3864]),
			.E(gen[3866]),

			.SO(gen[3959]),
			.S(gen[3960]),
			.SE(gen[3961]),

			.SELF(gen[3865]),
			.cell_state(gen[3865])
		); 

/******************* CELL 3866 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3866 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3770]),
			.N(gen[3771]),
			.NE(gen[3772]),

			.O(gen[3865]),
			.E(gen[3867]),

			.SO(gen[3960]),
			.S(gen[3961]),
			.SE(gen[3962]),

			.SELF(gen[3866]),
			.cell_state(gen[3866])
		); 

/******************* CELL 3867 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3867 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3771]),
			.N(gen[3772]),
			.NE(gen[3773]),

			.O(gen[3866]),
			.E(gen[3868]),

			.SO(gen[3961]),
			.S(gen[3962]),
			.SE(gen[3963]),

			.SELF(gen[3867]),
			.cell_state(gen[3867])
		); 

/******************* CELL 3868 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3868 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3772]),
			.N(gen[3773]),
			.NE(gen[3774]),

			.O(gen[3867]),
			.E(gen[3869]),

			.SO(gen[3962]),
			.S(gen[3963]),
			.SE(gen[3964]),

			.SELF(gen[3868]),
			.cell_state(gen[3868])
		); 

/******************* CELL 3869 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3869 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3773]),
			.N(gen[3774]),
			.NE(gen[3775]),

			.O(gen[3868]),
			.E(gen[3870]),

			.SO(gen[3963]),
			.S(gen[3964]),
			.SE(gen[3965]),

			.SELF(gen[3869]),
			.cell_state(gen[3869])
		); 

/******************* CELL 3870 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3870 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3774]),
			.N(gen[3775]),
			.NE(gen[3776]),

			.O(gen[3869]),
			.E(gen[3871]),

			.SO(gen[3964]),
			.S(gen[3965]),
			.SE(gen[3966]),

			.SELF(gen[3870]),
			.cell_state(gen[3870])
		); 

/******************* CELL 3871 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3871 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3775]),
			.N(gen[3776]),
			.NE(gen[3777]),

			.O(gen[3870]),
			.E(gen[3872]),

			.SO(gen[3965]),
			.S(gen[3966]),
			.SE(gen[3967]),

			.SELF(gen[3871]),
			.cell_state(gen[3871])
		); 

/******************* CELL 3872 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3872 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3776]),
			.N(gen[3777]),
			.NE(gen[3778]),

			.O(gen[3871]),
			.E(gen[3873]),

			.SO(gen[3966]),
			.S(gen[3967]),
			.SE(gen[3968]),

			.SELF(gen[3872]),
			.cell_state(gen[3872])
		); 

/******************* CELL 3873 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3873 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3777]),
			.N(gen[3778]),
			.NE(gen[3779]),

			.O(gen[3872]),
			.E(gen[3874]),

			.SO(gen[3967]),
			.S(gen[3968]),
			.SE(gen[3969]),

			.SELF(gen[3873]),
			.cell_state(gen[3873])
		); 

/******************* CELL 3874 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3874 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3778]),
			.N(gen[3779]),
			.NE(gen[3780]),

			.O(gen[3873]),
			.E(gen[3875]),

			.SO(gen[3968]),
			.S(gen[3969]),
			.SE(gen[3970]),

			.SELF(gen[3874]),
			.cell_state(gen[3874])
		); 

/******************* CELL 3875 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3875 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3779]),
			.N(gen[3780]),
			.NE(gen[3781]),

			.O(gen[3874]),
			.E(gen[3876]),

			.SO(gen[3969]),
			.S(gen[3970]),
			.SE(gen[3971]),

			.SELF(gen[3875]),
			.cell_state(gen[3875])
		); 

/******************* CELL 3876 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3876 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3780]),
			.N(gen[3781]),
			.NE(gen[3782]),

			.O(gen[3875]),
			.E(gen[3877]),

			.SO(gen[3970]),
			.S(gen[3971]),
			.SE(gen[3972]),

			.SELF(gen[3876]),
			.cell_state(gen[3876])
		); 

/******************* CELL 3877 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3877 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3781]),
			.N(gen[3782]),
			.NE(gen[3783]),

			.O(gen[3876]),
			.E(gen[3878]),

			.SO(gen[3971]),
			.S(gen[3972]),
			.SE(gen[3973]),

			.SELF(gen[3877]),
			.cell_state(gen[3877])
		); 

/******************* CELL 3878 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3878 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3782]),
			.N(gen[3783]),
			.NE(gen[3784]),

			.O(gen[3877]),
			.E(gen[3879]),

			.SO(gen[3972]),
			.S(gen[3973]),
			.SE(gen[3974]),

			.SELF(gen[3878]),
			.cell_state(gen[3878])
		); 

/******************* CELL 3879 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3879 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3783]),
			.N(gen[3784]),
			.NE(gen[3785]),

			.O(gen[3878]),
			.E(gen[3880]),

			.SO(gen[3973]),
			.S(gen[3974]),
			.SE(gen[3975]),

			.SELF(gen[3879]),
			.cell_state(gen[3879])
		); 

/******************* CELL 3880 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3880 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3784]),
			.N(gen[3785]),
			.NE(gen[3786]),

			.O(gen[3879]),
			.E(gen[3881]),

			.SO(gen[3974]),
			.S(gen[3975]),
			.SE(gen[3976]),

			.SELF(gen[3880]),
			.cell_state(gen[3880])
		); 

/******************* CELL 3881 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3881 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3785]),
			.N(gen[3786]),
			.NE(gen[3787]),

			.O(gen[3880]),
			.E(gen[3882]),

			.SO(gen[3975]),
			.S(gen[3976]),
			.SE(gen[3977]),

			.SELF(gen[3881]),
			.cell_state(gen[3881])
		); 

/******************* CELL 3882 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3882 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3786]),
			.N(gen[3787]),
			.NE(gen[3788]),

			.O(gen[3881]),
			.E(gen[3883]),

			.SO(gen[3976]),
			.S(gen[3977]),
			.SE(gen[3978]),

			.SELF(gen[3882]),
			.cell_state(gen[3882])
		); 

/******************* CELL 3883 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3883 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3787]),
			.N(gen[3788]),
			.NE(gen[3789]),

			.O(gen[3882]),
			.E(gen[3884]),

			.SO(gen[3977]),
			.S(gen[3978]),
			.SE(gen[3979]),

			.SELF(gen[3883]),
			.cell_state(gen[3883])
		); 

/******************* CELL 3884 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3884 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3788]),
			.N(gen[3789]),
			.NE(gen[3790]),

			.O(gen[3883]),
			.E(gen[3885]),

			.SO(gen[3978]),
			.S(gen[3979]),
			.SE(gen[3980]),

			.SELF(gen[3884]),
			.cell_state(gen[3884])
		); 

/******************* CELL 3885 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3885 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3789]),
			.N(gen[3790]),
			.NE(gen[3791]),

			.O(gen[3884]),
			.E(gen[3886]),

			.SO(gen[3979]),
			.S(gen[3980]),
			.SE(gen[3981]),

			.SELF(gen[3885]),
			.cell_state(gen[3885])
		); 

/******************* CELL 3886 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3886 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3790]),
			.N(gen[3791]),
			.NE(gen[3792]),

			.O(gen[3885]),
			.E(gen[3887]),

			.SO(gen[3980]),
			.S(gen[3981]),
			.SE(gen[3982]),

			.SELF(gen[3886]),
			.cell_state(gen[3886])
		); 

/******************* CELL 3887 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3887 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3791]),
			.N(gen[3792]),
			.NE(gen[3793]),

			.O(gen[3886]),
			.E(gen[3888]),

			.SO(gen[3981]),
			.S(gen[3982]),
			.SE(gen[3983]),

			.SELF(gen[3887]),
			.cell_state(gen[3887])
		); 

/******************* CELL 3888 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3888 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3792]),
			.N(gen[3793]),
			.NE(gen[3794]),

			.O(gen[3887]),
			.E(gen[3889]),

			.SO(gen[3982]),
			.S(gen[3983]),
			.SE(gen[3984]),

			.SELF(gen[3888]),
			.cell_state(gen[3888])
		); 

/******************* CELL 3889 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3889 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3793]),
			.N(gen[3794]),
			.NE(gen[3795]),

			.O(gen[3888]),
			.E(gen[3890]),

			.SO(gen[3983]),
			.S(gen[3984]),
			.SE(gen[3985]),

			.SELF(gen[3889]),
			.cell_state(gen[3889])
		); 

/******************* CELL 3890 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3890 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3794]),
			.N(gen[3795]),
			.NE(gen[3796]),

			.O(gen[3889]),
			.E(gen[3891]),

			.SO(gen[3984]),
			.S(gen[3985]),
			.SE(gen[3986]),

			.SELF(gen[3890]),
			.cell_state(gen[3890])
		); 

/******************* CELL 3891 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3891 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3795]),
			.N(gen[3796]),
			.NE(gen[3797]),

			.O(gen[3890]),
			.E(gen[3892]),

			.SO(gen[3985]),
			.S(gen[3986]),
			.SE(gen[3987]),

			.SELF(gen[3891]),
			.cell_state(gen[3891])
		); 

/******************* CELL 3892 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3892 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3796]),
			.N(gen[3797]),
			.NE(gen[3798]),

			.O(gen[3891]),
			.E(gen[3893]),

			.SO(gen[3986]),
			.S(gen[3987]),
			.SE(gen[3988]),

			.SELF(gen[3892]),
			.cell_state(gen[3892])
		); 

/******************* CELL 3893 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3893 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3797]),
			.N(gen[3798]),
			.NE(gen[3799]),

			.O(gen[3892]),
			.E(gen[3894]),

			.SO(gen[3987]),
			.S(gen[3988]),
			.SE(gen[3989]),

			.SELF(gen[3893]),
			.cell_state(gen[3893])
		); 

/******************* CELL 3894 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3894 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3798]),
			.N(gen[3799]),
			.NE(gen[3798]),

			.O(gen[3893]),
			.E(gen[3893]),

			.SO(gen[3988]),
			.S(gen[3989]),
			.SE(gen[3988]),

			.SELF(gen[3894]),
			.cell_state(gen[3894])
		); 

/******************* CELL 3895 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3895 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3801]),
			.N(gen[3800]),
			.NE(gen[3801]),

			.O(gen[3896]),
			.E(gen[3896]),

			.SO(gen[3991]),
			.S(gen[3990]),
			.SE(gen[3991]),

			.SELF(gen[3895]),
			.cell_state(gen[3895])
		); 

/******************* CELL 3896 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3896 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3800]),
			.N(gen[3801]),
			.NE(gen[3802]),

			.O(gen[3895]),
			.E(gen[3897]),

			.SO(gen[3990]),
			.S(gen[3991]),
			.SE(gen[3992]),

			.SELF(gen[3896]),
			.cell_state(gen[3896])
		); 

/******************* CELL 3897 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3897 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3801]),
			.N(gen[3802]),
			.NE(gen[3803]),

			.O(gen[3896]),
			.E(gen[3898]),

			.SO(gen[3991]),
			.S(gen[3992]),
			.SE(gen[3993]),

			.SELF(gen[3897]),
			.cell_state(gen[3897])
		); 

/******************* CELL 3898 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3898 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3802]),
			.N(gen[3803]),
			.NE(gen[3804]),

			.O(gen[3897]),
			.E(gen[3899]),

			.SO(gen[3992]),
			.S(gen[3993]),
			.SE(gen[3994]),

			.SELF(gen[3898]),
			.cell_state(gen[3898])
		); 

/******************* CELL 3899 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3899 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3803]),
			.N(gen[3804]),
			.NE(gen[3805]),

			.O(gen[3898]),
			.E(gen[3900]),

			.SO(gen[3993]),
			.S(gen[3994]),
			.SE(gen[3995]),

			.SELF(gen[3899]),
			.cell_state(gen[3899])
		); 

/******************* CELL 3900 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3900 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3804]),
			.N(gen[3805]),
			.NE(gen[3806]),

			.O(gen[3899]),
			.E(gen[3901]),

			.SO(gen[3994]),
			.S(gen[3995]),
			.SE(gen[3996]),

			.SELF(gen[3900]),
			.cell_state(gen[3900])
		); 

/******************* CELL 3901 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3901 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3805]),
			.N(gen[3806]),
			.NE(gen[3807]),

			.O(gen[3900]),
			.E(gen[3902]),

			.SO(gen[3995]),
			.S(gen[3996]),
			.SE(gen[3997]),

			.SELF(gen[3901]),
			.cell_state(gen[3901])
		); 

/******************* CELL 3902 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3902 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3806]),
			.N(gen[3807]),
			.NE(gen[3808]),

			.O(gen[3901]),
			.E(gen[3903]),

			.SO(gen[3996]),
			.S(gen[3997]),
			.SE(gen[3998]),

			.SELF(gen[3902]),
			.cell_state(gen[3902])
		); 

/******************* CELL 3903 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3903 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3807]),
			.N(gen[3808]),
			.NE(gen[3809]),

			.O(gen[3902]),
			.E(gen[3904]),

			.SO(gen[3997]),
			.S(gen[3998]),
			.SE(gen[3999]),

			.SELF(gen[3903]),
			.cell_state(gen[3903])
		); 

/******************* CELL 3904 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3904 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3808]),
			.N(gen[3809]),
			.NE(gen[3810]),

			.O(gen[3903]),
			.E(gen[3905]),

			.SO(gen[3998]),
			.S(gen[3999]),
			.SE(gen[4000]),

			.SELF(gen[3904]),
			.cell_state(gen[3904])
		); 

/******************* CELL 3905 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3905 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3809]),
			.N(gen[3810]),
			.NE(gen[3811]),

			.O(gen[3904]),
			.E(gen[3906]),

			.SO(gen[3999]),
			.S(gen[4000]),
			.SE(gen[4001]),

			.SELF(gen[3905]),
			.cell_state(gen[3905])
		); 

/******************* CELL 3906 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3906 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3810]),
			.N(gen[3811]),
			.NE(gen[3812]),

			.O(gen[3905]),
			.E(gen[3907]),

			.SO(gen[4000]),
			.S(gen[4001]),
			.SE(gen[4002]),

			.SELF(gen[3906]),
			.cell_state(gen[3906])
		); 

/******************* CELL 3907 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3907 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3811]),
			.N(gen[3812]),
			.NE(gen[3813]),

			.O(gen[3906]),
			.E(gen[3908]),

			.SO(gen[4001]),
			.S(gen[4002]),
			.SE(gen[4003]),

			.SELF(gen[3907]),
			.cell_state(gen[3907])
		); 

/******************* CELL 3908 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3908 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3812]),
			.N(gen[3813]),
			.NE(gen[3814]),

			.O(gen[3907]),
			.E(gen[3909]),

			.SO(gen[4002]),
			.S(gen[4003]),
			.SE(gen[4004]),

			.SELF(gen[3908]),
			.cell_state(gen[3908])
		); 

/******************* CELL 3909 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3909 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3813]),
			.N(gen[3814]),
			.NE(gen[3815]),

			.O(gen[3908]),
			.E(gen[3910]),

			.SO(gen[4003]),
			.S(gen[4004]),
			.SE(gen[4005]),

			.SELF(gen[3909]),
			.cell_state(gen[3909])
		); 

/******************* CELL 3910 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3910 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3814]),
			.N(gen[3815]),
			.NE(gen[3816]),

			.O(gen[3909]),
			.E(gen[3911]),

			.SO(gen[4004]),
			.S(gen[4005]),
			.SE(gen[4006]),

			.SELF(gen[3910]),
			.cell_state(gen[3910])
		); 

/******************* CELL 3911 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3911 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3815]),
			.N(gen[3816]),
			.NE(gen[3817]),

			.O(gen[3910]),
			.E(gen[3912]),

			.SO(gen[4005]),
			.S(gen[4006]),
			.SE(gen[4007]),

			.SELF(gen[3911]),
			.cell_state(gen[3911])
		); 

/******************* CELL 3912 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3912 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3816]),
			.N(gen[3817]),
			.NE(gen[3818]),

			.O(gen[3911]),
			.E(gen[3913]),

			.SO(gen[4006]),
			.S(gen[4007]),
			.SE(gen[4008]),

			.SELF(gen[3912]),
			.cell_state(gen[3912])
		); 

/******************* CELL 3913 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3913 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3817]),
			.N(gen[3818]),
			.NE(gen[3819]),

			.O(gen[3912]),
			.E(gen[3914]),

			.SO(gen[4007]),
			.S(gen[4008]),
			.SE(gen[4009]),

			.SELF(gen[3913]),
			.cell_state(gen[3913])
		); 

/******************* CELL 3914 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3914 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3818]),
			.N(gen[3819]),
			.NE(gen[3820]),

			.O(gen[3913]),
			.E(gen[3915]),

			.SO(gen[4008]),
			.S(gen[4009]),
			.SE(gen[4010]),

			.SELF(gen[3914]),
			.cell_state(gen[3914])
		); 

/******************* CELL 3915 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3915 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3819]),
			.N(gen[3820]),
			.NE(gen[3821]),

			.O(gen[3914]),
			.E(gen[3916]),

			.SO(gen[4009]),
			.S(gen[4010]),
			.SE(gen[4011]),

			.SELF(gen[3915]),
			.cell_state(gen[3915])
		); 

/******************* CELL 3916 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3916 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3820]),
			.N(gen[3821]),
			.NE(gen[3822]),

			.O(gen[3915]),
			.E(gen[3917]),

			.SO(gen[4010]),
			.S(gen[4011]),
			.SE(gen[4012]),

			.SELF(gen[3916]),
			.cell_state(gen[3916])
		); 

/******************* CELL 3917 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3917 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3821]),
			.N(gen[3822]),
			.NE(gen[3823]),

			.O(gen[3916]),
			.E(gen[3918]),

			.SO(gen[4011]),
			.S(gen[4012]),
			.SE(gen[4013]),

			.SELF(gen[3917]),
			.cell_state(gen[3917])
		); 

/******************* CELL 3918 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3918 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3822]),
			.N(gen[3823]),
			.NE(gen[3824]),

			.O(gen[3917]),
			.E(gen[3919]),

			.SO(gen[4012]),
			.S(gen[4013]),
			.SE(gen[4014]),

			.SELF(gen[3918]),
			.cell_state(gen[3918])
		); 

/******************* CELL 3919 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3919 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3823]),
			.N(gen[3824]),
			.NE(gen[3825]),

			.O(gen[3918]),
			.E(gen[3920]),

			.SO(gen[4013]),
			.S(gen[4014]),
			.SE(gen[4015]),

			.SELF(gen[3919]),
			.cell_state(gen[3919])
		); 

/******************* CELL 3920 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3920 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3824]),
			.N(gen[3825]),
			.NE(gen[3826]),

			.O(gen[3919]),
			.E(gen[3921]),

			.SO(gen[4014]),
			.S(gen[4015]),
			.SE(gen[4016]),

			.SELF(gen[3920]),
			.cell_state(gen[3920])
		); 

/******************* CELL 3921 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3921 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3825]),
			.N(gen[3826]),
			.NE(gen[3827]),

			.O(gen[3920]),
			.E(gen[3922]),

			.SO(gen[4015]),
			.S(gen[4016]),
			.SE(gen[4017]),

			.SELF(gen[3921]),
			.cell_state(gen[3921])
		); 

/******************* CELL 3922 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3922 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3826]),
			.N(gen[3827]),
			.NE(gen[3828]),

			.O(gen[3921]),
			.E(gen[3923]),

			.SO(gen[4016]),
			.S(gen[4017]),
			.SE(gen[4018]),

			.SELF(gen[3922]),
			.cell_state(gen[3922])
		); 

/******************* CELL 3923 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3923 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3827]),
			.N(gen[3828]),
			.NE(gen[3829]),

			.O(gen[3922]),
			.E(gen[3924]),

			.SO(gen[4017]),
			.S(gen[4018]),
			.SE(gen[4019]),

			.SELF(gen[3923]),
			.cell_state(gen[3923])
		); 

/******************* CELL 3924 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3924 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3828]),
			.N(gen[3829]),
			.NE(gen[3830]),

			.O(gen[3923]),
			.E(gen[3925]),

			.SO(gen[4018]),
			.S(gen[4019]),
			.SE(gen[4020]),

			.SELF(gen[3924]),
			.cell_state(gen[3924])
		); 

/******************* CELL 3925 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3925 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3829]),
			.N(gen[3830]),
			.NE(gen[3831]),

			.O(gen[3924]),
			.E(gen[3926]),

			.SO(gen[4019]),
			.S(gen[4020]),
			.SE(gen[4021]),

			.SELF(gen[3925]),
			.cell_state(gen[3925])
		); 

/******************* CELL 3926 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3926 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3830]),
			.N(gen[3831]),
			.NE(gen[3832]),

			.O(gen[3925]),
			.E(gen[3927]),

			.SO(gen[4020]),
			.S(gen[4021]),
			.SE(gen[4022]),

			.SELF(gen[3926]),
			.cell_state(gen[3926])
		); 

/******************* CELL 3927 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3927 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3831]),
			.N(gen[3832]),
			.NE(gen[3833]),

			.O(gen[3926]),
			.E(gen[3928]),

			.SO(gen[4021]),
			.S(gen[4022]),
			.SE(gen[4023]),

			.SELF(gen[3927]),
			.cell_state(gen[3927])
		); 

/******************* CELL 3928 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3928 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3832]),
			.N(gen[3833]),
			.NE(gen[3834]),

			.O(gen[3927]),
			.E(gen[3929]),

			.SO(gen[4022]),
			.S(gen[4023]),
			.SE(gen[4024]),

			.SELF(gen[3928]),
			.cell_state(gen[3928])
		); 

/******************* CELL 3929 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3929 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3833]),
			.N(gen[3834]),
			.NE(gen[3835]),

			.O(gen[3928]),
			.E(gen[3930]),

			.SO(gen[4023]),
			.S(gen[4024]),
			.SE(gen[4025]),

			.SELF(gen[3929]),
			.cell_state(gen[3929])
		); 

/******************* CELL 3930 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3930 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3834]),
			.N(gen[3835]),
			.NE(gen[3836]),

			.O(gen[3929]),
			.E(gen[3931]),

			.SO(gen[4024]),
			.S(gen[4025]),
			.SE(gen[4026]),

			.SELF(gen[3930]),
			.cell_state(gen[3930])
		); 

/******************* CELL 3931 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3931 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3835]),
			.N(gen[3836]),
			.NE(gen[3837]),

			.O(gen[3930]),
			.E(gen[3932]),

			.SO(gen[4025]),
			.S(gen[4026]),
			.SE(gen[4027]),

			.SELF(gen[3931]),
			.cell_state(gen[3931])
		); 

/******************* CELL 3932 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3932 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3836]),
			.N(gen[3837]),
			.NE(gen[3838]),

			.O(gen[3931]),
			.E(gen[3933]),

			.SO(gen[4026]),
			.S(gen[4027]),
			.SE(gen[4028]),

			.SELF(gen[3932]),
			.cell_state(gen[3932])
		); 

/******************* CELL 3933 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3933 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3837]),
			.N(gen[3838]),
			.NE(gen[3839]),

			.O(gen[3932]),
			.E(gen[3934]),

			.SO(gen[4027]),
			.S(gen[4028]),
			.SE(gen[4029]),

			.SELF(gen[3933]),
			.cell_state(gen[3933])
		); 

/******************* CELL 3934 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3934 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3838]),
			.N(gen[3839]),
			.NE(gen[3840]),

			.O(gen[3933]),
			.E(gen[3935]),

			.SO(gen[4028]),
			.S(gen[4029]),
			.SE(gen[4030]),

			.SELF(gen[3934]),
			.cell_state(gen[3934])
		); 

/******************* CELL 3935 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3935 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3839]),
			.N(gen[3840]),
			.NE(gen[3841]),

			.O(gen[3934]),
			.E(gen[3936]),

			.SO(gen[4029]),
			.S(gen[4030]),
			.SE(gen[4031]),

			.SELF(gen[3935]),
			.cell_state(gen[3935])
		); 

/******************* CELL 3936 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3936 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3840]),
			.N(gen[3841]),
			.NE(gen[3842]),

			.O(gen[3935]),
			.E(gen[3937]),

			.SO(gen[4030]),
			.S(gen[4031]),
			.SE(gen[4032]),

			.SELF(gen[3936]),
			.cell_state(gen[3936])
		); 

/******************* CELL 3937 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3937 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3841]),
			.N(gen[3842]),
			.NE(gen[3843]),

			.O(gen[3936]),
			.E(gen[3938]),

			.SO(gen[4031]),
			.S(gen[4032]),
			.SE(gen[4033]),

			.SELF(gen[3937]),
			.cell_state(gen[3937])
		); 

/******************* CELL 3938 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3938 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3842]),
			.N(gen[3843]),
			.NE(gen[3844]),

			.O(gen[3937]),
			.E(gen[3939]),

			.SO(gen[4032]),
			.S(gen[4033]),
			.SE(gen[4034]),

			.SELF(gen[3938]),
			.cell_state(gen[3938])
		); 

/******************* CELL 3939 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3939 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3843]),
			.N(gen[3844]),
			.NE(gen[3845]),

			.O(gen[3938]),
			.E(gen[3940]),

			.SO(gen[4033]),
			.S(gen[4034]),
			.SE(gen[4035]),

			.SELF(gen[3939]),
			.cell_state(gen[3939])
		); 

/******************* CELL 3940 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3940 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3844]),
			.N(gen[3845]),
			.NE(gen[3846]),

			.O(gen[3939]),
			.E(gen[3941]),

			.SO(gen[4034]),
			.S(gen[4035]),
			.SE(gen[4036]),

			.SELF(gen[3940]),
			.cell_state(gen[3940])
		); 

/******************* CELL 3941 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3941 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3845]),
			.N(gen[3846]),
			.NE(gen[3847]),

			.O(gen[3940]),
			.E(gen[3942]),

			.SO(gen[4035]),
			.S(gen[4036]),
			.SE(gen[4037]),

			.SELF(gen[3941]),
			.cell_state(gen[3941])
		); 

/******************* CELL 3942 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3942 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3846]),
			.N(gen[3847]),
			.NE(gen[3848]),

			.O(gen[3941]),
			.E(gen[3943]),

			.SO(gen[4036]),
			.S(gen[4037]),
			.SE(gen[4038]),

			.SELF(gen[3942]),
			.cell_state(gen[3942])
		); 

/******************* CELL 3943 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3943 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3847]),
			.N(gen[3848]),
			.NE(gen[3849]),

			.O(gen[3942]),
			.E(gen[3944]),

			.SO(gen[4037]),
			.S(gen[4038]),
			.SE(gen[4039]),

			.SELF(gen[3943]),
			.cell_state(gen[3943])
		); 

/******************* CELL 3944 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3944 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3848]),
			.N(gen[3849]),
			.NE(gen[3850]),

			.O(gen[3943]),
			.E(gen[3945]),

			.SO(gen[4038]),
			.S(gen[4039]),
			.SE(gen[4040]),

			.SELF(gen[3944]),
			.cell_state(gen[3944])
		); 

/******************* CELL 3945 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3945 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3849]),
			.N(gen[3850]),
			.NE(gen[3851]),

			.O(gen[3944]),
			.E(gen[3946]),

			.SO(gen[4039]),
			.S(gen[4040]),
			.SE(gen[4041]),

			.SELF(gen[3945]),
			.cell_state(gen[3945])
		); 

/******************* CELL 3946 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3946 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3850]),
			.N(gen[3851]),
			.NE(gen[3852]),

			.O(gen[3945]),
			.E(gen[3947]),

			.SO(gen[4040]),
			.S(gen[4041]),
			.SE(gen[4042]),

			.SELF(gen[3946]),
			.cell_state(gen[3946])
		); 

/******************* CELL 3947 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3947 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3851]),
			.N(gen[3852]),
			.NE(gen[3853]),

			.O(gen[3946]),
			.E(gen[3948]),

			.SO(gen[4041]),
			.S(gen[4042]),
			.SE(gen[4043]),

			.SELF(gen[3947]),
			.cell_state(gen[3947])
		); 

/******************* CELL 3948 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3948 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3852]),
			.N(gen[3853]),
			.NE(gen[3854]),

			.O(gen[3947]),
			.E(gen[3949]),

			.SO(gen[4042]),
			.S(gen[4043]),
			.SE(gen[4044]),

			.SELF(gen[3948]),
			.cell_state(gen[3948])
		); 

/******************* CELL 3949 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3949 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3853]),
			.N(gen[3854]),
			.NE(gen[3855]),

			.O(gen[3948]),
			.E(gen[3950]),

			.SO(gen[4043]),
			.S(gen[4044]),
			.SE(gen[4045]),

			.SELF(gen[3949]),
			.cell_state(gen[3949])
		); 

/******************* CELL 3950 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3950 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3854]),
			.N(gen[3855]),
			.NE(gen[3856]),

			.O(gen[3949]),
			.E(gen[3951]),

			.SO(gen[4044]),
			.S(gen[4045]),
			.SE(gen[4046]),

			.SELF(gen[3950]),
			.cell_state(gen[3950])
		); 

/******************* CELL 3951 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3951 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3855]),
			.N(gen[3856]),
			.NE(gen[3857]),

			.O(gen[3950]),
			.E(gen[3952]),

			.SO(gen[4045]),
			.S(gen[4046]),
			.SE(gen[4047]),

			.SELF(gen[3951]),
			.cell_state(gen[3951])
		); 

/******************* CELL 3952 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3952 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3856]),
			.N(gen[3857]),
			.NE(gen[3858]),

			.O(gen[3951]),
			.E(gen[3953]),

			.SO(gen[4046]),
			.S(gen[4047]),
			.SE(gen[4048]),

			.SELF(gen[3952]),
			.cell_state(gen[3952])
		); 

/******************* CELL 3953 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3953 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3857]),
			.N(gen[3858]),
			.NE(gen[3859]),

			.O(gen[3952]),
			.E(gen[3954]),

			.SO(gen[4047]),
			.S(gen[4048]),
			.SE(gen[4049]),

			.SELF(gen[3953]),
			.cell_state(gen[3953])
		); 

/******************* CELL 3954 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3954 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3858]),
			.N(gen[3859]),
			.NE(gen[3860]),

			.O(gen[3953]),
			.E(gen[3955]),

			.SO(gen[4048]),
			.S(gen[4049]),
			.SE(gen[4050]),

			.SELF(gen[3954]),
			.cell_state(gen[3954])
		); 

/******************* CELL 3955 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3955 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3859]),
			.N(gen[3860]),
			.NE(gen[3861]),

			.O(gen[3954]),
			.E(gen[3956]),

			.SO(gen[4049]),
			.S(gen[4050]),
			.SE(gen[4051]),

			.SELF(gen[3955]),
			.cell_state(gen[3955])
		); 

/******************* CELL 3956 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3956 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3860]),
			.N(gen[3861]),
			.NE(gen[3862]),

			.O(gen[3955]),
			.E(gen[3957]),

			.SO(gen[4050]),
			.S(gen[4051]),
			.SE(gen[4052]),

			.SELF(gen[3956]),
			.cell_state(gen[3956])
		); 

/******************* CELL 3957 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3957 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3861]),
			.N(gen[3862]),
			.NE(gen[3863]),

			.O(gen[3956]),
			.E(gen[3958]),

			.SO(gen[4051]),
			.S(gen[4052]),
			.SE(gen[4053]),

			.SELF(gen[3957]),
			.cell_state(gen[3957])
		); 

/******************* CELL 3958 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3958 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3862]),
			.N(gen[3863]),
			.NE(gen[3864]),

			.O(gen[3957]),
			.E(gen[3959]),

			.SO(gen[4052]),
			.S(gen[4053]),
			.SE(gen[4054]),

			.SELF(gen[3958]),
			.cell_state(gen[3958])
		); 

/******************* CELL 3959 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3959 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3863]),
			.N(gen[3864]),
			.NE(gen[3865]),

			.O(gen[3958]),
			.E(gen[3960]),

			.SO(gen[4053]),
			.S(gen[4054]),
			.SE(gen[4055]),

			.SELF(gen[3959]),
			.cell_state(gen[3959])
		); 

/******************* CELL 3960 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3960 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3864]),
			.N(gen[3865]),
			.NE(gen[3866]),

			.O(gen[3959]),
			.E(gen[3961]),

			.SO(gen[4054]),
			.S(gen[4055]),
			.SE(gen[4056]),

			.SELF(gen[3960]),
			.cell_state(gen[3960])
		); 

/******************* CELL 3961 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3961 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3865]),
			.N(gen[3866]),
			.NE(gen[3867]),

			.O(gen[3960]),
			.E(gen[3962]),

			.SO(gen[4055]),
			.S(gen[4056]),
			.SE(gen[4057]),

			.SELF(gen[3961]),
			.cell_state(gen[3961])
		); 

/******************* CELL 3962 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3962 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3866]),
			.N(gen[3867]),
			.NE(gen[3868]),

			.O(gen[3961]),
			.E(gen[3963]),

			.SO(gen[4056]),
			.S(gen[4057]),
			.SE(gen[4058]),

			.SELF(gen[3962]),
			.cell_state(gen[3962])
		); 

/******************* CELL 3963 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3963 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3867]),
			.N(gen[3868]),
			.NE(gen[3869]),

			.O(gen[3962]),
			.E(gen[3964]),

			.SO(gen[4057]),
			.S(gen[4058]),
			.SE(gen[4059]),

			.SELF(gen[3963]),
			.cell_state(gen[3963])
		); 

/******************* CELL 3964 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3964 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3868]),
			.N(gen[3869]),
			.NE(gen[3870]),

			.O(gen[3963]),
			.E(gen[3965]),

			.SO(gen[4058]),
			.S(gen[4059]),
			.SE(gen[4060]),

			.SELF(gen[3964]),
			.cell_state(gen[3964])
		); 

/******************* CELL 3965 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3965 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3869]),
			.N(gen[3870]),
			.NE(gen[3871]),

			.O(gen[3964]),
			.E(gen[3966]),

			.SO(gen[4059]),
			.S(gen[4060]),
			.SE(gen[4061]),

			.SELF(gen[3965]),
			.cell_state(gen[3965])
		); 

/******************* CELL 3966 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3966 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3870]),
			.N(gen[3871]),
			.NE(gen[3872]),

			.O(gen[3965]),
			.E(gen[3967]),

			.SO(gen[4060]),
			.S(gen[4061]),
			.SE(gen[4062]),

			.SELF(gen[3966]),
			.cell_state(gen[3966])
		); 

/******************* CELL 3967 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3967 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3871]),
			.N(gen[3872]),
			.NE(gen[3873]),

			.O(gen[3966]),
			.E(gen[3968]),

			.SO(gen[4061]),
			.S(gen[4062]),
			.SE(gen[4063]),

			.SELF(gen[3967]),
			.cell_state(gen[3967])
		); 

/******************* CELL 3968 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3968 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3872]),
			.N(gen[3873]),
			.NE(gen[3874]),

			.O(gen[3967]),
			.E(gen[3969]),

			.SO(gen[4062]),
			.S(gen[4063]),
			.SE(gen[4064]),

			.SELF(gen[3968]),
			.cell_state(gen[3968])
		); 

/******************* CELL 3969 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3969 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3873]),
			.N(gen[3874]),
			.NE(gen[3875]),

			.O(gen[3968]),
			.E(gen[3970]),

			.SO(gen[4063]),
			.S(gen[4064]),
			.SE(gen[4065]),

			.SELF(gen[3969]),
			.cell_state(gen[3969])
		); 

/******************* CELL 3970 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3970 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3874]),
			.N(gen[3875]),
			.NE(gen[3876]),

			.O(gen[3969]),
			.E(gen[3971]),

			.SO(gen[4064]),
			.S(gen[4065]),
			.SE(gen[4066]),

			.SELF(gen[3970]),
			.cell_state(gen[3970])
		); 

/******************* CELL 3971 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3971 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3875]),
			.N(gen[3876]),
			.NE(gen[3877]),

			.O(gen[3970]),
			.E(gen[3972]),

			.SO(gen[4065]),
			.S(gen[4066]),
			.SE(gen[4067]),

			.SELF(gen[3971]),
			.cell_state(gen[3971])
		); 

/******************* CELL 3972 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3972 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3876]),
			.N(gen[3877]),
			.NE(gen[3878]),

			.O(gen[3971]),
			.E(gen[3973]),

			.SO(gen[4066]),
			.S(gen[4067]),
			.SE(gen[4068]),

			.SELF(gen[3972]),
			.cell_state(gen[3972])
		); 

/******************* CELL 3973 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3973 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3877]),
			.N(gen[3878]),
			.NE(gen[3879]),

			.O(gen[3972]),
			.E(gen[3974]),

			.SO(gen[4067]),
			.S(gen[4068]),
			.SE(gen[4069]),

			.SELF(gen[3973]),
			.cell_state(gen[3973])
		); 

/******************* CELL 3974 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3974 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3878]),
			.N(gen[3879]),
			.NE(gen[3880]),

			.O(gen[3973]),
			.E(gen[3975]),

			.SO(gen[4068]),
			.S(gen[4069]),
			.SE(gen[4070]),

			.SELF(gen[3974]),
			.cell_state(gen[3974])
		); 

/******************* CELL 3975 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3975 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3879]),
			.N(gen[3880]),
			.NE(gen[3881]),

			.O(gen[3974]),
			.E(gen[3976]),

			.SO(gen[4069]),
			.S(gen[4070]),
			.SE(gen[4071]),

			.SELF(gen[3975]),
			.cell_state(gen[3975])
		); 

/******************* CELL 3976 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3976 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3880]),
			.N(gen[3881]),
			.NE(gen[3882]),

			.O(gen[3975]),
			.E(gen[3977]),

			.SO(gen[4070]),
			.S(gen[4071]),
			.SE(gen[4072]),

			.SELF(gen[3976]),
			.cell_state(gen[3976])
		); 

/******************* CELL 3977 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3977 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3881]),
			.N(gen[3882]),
			.NE(gen[3883]),

			.O(gen[3976]),
			.E(gen[3978]),

			.SO(gen[4071]),
			.S(gen[4072]),
			.SE(gen[4073]),

			.SELF(gen[3977]),
			.cell_state(gen[3977])
		); 

/******************* CELL 3978 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3978 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3882]),
			.N(gen[3883]),
			.NE(gen[3884]),

			.O(gen[3977]),
			.E(gen[3979]),

			.SO(gen[4072]),
			.S(gen[4073]),
			.SE(gen[4074]),

			.SELF(gen[3978]),
			.cell_state(gen[3978])
		); 

/******************* CELL 3979 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3979 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3883]),
			.N(gen[3884]),
			.NE(gen[3885]),

			.O(gen[3978]),
			.E(gen[3980]),

			.SO(gen[4073]),
			.S(gen[4074]),
			.SE(gen[4075]),

			.SELF(gen[3979]),
			.cell_state(gen[3979])
		); 

/******************* CELL 3980 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3980 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3884]),
			.N(gen[3885]),
			.NE(gen[3886]),

			.O(gen[3979]),
			.E(gen[3981]),

			.SO(gen[4074]),
			.S(gen[4075]),
			.SE(gen[4076]),

			.SELF(gen[3980]),
			.cell_state(gen[3980])
		); 

/******************* CELL 3981 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3981 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3885]),
			.N(gen[3886]),
			.NE(gen[3887]),

			.O(gen[3980]),
			.E(gen[3982]),

			.SO(gen[4075]),
			.S(gen[4076]),
			.SE(gen[4077]),

			.SELF(gen[3981]),
			.cell_state(gen[3981])
		); 

/******************* CELL 3982 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3982 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3886]),
			.N(gen[3887]),
			.NE(gen[3888]),

			.O(gen[3981]),
			.E(gen[3983]),

			.SO(gen[4076]),
			.S(gen[4077]),
			.SE(gen[4078]),

			.SELF(gen[3982]),
			.cell_state(gen[3982])
		); 

/******************* CELL 3983 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3983 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3887]),
			.N(gen[3888]),
			.NE(gen[3889]),

			.O(gen[3982]),
			.E(gen[3984]),

			.SO(gen[4077]),
			.S(gen[4078]),
			.SE(gen[4079]),

			.SELF(gen[3983]),
			.cell_state(gen[3983])
		); 

/******************* CELL 3984 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3984 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3888]),
			.N(gen[3889]),
			.NE(gen[3890]),

			.O(gen[3983]),
			.E(gen[3985]),

			.SO(gen[4078]),
			.S(gen[4079]),
			.SE(gen[4080]),

			.SELF(gen[3984]),
			.cell_state(gen[3984])
		); 

/******************* CELL 3985 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3985 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3889]),
			.N(gen[3890]),
			.NE(gen[3891]),

			.O(gen[3984]),
			.E(gen[3986]),

			.SO(gen[4079]),
			.S(gen[4080]),
			.SE(gen[4081]),

			.SELF(gen[3985]),
			.cell_state(gen[3985])
		); 

/******************* CELL 3986 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3986 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3890]),
			.N(gen[3891]),
			.NE(gen[3892]),

			.O(gen[3985]),
			.E(gen[3987]),

			.SO(gen[4080]),
			.S(gen[4081]),
			.SE(gen[4082]),

			.SELF(gen[3986]),
			.cell_state(gen[3986])
		); 

/******************* CELL 3987 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3987 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3891]),
			.N(gen[3892]),
			.NE(gen[3893]),

			.O(gen[3986]),
			.E(gen[3988]),

			.SO(gen[4081]),
			.S(gen[4082]),
			.SE(gen[4083]),

			.SELF(gen[3987]),
			.cell_state(gen[3987])
		); 

/******************* CELL 3988 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3988 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3892]),
			.N(gen[3893]),
			.NE(gen[3894]),

			.O(gen[3987]),
			.E(gen[3989]),

			.SO(gen[4082]),
			.S(gen[4083]),
			.SE(gen[4084]),

			.SELF(gen[3988]),
			.cell_state(gen[3988])
		); 

/******************* CELL 3989 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3989 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3893]),
			.N(gen[3894]),
			.NE(gen[3893]),

			.O(gen[3988]),
			.E(gen[3988]),

			.SO(gen[4083]),
			.S(gen[4084]),
			.SE(gen[4083]),

			.SELF(gen[3989]),
			.cell_state(gen[3989])
		); 

/******************* CELL 3990 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3990 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3896]),
			.N(gen[3895]),
			.NE(gen[3896]),

			.O(gen[3991]),
			.E(gen[3991]),

			.SO(gen[4086]),
			.S(gen[4085]),
			.SE(gen[4086]),

			.SELF(gen[3990]),
			.cell_state(gen[3990])
		); 

/******************* CELL 3991 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3991 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3895]),
			.N(gen[3896]),
			.NE(gen[3897]),

			.O(gen[3990]),
			.E(gen[3992]),

			.SO(gen[4085]),
			.S(gen[4086]),
			.SE(gen[4087]),

			.SELF(gen[3991]),
			.cell_state(gen[3991])
		); 

/******************* CELL 3992 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3992 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3896]),
			.N(gen[3897]),
			.NE(gen[3898]),

			.O(gen[3991]),
			.E(gen[3993]),

			.SO(gen[4086]),
			.S(gen[4087]),
			.SE(gen[4088]),

			.SELF(gen[3992]),
			.cell_state(gen[3992])
		); 

/******************* CELL 3993 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3993 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3897]),
			.N(gen[3898]),
			.NE(gen[3899]),

			.O(gen[3992]),
			.E(gen[3994]),

			.SO(gen[4087]),
			.S(gen[4088]),
			.SE(gen[4089]),

			.SELF(gen[3993]),
			.cell_state(gen[3993])
		); 

/******************* CELL 3994 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3994 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3898]),
			.N(gen[3899]),
			.NE(gen[3900]),

			.O(gen[3993]),
			.E(gen[3995]),

			.SO(gen[4088]),
			.S(gen[4089]),
			.SE(gen[4090]),

			.SELF(gen[3994]),
			.cell_state(gen[3994])
		); 

/******************* CELL 3995 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3995 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3899]),
			.N(gen[3900]),
			.NE(gen[3901]),

			.O(gen[3994]),
			.E(gen[3996]),

			.SO(gen[4089]),
			.S(gen[4090]),
			.SE(gen[4091]),

			.SELF(gen[3995]),
			.cell_state(gen[3995])
		); 

/******************* CELL 3996 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3996 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3900]),
			.N(gen[3901]),
			.NE(gen[3902]),

			.O(gen[3995]),
			.E(gen[3997]),

			.SO(gen[4090]),
			.S(gen[4091]),
			.SE(gen[4092]),

			.SELF(gen[3996]),
			.cell_state(gen[3996])
		); 

/******************* CELL 3997 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3997 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3901]),
			.N(gen[3902]),
			.NE(gen[3903]),

			.O(gen[3996]),
			.E(gen[3998]),

			.SO(gen[4091]),
			.S(gen[4092]),
			.SE(gen[4093]),

			.SELF(gen[3997]),
			.cell_state(gen[3997])
		); 

/******************* CELL 3998 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3998 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3902]),
			.N(gen[3903]),
			.NE(gen[3904]),

			.O(gen[3997]),
			.E(gen[3999]),

			.SO(gen[4092]),
			.S(gen[4093]),
			.SE(gen[4094]),

			.SELF(gen[3998]),
			.cell_state(gen[3998])
		); 

/******************* CELL 3999 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3999 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3903]),
			.N(gen[3904]),
			.NE(gen[3905]),

			.O(gen[3998]),
			.E(gen[4000]),

			.SO(gen[4093]),
			.S(gen[4094]),
			.SE(gen[4095]),

			.SELF(gen[3999]),
			.cell_state(gen[3999])
		); 

/******************* CELL 4000 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4000 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3904]),
			.N(gen[3905]),
			.NE(gen[3906]),

			.O(gen[3999]),
			.E(gen[4001]),

			.SO(gen[4094]),
			.S(gen[4095]),
			.SE(gen[4096]),

			.SELF(gen[4000]),
			.cell_state(gen[4000])
		); 

/******************* CELL 4001 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4001 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3905]),
			.N(gen[3906]),
			.NE(gen[3907]),

			.O(gen[4000]),
			.E(gen[4002]),

			.SO(gen[4095]),
			.S(gen[4096]),
			.SE(gen[4097]),

			.SELF(gen[4001]),
			.cell_state(gen[4001])
		); 

/******************* CELL 4002 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4002 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3906]),
			.N(gen[3907]),
			.NE(gen[3908]),

			.O(gen[4001]),
			.E(gen[4003]),

			.SO(gen[4096]),
			.S(gen[4097]),
			.SE(gen[4098]),

			.SELF(gen[4002]),
			.cell_state(gen[4002])
		); 

/******************* CELL 4003 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4003 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3907]),
			.N(gen[3908]),
			.NE(gen[3909]),

			.O(gen[4002]),
			.E(gen[4004]),

			.SO(gen[4097]),
			.S(gen[4098]),
			.SE(gen[4099]),

			.SELF(gen[4003]),
			.cell_state(gen[4003])
		); 

/******************* CELL 4004 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4004 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3908]),
			.N(gen[3909]),
			.NE(gen[3910]),

			.O(gen[4003]),
			.E(gen[4005]),

			.SO(gen[4098]),
			.S(gen[4099]),
			.SE(gen[4100]),

			.SELF(gen[4004]),
			.cell_state(gen[4004])
		); 

/******************* CELL 4005 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4005 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3909]),
			.N(gen[3910]),
			.NE(gen[3911]),

			.O(gen[4004]),
			.E(gen[4006]),

			.SO(gen[4099]),
			.S(gen[4100]),
			.SE(gen[4101]),

			.SELF(gen[4005]),
			.cell_state(gen[4005])
		); 

/******************* CELL 4006 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4006 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3910]),
			.N(gen[3911]),
			.NE(gen[3912]),

			.O(gen[4005]),
			.E(gen[4007]),

			.SO(gen[4100]),
			.S(gen[4101]),
			.SE(gen[4102]),

			.SELF(gen[4006]),
			.cell_state(gen[4006])
		); 

/******************* CELL 4007 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4007 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3911]),
			.N(gen[3912]),
			.NE(gen[3913]),

			.O(gen[4006]),
			.E(gen[4008]),

			.SO(gen[4101]),
			.S(gen[4102]),
			.SE(gen[4103]),

			.SELF(gen[4007]),
			.cell_state(gen[4007])
		); 

/******************* CELL 4008 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4008 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3912]),
			.N(gen[3913]),
			.NE(gen[3914]),

			.O(gen[4007]),
			.E(gen[4009]),

			.SO(gen[4102]),
			.S(gen[4103]),
			.SE(gen[4104]),

			.SELF(gen[4008]),
			.cell_state(gen[4008])
		); 

/******************* CELL 4009 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4009 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3913]),
			.N(gen[3914]),
			.NE(gen[3915]),

			.O(gen[4008]),
			.E(gen[4010]),

			.SO(gen[4103]),
			.S(gen[4104]),
			.SE(gen[4105]),

			.SELF(gen[4009]),
			.cell_state(gen[4009])
		); 

/******************* CELL 4010 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4010 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3914]),
			.N(gen[3915]),
			.NE(gen[3916]),

			.O(gen[4009]),
			.E(gen[4011]),

			.SO(gen[4104]),
			.S(gen[4105]),
			.SE(gen[4106]),

			.SELF(gen[4010]),
			.cell_state(gen[4010])
		); 

/******************* CELL 4011 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4011 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3915]),
			.N(gen[3916]),
			.NE(gen[3917]),

			.O(gen[4010]),
			.E(gen[4012]),

			.SO(gen[4105]),
			.S(gen[4106]),
			.SE(gen[4107]),

			.SELF(gen[4011]),
			.cell_state(gen[4011])
		); 

/******************* CELL 4012 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4012 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3916]),
			.N(gen[3917]),
			.NE(gen[3918]),

			.O(gen[4011]),
			.E(gen[4013]),

			.SO(gen[4106]),
			.S(gen[4107]),
			.SE(gen[4108]),

			.SELF(gen[4012]),
			.cell_state(gen[4012])
		); 

/******************* CELL 4013 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4013 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3917]),
			.N(gen[3918]),
			.NE(gen[3919]),

			.O(gen[4012]),
			.E(gen[4014]),

			.SO(gen[4107]),
			.S(gen[4108]),
			.SE(gen[4109]),

			.SELF(gen[4013]),
			.cell_state(gen[4013])
		); 

/******************* CELL 4014 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4014 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3918]),
			.N(gen[3919]),
			.NE(gen[3920]),

			.O(gen[4013]),
			.E(gen[4015]),

			.SO(gen[4108]),
			.S(gen[4109]),
			.SE(gen[4110]),

			.SELF(gen[4014]),
			.cell_state(gen[4014])
		); 

/******************* CELL 4015 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4015 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3919]),
			.N(gen[3920]),
			.NE(gen[3921]),

			.O(gen[4014]),
			.E(gen[4016]),

			.SO(gen[4109]),
			.S(gen[4110]),
			.SE(gen[4111]),

			.SELF(gen[4015]),
			.cell_state(gen[4015])
		); 

/******************* CELL 4016 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4016 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3920]),
			.N(gen[3921]),
			.NE(gen[3922]),

			.O(gen[4015]),
			.E(gen[4017]),

			.SO(gen[4110]),
			.S(gen[4111]),
			.SE(gen[4112]),

			.SELF(gen[4016]),
			.cell_state(gen[4016])
		); 

/******************* CELL 4017 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4017 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3921]),
			.N(gen[3922]),
			.NE(gen[3923]),

			.O(gen[4016]),
			.E(gen[4018]),

			.SO(gen[4111]),
			.S(gen[4112]),
			.SE(gen[4113]),

			.SELF(gen[4017]),
			.cell_state(gen[4017])
		); 

/******************* CELL 4018 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4018 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3922]),
			.N(gen[3923]),
			.NE(gen[3924]),

			.O(gen[4017]),
			.E(gen[4019]),

			.SO(gen[4112]),
			.S(gen[4113]),
			.SE(gen[4114]),

			.SELF(gen[4018]),
			.cell_state(gen[4018])
		); 

/******************* CELL 4019 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4019 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3923]),
			.N(gen[3924]),
			.NE(gen[3925]),

			.O(gen[4018]),
			.E(gen[4020]),

			.SO(gen[4113]),
			.S(gen[4114]),
			.SE(gen[4115]),

			.SELF(gen[4019]),
			.cell_state(gen[4019])
		); 

/******************* CELL 4020 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4020 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3924]),
			.N(gen[3925]),
			.NE(gen[3926]),

			.O(gen[4019]),
			.E(gen[4021]),

			.SO(gen[4114]),
			.S(gen[4115]),
			.SE(gen[4116]),

			.SELF(gen[4020]),
			.cell_state(gen[4020])
		); 

/******************* CELL 4021 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4021 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3925]),
			.N(gen[3926]),
			.NE(gen[3927]),

			.O(gen[4020]),
			.E(gen[4022]),

			.SO(gen[4115]),
			.S(gen[4116]),
			.SE(gen[4117]),

			.SELF(gen[4021]),
			.cell_state(gen[4021])
		); 

/******************* CELL 4022 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4022 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3926]),
			.N(gen[3927]),
			.NE(gen[3928]),

			.O(gen[4021]),
			.E(gen[4023]),

			.SO(gen[4116]),
			.S(gen[4117]),
			.SE(gen[4118]),

			.SELF(gen[4022]),
			.cell_state(gen[4022])
		); 

/******************* CELL 4023 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4023 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3927]),
			.N(gen[3928]),
			.NE(gen[3929]),

			.O(gen[4022]),
			.E(gen[4024]),

			.SO(gen[4117]),
			.S(gen[4118]),
			.SE(gen[4119]),

			.SELF(gen[4023]),
			.cell_state(gen[4023])
		); 

/******************* CELL 4024 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4024 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3928]),
			.N(gen[3929]),
			.NE(gen[3930]),

			.O(gen[4023]),
			.E(gen[4025]),

			.SO(gen[4118]),
			.S(gen[4119]),
			.SE(gen[4120]),

			.SELF(gen[4024]),
			.cell_state(gen[4024])
		); 

/******************* CELL 4025 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4025 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3929]),
			.N(gen[3930]),
			.NE(gen[3931]),

			.O(gen[4024]),
			.E(gen[4026]),

			.SO(gen[4119]),
			.S(gen[4120]),
			.SE(gen[4121]),

			.SELF(gen[4025]),
			.cell_state(gen[4025])
		); 

/******************* CELL 4026 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4026 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3930]),
			.N(gen[3931]),
			.NE(gen[3932]),

			.O(gen[4025]),
			.E(gen[4027]),

			.SO(gen[4120]),
			.S(gen[4121]),
			.SE(gen[4122]),

			.SELF(gen[4026]),
			.cell_state(gen[4026])
		); 

/******************* CELL 4027 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4027 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3931]),
			.N(gen[3932]),
			.NE(gen[3933]),

			.O(gen[4026]),
			.E(gen[4028]),

			.SO(gen[4121]),
			.S(gen[4122]),
			.SE(gen[4123]),

			.SELF(gen[4027]),
			.cell_state(gen[4027])
		); 

/******************* CELL 4028 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4028 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3932]),
			.N(gen[3933]),
			.NE(gen[3934]),

			.O(gen[4027]),
			.E(gen[4029]),

			.SO(gen[4122]),
			.S(gen[4123]),
			.SE(gen[4124]),

			.SELF(gen[4028]),
			.cell_state(gen[4028])
		); 

/******************* CELL 4029 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4029 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3933]),
			.N(gen[3934]),
			.NE(gen[3935]),

			.O(gen[4028]),
			.E(gen[4030]),

			.SO(gen[4123]),
			.S(gen[4124]),
			.SE(gen[4125]),

			.SELF(gen[4029]),
			.cell_state(gen[4029])
		); 

/******************* CELL 4030 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4030 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3934]),
			.N(gen[3935]),
			.NE(gen[3936]),

			.O(gen[4029]),
			.E(gen[4031]),

			.SO(gen[4124]),
			.S(gen[4125]),
			.SE(gen[4126]),

			.SELF(gen[4030]),
			.cell_state(gen[4030])
		); 

/******************* CELL 4031 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4031 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3935]),
			.N(gen[3936]),
			.NE(gen[3937]),

			.O(gen[4030]),
			.E(gen[4032]),

			.SO(gen[4125]),
			.S(gen[4126]),
			.SE(gen[4127]),

			.SELF(gen[4031]),
			.cell_state(gen[4031])
		); 

/******************* CELL 4032 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4032 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3936]),
			.N(gen[3937]),
			.NE(gen[3938]),

			.O(gen[4031]),
			.E(gen[4033]),

			.SO(gen[4126]),
			.S(gen[4127]),
			.SE(gen[4128]),

			.SELF(gen[4032]),
			.cell_state(gen[4032])
		); 

/******************* CELL 4033 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4033 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3937]),
			.N(gen[3938]),
			.NE(gen[3939]),

			.O(gen[4032]),
			.E(gen[4034]),

			.SO(gen[4127]),
			.S(gen[4128]),
			.SE(gen[4129]),

			.SELF(gen[4033]),
			.cell_state(gen[4033])
		); 

/******************* CELL 4034 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4034 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3938]),
			.N(gen[3939]),
			.NE(gen[3940]),

			.O(gen[4033]),
			.E(gen[4035]),

			.SO(gen[4128]),
			.S(gen[4129]),
			.SE(gen[4130]),

			.SELF(gen[4034]),
			.cell_state(gen[4034])
		); 

/******************* CELL 4035 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4035 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3939]),
			.N(gen[3940]),
			.NE(gen[3941]),

			.O(gen[4034]),
			.E(gen[4036]),

			.SO(gen[4129]),
			.S(gen[4130]),
			.SE(gen[4131]),

			.SELF(gen[4035]),
			.cell_state(gen[4035])
		); 

/******************* CELL 4036 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4036 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3940]),
			.N(gen[3941]),
			.NE(gen[3942]),

			.O(gen[4035]),
			.E(gen[4037]),

			.SO(gen[4130]),
			.S(gen[4131]),
			.SE(gen[4132]),

			.SELF(gen[4036]),
			.cell_state(gen[4036])
		); 

/******************* CELL 4037 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4037 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3941]),
			.N(gen[3942]),
			.NE(gen[3943]),

			.O(gen[4036]),
			.E(gen[4038]),

			.SO(gen[4131]),
			.S(gen[4132]),
			.SE(gen[4133]),

			.SELF(gen[4037]),
			.cell_state(gen[4037])
		); 

/******************* CELL 4038 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4038 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3942]),
			.N(gen[3943]),
			.NE(gen[3944]),

			.O(gen[4037]),
			.E(gen[4039]),

			.SO(gen[4132]),
			.S(gen[4133]),
			.SE(gen[4134]),

			.SELF(gen[4038]),
			.cell_state(gen[4038])
		); 

/******************* CELL 4039 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4039 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3943]),
			.N(gen[3944]),
			.NE(gen[3945]),

			.O(gen[4038]),
			.E(gen[4040]),

			.SO(gen[4133]),
			.S(gen[4134]),
			.SE(gen[4135]),

			.SELF(gen[4039]),
			.cell_state(gen[4039])
		); 

/******************* CELL 4040 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4040 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3944]),
			.N(gen[3945]),
			.NE(gen[3946]),

			.O(gen[4039]),
			.E(gen[4041]),

			.SO(gen[4134]),
			.S(gen[4135]),
			.SE(gen[4136]),

			.SELF(gen[4040]),
			.cell_state(gen[4040])
		); 

/******************* CELL 4041 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4041 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3945]),
			.N(gen[3946]),
			.NE(gen[3947]),

			.O(gen[4040]),
			.E(gen[4042]),

			.SO(gen[4135]),
			.S(gen[4136]),
			.SE(gen[4137]),

			.SELF(gen[4041]),
			.cell_state(gen[4041])
		); 

/******************* CELL 4042 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4042 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3946]),
			.N(gen[3947]),
			.NE(gen[3948]),

			.O(gen[4041]),
			.E(gen[4043]),

			.SO(gen[4136]),
			.S(gen[4137]),
			.SE(gen[4138]),

			.SELF(gen[4042]),
			.cell_state(gen[4042])
		); 

/******************* CELL 4043 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4043 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3947]),
			.N(gen[3948]),
			.NE(gen[3949]),

			.O(gen[4042]),
			.E(gen[4044]),

			.SO(gen[4137]),
			.S(gen[4138]),
			.SE(gen[4139]),

			.SELF(gen[4043]),
			.cell_state(gen[4043])
		); 

/******************* CELL 4044 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4044 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3948]),
			.N(gen[3949]),
			.NE(gen[3950]),

			.O(gen[4043]),
			.E(gen[4045]),

			.SO(gen[4138]),
			.S(gen[4139]),
			.SE(gen[4140]),

			.SELF(gen[4044]),
			.cell_state(gen[4044])
		); 

/******************* CELL 4045 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4045 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3949]),
			.N(gen[3950]),
			.NE(gen[3951]),

			.O(gen[4044]),
			.E(gen[4046]),

			.SO(gen[4139]),
			.S(gen[4140]),
			.SE(gen[4141]),

			.SELF(gen[4045]),
			.cell_state(gen[4045])
		); 

/******************* CELL 4046 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4046 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3950]),
			.N(gen[3951]),
			.NE(gen[3952]),

			.O(gen[4045]),
			.E(gen[4047]),

			.SO(gen[4140]),
			.S(gen[4141]),
			.SE(gen[4142]),

			.SELF(gen[4046]),
			.cell_state(gen[4046])
		); 

/******************* CELL 4047 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4047 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3951]),
			.N(gen[3952]),
			.NE(gen[3953]),

			.O(gen[4046]),
			.E(gen[4048]),

			.SO(gen[4141]),
			.S(gen[4142]),
			.SE(gen[4143]),

			.SELF(gen[4047]),
			.cell_state(gen[4047])
		); 

/******************* CELL 4048 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4048 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3952]),
			.N(gen[3953]),
			.NE(gen[3954]),

			.O(gen[4047]),
			.E(gen[4049]),

			.SO(gen[4142]),
			.S(gen[4143]),
			.SE(gen[4144]),

			.SELF(gen[4048]),
			.cell_state(gen[4048])
		); 

/******************* CELL 4049 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4049 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3953]),
			.N(gen[3954]),
			.NE(gen[3955]),

			.O(gen[4048]),
			.E(gen[4050]),

			.SO(gen[4143]),
			.S(gen[4144]),
			.SE(gen[4145]),

			.SELF(gen[4049]),
			.cell_state(gen[4049])
		); 

/******************* CELL 4050 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4050 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3954]),
			.N(gen[3955]),
			.NE(gen[3956]),

			.O(gen[4049]),
			.E(gen[4051]),

			.SO(gen[4144]),
			.S(gen[4145]),
			.SE(gen[4146]),

			.SELF(gen[4050]),
			.cell_state(gen[4050])
		); 

/******************* CELL 4051 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4051 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3955]),
			.N(gen[3956]),
			.NE(gen[3957]),

			.O(gen[4050]),
			.E(gen[4052]),

			.SO(gen[4145]),
			.S(gen[4146]),
			.SE(gen[4147]),

			.SELF(gen[4051]),
			.cell_state(gen[4051])
		); 

/******************* CELL 4052 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4052 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3956]),
			.N(gen[3957]),
			.NE(gen[3958]),

			.O(gen[4051]),
			.E(gen[4053]),

			.SO(gen[4146]),
			.S(gen[4147]),
			.SE(gen[4148]),

			.SELF(gen[4052]),
			.cell_state(gen[4052])
		); 

/******************* CELL 4053 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4053 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3957]),
			.N(gen[3958]),
			.NE(gen[3959]),

			.O(gen[4052]),
			.E(gen[4054]),

			.SO(gen[4147]),
			.S(gen[4148]),
			.SE(gen[4149]),

			.SELF(gen[4053]),
			.cell_state(gen[4053])
		); 

/******************* CELL 4054 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4054 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3958]),
			.N(gen[3959]),
			.NE(gen[3960]),

			.O(gen[4053]),
			.E(gen[4055]),

			.SO(gen[4148]),
			.S(gen[4149]),
			.SE(gen[4150]),

			.SELF(gen[4054]),
			.cell_state(gen[4054])
		); 

/******************* CELL 4055 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4055 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3959]),
			.N(gen[3960]),
			.NE(gen[3961]),

			.O(gen[4054]),
			.E(gen[4056]),

			.SO(gen[4149]),
			.S(gen[4150]),
			.SE(gen[4151]),

			.SELF(gen[4055]),
			.cell_state(gen[4055])
		); 

/******************* CELL 4056 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4056 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3960]),
			.N(gen[3961]),
			.NE(gen[3962]),

			.O(gen[4055]),
			.E(gen[4057]),

			.SO(gen[4150]),
			.S(gen[4151]),
			.SE(gen[4152]),

			.SELF(gen[4056]),
			.cell_state(gen[4056])
		); 

/******************* CELL 4057 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4057 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3961]),
			.N(gen[3962]),
			.NE(gen[3963]),

			.O(gen[4056]),
			.E(gen[4058]),

			.SO(gen[4151]),
			.S(gen[4152]),
			.SE(gen[4153]),

			.SELF(gen[4057]),
			.cell_state(gen[4057])
		); 

/******************* CELL 4058 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4058 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3962]),
			.N(gen[3963]),
			.NE(gen[3964]),

			.O(gen[4057]),
			.E(gen[4059]),

			.SO(gen[4152]),
			.S(gen[4153]),
			.SE(gen[4154]),

			.SELF(gen[4058]),
			.cell_state(gen[4058])
		); 

/******************* CELL 4059 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4059 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3963]),
			.N(gen[3964]),
			.NE(gen[3965]),

			.O(gen[4058]),
			.E(gen[4060]),

			.SO(gen[4153]),
			.S(gen[4154]),
			.SE(gen[4155]),

			.SELF(gen[4059]),
			.cell_state(gen[4059])
		); 

/******************* CELL 4060 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4060 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3964]),
			.N(gen[3965]),
			.NE(gen[3966]),

			.O(gen[4059]),
			.E(gen[4061]),

			.SO(gen[4154]),
			.S(gen[4155]),
			.SE(gen[4156]),

			.SELF(gen[4060]),
			.cell_state(gen[4060])
		); 

/******************* CELL 4061 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4061 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3965]),
			.N(gen[3966]),
			.NE(gen[3967]),

			.O(gen[4060]),
			.E(gen[4062]),

			.SO(gen[4155]),
			.S(gen[4156]),
			.SE(gen[4157]),

			.SELF(gen[4061]),
			.cell_state(gen[4061])
		); 

/******************* CELL 4062 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4062 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3966]),
			.N(gen[3967]),
			.NE(gen[3968]),

			.O(gen[4061]),
			.E(gen[4063]),

			.SO(gen[4156]),
			.S(gen[4157]),
			.SE(gen[4158]),

			.SELF(gen[4062]),
			.cell_state(gen[4062])
		); 

/******************* CELL 4063 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4063 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3967]),
			.N(gen[3968]),
			.NE(gen[3969]),

			.O(gen[4062]),
			.E(gen[4064]),

			.SO(gen[4157]),
			.S(gen[4158]),
			.SE(gen[4159]),

			.SELF(gen[4063]),
			.cell_state(gen[4063])
		); 

/******************* CELL 4064 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4064 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3968]),
			.N(gen[3969]),
			.NE(gen[3970]),

			.O(gen[4063]),
			.E(gen[4065]),

			.SO(gen[4158]),
			.S(gen[4159]),
			.SE(gen[4160]),

			.SELF(gen[4064]),
			.cell_state(gen[4064])
		); 

/******************* CELL 4065 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4065 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3969]),
			.N(gen[3970]),
			.NE(gen[3971]),

			.O(gen[4064]),
			.E(gen[4066]),

			.SO(gen[4159]),
			.S(gen[4160]),
			.SE(gen[4161]),

			.SELF(gen[4065]),
			.cell_state(gen[4065])
		); 

/******************* CELL 4066 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4066 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3970]),
			.N(gen[3971]),
			.NE(gen[3972]),

			.O(gen[4065]),
			.E(gen[4067]),

			.SO(gen[4160]),
			.S(gen[4161]),
			.SE(gen[4162]),

			.SELF(gen[4066]),
			.cell_state(gen[4066])
		); 

/******************* CELL 4067 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4067 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3971]),
			.N(gen[3972]),
			.NE(gen[3973]),

			.O(gen[4066]),
			.E(gen[4068]),

			.SO(gen[4161]),
			.S(gen[4162]),
			.SE(gen[4163]),

			.SELF(gen[4067]),
			.cell_state(gen[4067])
		); 

/******************* CELL 4068 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4068 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3972]),
			.N(gen[3973]),
			.NE(gen[3974]),

			.O(gen[4067]),
			.E(gen[4069]),

			.SO(gen[4162]),
			.S(gen[4163]),
			.SE(gen[4164]),

			.SELF(gen[4068]),
			.cell_state(gen[4068])
		); 

/******************* CELL 4069 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4069 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3973]),
			.N(gen[3974]),
			.NE(gen[3975]),

			.O(gen[4068]),
			.E(gen[4070]),

			.SO(gen[4163]),
			.S(gen[4164]),
			.SE(gen[4165]),

			.SELF(gen[4069]),
			.cell_state(gen[4069])
		); 

/******************* CELL 4070 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4070 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3974]),
			.N(gen[3975]),
			.NE(gen[3976]),

			.O(gen[4069]),
			.E(gen[4071]),

			.SO(gen[4164]),
			.S(gen[4165]),
			.SE(gen[4166]),

			.SELF(gen[4070]),
			.cell_state(gen[4070])
		); 

/******************* CELL 4071 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4071 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3975]),
			.N(gen[3976]),
			.NE(gen[3977]),

			.O(gen[4070]),
			.E(gen[4072]),

			.SO(gen[4165]),
			.S(gen[4166]),
			.SE(gen[4167]),

			.SELF(gen[4071]),
			.cell_state(gen[4071])
		); 

/******************* CELL 4072 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4072 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3976]),
			.N(gen[3977]),
			.NE(gen[3978]),

			.O(gen[4071]),
			.E(gen[4073]),

			.SO(gen[4166]),
			.S(gen[4167]),
			.SE(gen[4168]),

			.SELF(gen[4072]),
			.cell_state(gen[4072])
		); 

/******************* CELL 4073 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4073 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3977]),
			.N(gen[3978]),
			.NE(gen[3979]),

			.O(gen[4072]),
			.E(gen[4074]),

			.SO(gen[4167]),
			.S(gen[4168]),
			.SE(gen[4169]),

			.SELF(gen[4073]),
			.cell_state(gen[4073])
		); 

/******************* CELL 4074 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4074 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3978]),
			.N(gen[3979]),
			.NE(gen[3980]),

			.O(gen[4073]),
			.E(gen[4075]),

			.SO(gen[4168]),
			.S(gen[4169]),
			.SE(gen[4170]),

			.SELF(gen[4074]),
			.cell_state(gen[4074])
		); 

/******************* CELL 4075 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4075 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3979]),
			.N(gen[3980]),
			.NE(gen[3981]),

			.O(gen[4074]),
			.E(gen[4076]),

			.SO(gen[4169]),
			.S(gen[4170]),
			.SE(gen[4171]),

			.SELF(gen[4075]),
			.cell_state(gen[4075])
		); 

/******************* CELL 4076 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4076 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3980]),
			.N(gen[3981]),
			.NE(gen[3982]),

			.O(gen[4075]),
			.E(gen[4077]),

			.SO(gen[4170]),
			.S(gen[4171]),
			.SE(gen[4172]),

			.SELF(gen[4076]),
			.cell_state(gen[4076])
		); 

/******************* CELL 4077 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4077 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3981]),
			.N(gen[3982]),
			.NE(gen[3983]),

			.O(gen[4076]),
			.E(gen[4078]),

			.SO(gen[4171]),
			.S(gen[4172]),
			.SE(gen[4173]),

			.SELF(gen[4077]),
			.cell_state(gen[4077])
		); 

/******************* CELL 4078 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4078 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3982]),
			.N(gen[3983]),
			.NE(gen[3984]),

			.O(gen[4077]),
			.E(gen[4079]),

			.SO(gen[4172]),
			.S(gen[4173]),
			.SE(gen[4174]),

			.SELF(gen[4078]),
			.cell_state(gen[4078])
		); 

/******************* CELL 4079 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4079 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3983]),
			.N(gen[3984]),
			.NE(gen[3985]),

			.O(gen[4078]),
			.E(gen[4080]),

			.SO(gen[4173]),
			.S(gen[4174]),
			.SE(gen[4175]),

			.SELF(gen[4079]),
			.cell_state(gen[4079])
		); 

/******************* CELL 4080 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4080 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3984]),
			.N(gen[3985]),
			.NE(gen[3986]),

			.O(gen[4079]),
			.E(gen[4081]),

			.SO(gen[4174]),
			.S(gen[4175]),
			.SE(gen[4176]),

			.SELF(gen[4080]),
			.cell_state(gen[4080])
		); 

/******************* CELL 4081 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4081 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3985]),
			.N(gen[3986]),
			.NE(gen[3987]),

			.O(gen[4080]),
			.E(gen[4082]),

			.SO(gen[4175]),
			.S(gen[4176]),
			.SE(gen[4177]),

			.SELF(gen[4081]),
			.cell_state(gen[4081])
		); 

/******************* CELL 4082 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4082 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3986]),
			.N(gen[3987]),
			.NE(gen[3988]),

			.O(gen[4081]),
			.E(gen[4083]),

			.SO(gen[4176]),
			.S(gen[4177]),
			.SE(gen[4178]),

			.SELF(gen[4082]),
			.cell_state(gen[4082])
		); 

/******************* CELL 4083 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4083 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3987]),
			.N(gen[3988]),
			.NE(gen[3989]),

			.O(gen[4082]),
			.E(gen[4084]),

			.SO(gen[4177]),
			.S(gen[4178]),
			.SE(gen[4179]),

			.SELF(gen[4083]),
			.cell_state(gen[4083])
		); 

/******************* CELL 4084 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4084 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3988]),
			.N(gen[3989]),
			.NE(gen[3988]),

			.O(gen[4083]),
			.E(gen[4083]),

			.SO(gen[4178]),
			.S(gen[4179]),
			.SE(gen[4178]),

			.SELF(gen[4084]),
			.cell_state(gen[4084])
		); 

/******************* CELL 4085 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4085 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3991]),
			.N(gen[3990]),
			.NE(gen[3991]),

			.O(gen[4086]),
			.E(gen[4086]),

			.SO(gen[4181]),
			.S(gen[4180]),
			.SE(gen[4181]),

			.SELF(gen[4085]),
			.cell_state(gen[4085])
		); 

/******************* CELL 4086 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4086 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3990]),
			.N(gen[3991]),
			.NE(gen[3992]),

			.O(gen[4085]),
			.E(gen[4087]),

			.SO(gen[4180]),
			.S(gen[4181]),
			.SE(gen[4182]),

			.SELF(gen[4086]),
			.cell_state(gen[4086])
		); 

/******************* CELL 4087 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4087 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3991]),
			.N(gen[3992]),
			.NE(gen[3993]),

			.O(gen[4086]),
			.E(gen[4088]),

			.SO(gen[4181]),
			.S(gen[4182]),
			.SE(gen[4183]),

			.SELF(gen[4087]),
			.cell_state(gen[4087])
		); 

/******************* CELL 4088 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4088 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3992]),
			.N(gen[3993]),
			.NE(gen[3994]),

			.O(gen[4087]),
			.E(gen[4089]),

			.SO(gen[4182]),
			.S(gen[4183]),
			.SE(gen[4184]),

			.SELF(gen[4088]),
			.cell_state(gen[4088])
		); 

/******************* CELL 4089 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4089 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3993]),
			.N(gen[3994]),
			.NE(gen[3995]),

			.O(gen[4088]),
			.E(gen[4090]),

			.SO(gen[4183]),
			.S(gen[4184]),
			.SE(gen[4185]),

			.SELF(gen[4089]),
			.cell_state(gen[4089])
		); 

/******************* CELL 4090 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4090 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3994]),
			.N(gen[3995]),
			.NE(gen[3996]),

			.O(gen[4089]),
			.E(gen[4091]),

			.SO(gen[4184]),
			.S(gen[4185]),
			.SE(gen[4186]),

			.SELF(gen[4090]),
			.cell_state(gen[4090])
		); 

/******************* CELL 4091 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4091 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3995]),
			.N(gen[3996]),
			.NE(gen[3997]),

			.O(gen[4090]),
			.E(gen[4092]),

			.SO(gen[4185]),
			.S(gen[4186]),
			.SE(gen[4187]),

			.SELF(gen[4091]),
			.cell_state(gen[4091])
		); 

/******************* CELL 4092 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4092 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3996]),
			.N(gen[3997]),
			.NE(gen[3998]),

			.O(gen[4091]),
			.E(gen[4093]),

			.SO(gen[4186]),
			.S(gen[4187]),
			.SE(gen[4188]),

			.SELF(gen[4092]),
			.cell_state(gen[4092])
		); 

/******************* CELL 4093 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4093 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3997]),
			.N(gen[3998]),
			.NE(gen[3999]),

			.O(gen[4092]),
			.E(gen[4094]),

			.SO(gen[4187]),
			.S(gen[4188]),
			.SE(gen[4189]),

			.SELF(gen[4093]),
			.cell_state(gen[4093])
		); 

/******************* CELL 4094 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4094 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3998]),
			.N(gen[3999]),
			.NE(gen[4000]),

			.O(gen[4093]),
			.E(gen[4095]),

			.SO(gen[4188]),
			.S(gen[4189]),
			.SE(gen[4190]),

			.SELF(gen[4094]),
			.cell_state(gen[4094])
		); 

/******************* CELL 4095 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4095 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3999]),
			.N(gen[4000]),
			.NE(gen[4001]),

			.O(gen[4094]),
			.E(gen[4096]),

			.SO(gen[4189]),
			.S(gen[4190]),
			.SE(gen[4191]),

			.SELF(gen[4095]),
			.cell_state(gen[4095])
		); 

/******************* CELL 4096 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4096 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4000]),
			.N(gen[4001]),
			.NE(gen[4002]),

			.O(gen[4095]),
			.E(gen[4097]),

			.SO(gen[4190]),
			.S(gen[4191]),
			.SE(gen[4192]),

			.SELF(gen[4096]),
			.cell_state(gen[4096])
		); 

/******************* CELL 4097 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4097 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4001]),
			.N(gen[4002]),
			.NE(gen[4003]),

			.O(gen[4096]),
			.E(gen[4098]),

			.SO(gen[4191]),
			.S(gen[4192]),
			.SE(gen[4193]),

			.SELF(gen[4097]),
			.cell_state(gen[4097])
		); 

/******************* CELL 4098 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4098 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4002]),
			.N(gen[4003]),
			.NE(gen[4004]),

			.O(gen[4097]),
			.E(gen[4099]),

			.SO(gen[4192]),
			.S(gen[4193]),
			.SE(gen[4194]),

			.SELF(gen[4098]),
			.cell_state(gen[4098])
		); 

/******************* CELL 4099 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4099 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4003]),
			.N(gen[4004]),
			.NE(gen[4005]),

			.O(gen[4098]),
			.E(gen[4100]),

			.SO(gen[4193]),
			.S(gen[4194]),
			.SE(gen[4195]),

			.SELF(gen[4099]),
			.cell_state(gen[4099])
		); 

/******************* CELL 4100 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4100 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4004]),
			.N(gen[4005]),
			.NE(gen[4006]),

			.O(gen[4099]),
			.E(gen[4101]),

			.SO(gen[4194]),
			.S(gen[4195]),
			.SE(gen[4196]),

			.SELF(gen[4100]),
			.cell_state(gen[4100])
		); 

/******************* CELL 4101 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4101 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4005]),
			.N(gen[4006]),
			.NE(gen[4007]),

			.O(gen[4100]),
			.E(gen[4102]),

			.SO(gen[4195]),
			.S(gen[4196]),
			.SE(gen[4197]),

			.SELF(gen[4101]),
			.cell_state(gen[4101])
		); 

/******************* CELL 4102 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4102 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4006]),
			.N(gen[4007]),
			.NE(gen[4008]),

			.O(gen[4101]),
			.E(gen[4103]),

			.SO(gen[4196]),
			.S(gen[4197]),
			.SE(gen[4198]),

			.SELF(gen[4102]),
			.cell_state(gen[4102])
		); 

/******************* CELL 4103 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4103 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4007]),
			.N(gen[4008]),
			.NE(gen[4009]),

			.O(gen[4102]),
			.E(gen[4104]),

			.SO(gen[4197]),
			.S(gen[4198]),
			.SE(gen[4199]),

			.SELF(gen[4103]),
			.cell_state(gen[4103])
		); 

/******************* CELL 4104 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4104 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4008]),
			.N(gen[4009]),
			.NE(gen[4010]),

			.O(gen[4103]),
			.E(gen[4105]),

			.SO(gen[4198]),
			.S(gen[4199]),
			.SE(gen[4200]),

			.SELF(gen[4104]),
			.cell_state(gen[4104])
		); 

/******************* CELL 4105 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4105 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4009]),
			.N(gen[4010]),
			.NE(gen[4011]),

			.O(gen[4104]),
			.E(gen[4106]),

			.SO(gen[4199]),
			.S(gen[4200]),
			.SE(gen[4201]),

			.SELF(gen[4105]),
			.cell_state(gen[4105])
		); 

/******************* CELL 4106 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4106 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4010]),
			.N(gen[4011]),
			.NE(gen[4012]),

			.O(gen[4105]),
			.E(gen[4107]),

			.SO(gen[4200]),
			.S(gen[4201]),
			.SE(gen[4202]),

			.SELF(gen[4106]),
			.cell_state(gen[4106])
		); 

/******************* CELL 4107 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4107 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4011]),
			.N(gen[4012]),
			.NE(gen[4013]),

			.O(gen[4106]),
			.E(gen[4108]),

			.SO(gen[4201]),
			.S(gen[4202]),
			.SE(gen[4203]),

			.SELF(gen[4107]),
			.cell_state(gen[4107])
		); 

/******************* CELL 4108 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4108 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4012]),
			.N(gen[4013]),
			.NE(gen[4014]),

			.O(gen[4107]),
			.E(gen[4109]),

			.SO(gen[4202]),
			.S(gen[4203]),
			.SE(gen[4204]),

			.SELF(gen[4108]),
			.cell_state(gen[4108])
		); 

/******************* CELL 4109 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4109 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4013]),
			.N(gen[4014]),
			.NE(gen[4015]),

			.O(gen[4108]),
			.E(gen[4110]),

			.SO(gen[4203]),
			.S(gen[4204]),
			.SE(gen[4205]),

			.SELF(gen[4109]),
			.cell_state(gen[4109])
		); 

/******************* CELL 4110 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4110 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4014]),
			.N(gen[4015]),
			.NE(gen[4016]),

			.O(gen[4109]),
			.E(gen[4111]),

			.SO(gen[4204]),
			.S(gen[4205]),
			.SE(gen[4206]),

			.SELF(gen[4110]),
			.cell_state(gen[4110])
		); 

/******************* CELL 4111 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4111 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4015]),
			.N(gen[4016]),
			.NE(gen[4017]),

			.O(gen[4110]),
			.E(gen[4112]),

			.SO(gen[4205]),
			.S(gen[4206]),
			.SE(gen[4207]),

			.SELF(gen[4111]),
			.cell_state(gen[4111])
		); 

/******************* CELL 4112 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4112 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4016]),
			.N(gen[4017]),
			.NE(gen[4018]),

			.O(gen[4111]),
			.E(gen[4113]),

			.SO(gen[4206]),
			.S(gen[4207]),
			.SE(gen[4208]),

			.SELF(gen[4112]),
			.cell_state(gen[4112])
		); 

/******************* CELL 4113 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4113 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4017]),
			.N(gen[4018]),
			.NE(gen[4019]),

			.O(gen[4112]),
			.E(gen[4114]),

			.SO(gen[4207]),
			.S(gen[4208]),
			.SE(gen[4209]),

			.SELF(gen[4113]),
			.cell_state(gen[4113])
		); 

/******************* CELL 4114 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4114 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4018]),
			.N(gen[4019]),
			.NE(gen[4020]),

			.O(gen[4113]),
			.E(gen[4115]),

			.SO(gen[4208]),
			.S(gen[4209]),
			.SE(gen[4210]),

			.SELF(gen[4114]),
			.cell_state(gen[4114])
		); 

/******************* CELL 4115 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4115 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4019]),
			.N(gen[4020]),
			.NE(gen[4021]),

			.O(gen[4114]),
			.E(gen[4116]),

			.SO(gen[4209]),
			.S(gen[4210]),
			.SE(gen[4211]),

			.SELF(gen[4115]),
			.cell_state(gen[4115])
		); 

/******************* CELL 4116 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4116 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4020]),
			.N(gen[4021]),
			.NE(gen[4022]),

			.O(gen[4115]),
			.E(gen[4117]),

			.SO(gen[4210]),
			.S(gen[4211]),
			.SE(gen[4212]),

			.SELF(gen[4116]),
			.cell_state(gen[4116])
		); 

/******************* CELL 4117 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4117 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4021]),
			.N(gen[4022]),
			.NE(gen[4023]),

			.O(gen[4116]),
			.E(gen[4118]),

			.SO(gen[4211]),
			.S(gen[4212]),
			.SE(gen[4213]),

			.SELF(gen[4117]),
			.cell_state(gen[4117])
		); 

/******************* CELL 4118 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4118 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4022]),
			.N(gen[4023]),
			.NE(gen[4024]),

			.O(gen[4117]),
			.E(gen[4119]),

			.SO(gen[4212]),
			.S(gen[4213]),
			.SE(gen[4214]),

			.SELF(gen[4118]),
			.cell_state(gen[4118])
		); 

/******************* CELL 4119 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4119 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4023]),
			.N(gen[4024]),
			.NE(gen[4025]),

			.O(gen[4118]),
			.E(gen[4120]),

			.SO(gen[4213]),
			.S(gen[4214]),
			.SE(gen[4215]),

			.SELF(gen[4119]),
			.cell_state(gen[4119])
		); 

/******************* CELL 4120 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4120 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4024]),
			.N(gen[4025]),
			.NE(gen[4026]),

			.O(gen[4119]),
			.E(gen[4121]),

			.SO(gen[4214]),
			.S(gen[4215]),
			.SE(gen[4216]),

			.SELF(gen[4120]),
			.cell_state(gen[4120])
		); 

/******************* CELL 4121 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4121 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4025]),
			.N(gen[4026]),
			.NE(gen[4027]),

			.O(gen[4120]),
			.E(gen[4122]),

			.SO(gen[4215]),
			.S(gen[4216]),
			.SE(gen[4217]),

			.SELF(gen[4121]),
			.cell_state(gen[4121])
		); 

/******************* CELL 4122 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4122 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4026]),
			.N(gen[4027]),
			.NE(gen[4028]),

			.O(gen[4121]),
			.E(gen[4123]),

			.SO(gen[4216]),
			.S(gen[4217]),
			.SE(gen[4218]),

			.SELF(gen[4122]),
			.cell_state(gen[4122])
		); 

/******************* CELL 4123 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4123 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4027]),
			.N(gen[4028]),
			.NE(gen[4029]),

			.O(gen[4122]),
			.E(gen[4124]),

			.SO(gen[4217]),
			.S(gen[4218]),
			.SE(gen[4219]),

			.SELF(gen[4123]),
			.cell_state(gen[4123])
		); 

/******************* CELL 4124 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4124 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4028]),
			.N(gen[4029]),
			.NE(gen[4030]),

			.O(gen[4123]),
			.E(gen[4125]),

			.SO(gen[4218]),
			.S(gen[4219]),
			.SE(gen[4220]),

			.SELF(gen[4124]),
			.cell_state(gen[4124])
		); 

/******************* CELL 4125 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4125 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4029]),
			.N(gen[4030]),
			.NE(gen[4031]),

			.O(gen[4124]),
			.E(gen[4126]),

			.SO(gen[4219]),
			.S(gen[4220]),
			.SE(gen[4221]),

			.SELF(gen[4125]),
			.cell_state(gen[4125])
		); 

/******************* CELL 4126 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4126 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4030]),
			.N(gen[4031]),
			.NE(gen[4032]),

			.O(gen[4125]),
			.E(gen[4127]),

			.SO(gen[4220]),
			.S(gen[4221]),
			.SE(gen[4222]),

			.SELF(gen[4126]),
			.cell_state(gen[4126])
		); 

/******************* CELL 4127 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4127 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4031]),
			.N(gen[4032]),
			.NE(gen[4033]),

			.O(gen[4126]),
			.E(gen[4128]),

			.SO(gen[4221]),
			.S(gen[4222]),
			.SE(gen[4223]),

			.SELF(gen[4127]),
			.cell_state(gen[4127])
		); 

/******************* CELL 4128 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4128 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4032]),
			.N(gen[4033]),
			.NE(gen[4034]),

			.O(gen[4127]),
			.E(gen[4129]),

			.SO(gen[4222]),
			.S(gen[4223]),
			.SE(gen[4224]),

			.SELF(gen[4128]),
			.cell_state(gen[4128])
		); 

/******************* CELL 4129 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4129 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4033]),
			.N(gen[4034]),
			.NE(gen[4035]),

			.O(gen[4128]),
			.E(gen[4130]),

			.SO(gen[4223]),
			.S(gen[4224]),
			.SE(gen[4225]),

			.SELF(gen[4129]),
			.cell_state(gen[4129])
		); 

/******************* CELL 4130 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4130 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4034]),
			.N(gen[4035]),
			.NE(gen[4036]),

			.O(gen[4129]),
			.E(gen[4131]),

			.SO(gen[4224]),
			.S(gen[4225]),
			.SE(gen[4226]),

			.SELF(gen[4130]),
			.cell_state(gen[4130])
		); 

/******************* CELL 4131 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4131 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4035]),
			.N(gen[4036]),
			.NE(gen[4037]),

			.O(gen[4130]),
			.E(gen[4132]),

			.SO(gen[4225]),
			.S(gen[4226]),
			.SE(gen[4227]),

			.SELF(gen[4131]),
			.cell_state(gen[4131])
		); 

/******************* CELL 4132 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4132 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4036]),
			.N(gen[4037]),
			.NE(gen[4038]),

			.O(gen[4131]),
			.E(gen[4133]),

			.SO(gen[4226]),
			.S(gen[4227]),
			.SE(gen[4228]),

			.SELF(gen[4132]),
			.cell_state(gen[4132])
		); 

/******************* CELL 4133 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4133 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4037]),
			.N(gen[4038]),
			.NE(gen[4039]),

			.O(gen[4132]),
			.E(gen[4134]),

			.SO(gen[4227]),
			.S(gen[4228]),
			.SE(gen[4229]),

			.SELF(gen[4133]),
			.cell_state(gen[4133])
		); 

/******************* CELL 4134 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4134 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4038]),
			.N(gen[4039]),
			.NE(gen[4040]),

			.O(gen[4133]),
			.E(gen[4135]),

			.SO(gen[4228]),
			.S(gen[4229]),
			.SE(gen[4230]),

			.SELF(gen[4134]),
			.cell_state(gen[4134])
		); 

/******************* CELL 4135 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4135 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4039]),
			.N(gen[4040]),
			.NE(gen[4041]),

			.O(gen[4134]),
			.E(gen[4136]),

			.SO(gen[4229]),
			.S(gen[4230]),
			.SE(gen[4231]),

			.SELF(gen[4135]),
			.cell_state(gen[4135])
		); 

/******************* CELL 4136 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4136 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4040]),
			.N(gen[4041]),
			.NE(gen[4042]),

			.O(gen[4135]),
			.E(gen[4137]),

			.SO(gen[4230]),
			.S(gen[4231]),
			.SE(gen[4232]),

			.SELF(gen[4136]),
			.cell_state(gen[4136])
		); 

/******************* CELL 4137 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4137 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4041]),
			.N(gen[4042]),
			.NE(gen[4043]),

			.O(gen[4136]),
			.E(gen[4138]),

			.SO(gen[4231]),
			.S(gen[4232]),
			.SE(gen[4233]),

			.SELF(gen[4137]),
			.cell_state(gen[4137])
		); 

/******************* CELL 4138 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4138 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4042]),
			.N(gen[4043]),
			.NE(gen[4044]),

			.O(gen[4137]),
			.E(gen[4139]),

			.SO(gen[4232]),
			.S(gen[4233]),
			.SE(gen[4234]),

			.SELF(gen[4138]),
			.cell_state(gen[4138])
		); 

/******************* CELL 4139 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4139 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4043]),
			.N(gen[4044]),
			.NE(gen[4045]),

			.O(gen[4138]),
			.E(gen[4140]),

			.SO(gen[4233]),
			.S(gen[4234]),
			.SE(gen[4235]),

			.SELF(gen[4139]),
			.cell_state(gen[4139])
		); 

/******************* CELL 4140 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4140 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4044]),
			.N(gen[4045]),
			.NE(gen[4046]),

			.O(gen[4139]),
			.E(gen[4141]),

			.SO(gen[4234]),
			.S(gen[4235]),
			.SE(gen[4236]),

			.SELF(gen[4140]),
			.cell_state(gen[4140])
		); 

/******************* CELL 4141 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4141 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4045]),
			.N(gen[4046]),
			.NE(gen[4047]),

			.O(gen[4140]),
			.E(gen[4142]),

			.SO(gen[4235]),
			.S(gen[4236]),
			.SE(gen[4237]),

			.SELF(gen[4141]),
			.cell_state(gen[4141])
		); 

/******************* CELL 4142 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4142 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4046]),
			.N(gen[4047]),
			.NE(gen[4048]),

			.O(gen[4141]),
			.E(gen[4143]),

			.SO(gen[4236]),
			.S(gen[4237]),
			.SE(gen[4238]),

			.SELF(gen[4142]),
			.cell_state(gen[4142])
		); 

/******************* CELL 4143 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4143 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4047]),
			.N(gen[4048]),
			.NE(gen[4049]),

			.O(gen[4142]),
			.E(gen[4144]),

			.SO(gen[4237]),
			.S(gen[4238]),
			.SE(gen[4239]),

			.SELF(gen[4143]),
			.cell_state(gen[4143])
		); 

/******************* CELL 4144 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4144 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4048]),
			.N(gen[4049]),
			.NE(gen[4050]),

			.O(gen[4143]),
			.E(gen[4145]),

			.SO(gen[4238]),
			.S(gen[4239]),
			.SE(gen[4240]),

			.SELF(gen[4144]),
			.cell_state(gen[4144])
		); 

/******************* CELL 4145 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4145 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4049]),
			.N(gen[4050]),
			.NE(gen[4051]),

			.O(gen[4144]),
			.E(gen[4146]),

			.SO(gen[4239]),
			.S(gen[4240]),
			.SE(gen[4241]),

			.SELF(gen[4145]),
			.cell_state(gen[4145])
		); 

/******************* CELL 4146 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4146 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4050]),
			.N(gen[4051]),
			.NE(gen[4052]),

			.O(gen[4145]),
			.E(gen[4147]),

			.SO(gen[4240]),
			.S(gen[4241]),
			.SE(gen[4242]),

			.SELF(gen[4146]),
			.cell_state(gen[4146])
		); 

/******************* CELL 4147 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4147 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4051]),
			.N(gen[4052]),
			.NE(gen[4053]),

			.O(gen[4146]),
			.E(gen[4148]),

			.SO(gen[4241]),
			.S(gen[4242]),
			.SE(gen[4243]),

			.SELF(gen[4147]),
			.cell_state(gen[4147])
		); 

/******************* CELL 4148 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4148 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4052]),
			.N(gen[4053]),
			.NE(gen[4054]),

			.O(gen[4147]),
			.E(gen[4149]),

			.SO(gen[4242]),
			.S(gen[4243]),
			.SE(gen[4244]),

			.SELF(gen[4148]),
			.cell_state(gen[4148])
		); 

/******************* CELL 4149 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4149 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4053]),
			.N(gen[4054]),
			.NE(gen[4055]),

			.O(gen[4148]),
			.E(gen[4150]),

			.SO(gen[4243]),
			.S(gen[4244]),
			.SE(gen[4245]),

			.SELF(gen[4149]),
			.cell_state(gen[4149])
		); 

/******************* CELL 4150 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4150 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4054]),
			.N(gen[4055]),
			.NE(gen[4056]),

			.O(gen[4149]),
			.E(gen[4151]),

			.SO(gen[4244]),
			.S(gen[4245]),
			.SE(gen[4246]),

			.SELF(gen[4150]),
			.cell_state(gen[4150])
		); 

/******************* CELL 4151 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4151 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4055]),
			.N(gen[4056]),
			.NE(gen[4057]),

			.O(gen[4150]),
			.E(gen[4152]),

			.SO(gen[4245]),
			.S(gen[4246]),
			.SE(gen[4247]),

			.SELF(gen[4151]),
			.cell_state(gen[4151])
		); 

/******************* CELL 4152 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4152 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4056]),
			.N(gen[4057]),
			.NE(gen[4058]),

			.O(gen[4151]),
			.E(gen[4153]),

			.SO(gen[4246]),
			.S(gen[4247]),
			.SE(gen[4248]),

			.SELF(gen[4152]),
			.cell_state(gen[4152])
		); 

/******************* CELL 4153 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4153 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4057]),
			.N(gen[4058]),
			.NE(gen[4059]),

			.O(gen[4152]),
			.E(gen[4154]),

			.SO(gen[4247]),
			.S(gen[4248]),
			.SE(gen[4249]),

			.SELF(gen[4153]),
			.cell_state(gen[4153])
		); 

/******************* CELL 4154 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4154 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4058]),
			.N(gen[4059]),
			.NE(gen[4060]),

			.O(gen[4153]),
			.E(gen[4155]),

			.SO(gen[4248]),
			.S(gen[4249]),
			.SE(gen[4250]),

			.SELF(gen[4154]),
			.cell_state(gen[4154])
		); 

/******************* CELL 4155 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4155 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4059]),
			.N(gen[4060]),
			.NE(gen[4061]),

			.O(gen[4154]),
			.E(gen[4156]),

			.SO(gen[4249]),
			.S(gen[4250]),
			.SE(gen[4251]),

			.SELF(gen[4155]),
			.cell_state(gen[4155])
		); 

/******************* CELL 4156 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4156 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4060]),
			.N(gen[4061]),
			.NE(gen[4062]),

			.O(gen[4155]),
			.E(gen[4157]),

			.SO(gen[4250]),
			.S(gen[4251]),
			.SE(gen[4252]),

			.SELF(gen[4156]),
			.cell_state(gen[4156])
		); 

/******************* CELL 4157 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4157 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4061]),
			.N(gen[4062]),
			.NE(gen[4063]),

			.O(gen[4156]),
			.E(gen[4158]),

			.SO(gen[4251]),
			.S(gen[4252]),
			.SE(gen[4253]),

			.SELF(gen[4157]),
			.cell_state(gen[4157])
		); 

/******************* CELL 4158 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4158 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4062]),
			.N(gen[4063]),
			.NE(gen[4064]),

			.O(gen[4157]),
			.E(gen[4159]),

			.SO(gen[4252]),
			.S(gen[4253]),
			.SE(gen[4254]),

			.SELF(gen[4158]),
			.cell_state(gen[4158])
		); 

/******************* CELL 4159 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4159 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4063]),
			.N(gen[4064]),
			.NE(gen[4065]),

			.O(gen[4158]),
			.E(gen[4160]),

			.SO(gen[4253]),
			.S(gen[4254]),
			.SE(gen[4255]),

			.SELF(gen[4159]),
			.cell_state(gen[4159])
		); 

/******************* CELL 4160 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4160 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4064]),
			.N(gen[4065]),
			.NE(gen[4066]),

			.O(gen[4159]),
			.E(gen[4161]),

			.SO(gen[4254]),
			.S(gen[4255]),
			.SE(gen[4256]),

			.SELF(gen[4160]),
			.cell_state(gen[4160])
		); 

/******************* CELL 4161 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4161 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4065]),
			.N(gen[4066]),
			.NE(gen[4067]),

			.O(gen[4160]),
			.E(gen[4162]),

			.SO(gen[4255]),
			.S(gen[4256]),
			.SE(gen[4257]),

			.SELF(gen[4161]),
			.cell_state(gen[4161])
		); 

/******************* CELL 4162 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4162 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4066]),
			.N(gen[4067]),
			.NE(gen[4068]),

			.O(gen[4161]),
			.E(gen[4163]),

			.SO(gen[4256]),
			.S(gen[4257]),
			.SE(gen[4258]),

			.SELF(gen[4162]),
			.cell_state(gen[4162])
		); 

/******************* CELL 4163 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4163 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4067]),
			.N(gen[4068]),
			.NE(gen[4069]),

			.O(gen[4162]),
			.E(gen[4164]),

			.SO(gen[4257]),
			.S(gen[4258]),
			.SE(gen[4259]),

			.SELF(gen[4163]),
			.cell_state(gen[4163])
		); 

/******************* CELL 4164 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4164 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4068]),
			.N(gen[4069]),
			.NE(gen[4070]),

			.O(gen[4163]),
			.E(gen[4165]),

			.SO(gen[4258]),
			.S(gen[4259]),
			.SE(gen[4260]),

			.SELF(gen[4164]),
			.cell_state(gen[4164])
		); 

/******************* CELL 4165 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4165 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4069]),
			.N(gen[4070]),
			.NE(gen[4071]),

			.O(gen[4164]),
			.E(gen[4166]),

			.SO(gen[4259]),
			.S(gen[4260]),
			.SE(gen[4261]),

			.SELF(gen[4165]),
			.cell_state(gen[4165])
		); 

/******************* CELL 4166 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4166 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4070]),
			.N(gen[4071]),
			.NE(gen[4072]),

			.O(gen[4165]),
			.E(gen[4167]),

			.SO(gen[4260]),
			.S(gen[4261]),
			.SE(gen[4262]),

			.SELF(gen[4166]),
			.cell_state(gen[4166])
		); 

/******************* CELL 4167 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4167 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4071]),
			.N(gen[4072]),
			.NE(gen[4073]),

			.O(gen[4166]),
			.E(gen[4168]),

			.SO(gen[4261]),
			.S(gen[4262]),
			.SE(gen[4263]),

			.SELF(gen[4167]),
			.cell_state(gen[4167])
		); 

/******************* CELL 4168 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4168 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4072]),
			.N(gen[4073]),
			.NE(gen[4074]),

			.O(gen[4167]),
			.E(gen[4169]),

			.SO(gen[4262]),
			.S(gen[4263]),
			.SE(gen[4264]),

			.SELF(gen[4168]),
			.cell_state(gen[4168])
		); 

/******************* CELL 4169 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4169 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4073]),
			.N(gen[4074]),
			.NE(gen[4075]),

			.O(gen[4168]),
			.E(gen[4170]),

			.SO(gen[4263]),
			.S(gen[4264]),
			.SE(gen[4265]),

			.SELF(gen[4169]),
			.cell_state(gen[4169])
		); 

/******************* CELL 4170 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4170 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4074]),
			.N(gen[4075]),
			.NE(gen[4076]),

			.O(gen[4169]),
			.E(gen[4171]),

			.SO(gen[4264]),
			.S(gen[4265]),
			.SE(gen[4266]),

			.SELF(gen[4170]),
			.cell_state(gen[4170])
		); 

/******************* CELL 4171 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4171 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4075]),
			.N(gen[4076]),
			.NE(gen[4077]),

			.O(gen[4170]),
			.E(gen[4172]),

			.SO(gen[4265]),
			.S(gen[4266]),
			.SE(gen[4267]),

			.SELF(gen[4171]),
			.cell_state(gen[4171])
		); 

/******************* CELL 4172 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4172 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4076]),
			.N(gen[4077]),
			.NE(gen[4078]),

			.O(gen[4171]),
			.E(gen[4173]),

			.SO(gen[4266]),
			.S(gen[4267]),
			.SE(gen[4268]),

			.SELF(gen[4172]),
			.cell_state(gen[4172])
		); 

/******************* CELL 4173 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4173 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4077]),
			.N(gen[4078]),
			.NE(gen[4079]),

			.O(gen[4172]),
			.E(gen[4174]),

			.SO(gen[4267]),
			.S(gen[4268]),
			.SE(gen[4269]),

			.SELF(gen[4173]),
			.cell_state(gen[4173])
		); 

/******************* CELL 4174 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4174 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4078]),
			.N(gen[4079]),
			.NE(gen[4080]),

			.O(gen[4173]),
			.E(gen[4175]),

			.SO(gen[4268]),
			.S(gen[4269]),
			.SE(gen[4270]),

			.SELF(gen[4174]),
			.cell_state(gen[4174])
		); 

/******************* CELL 4175 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4175 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4079]),
			.N(gen[4080]),
			.NE(gen[4081]),

			.O(gen[4174]),
			.E(gen[4176]),

			.SO(gen[4269]),
			.S(gen[4270]),
			.SE(gen[4271]),

			.SELF(gen[4175]),
			.cell_state(gen[4175])
		); 

/******************* CELL 4176 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4176 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4080]),
			.N(gen[4081]),
			.NE(gen[4082]),

			.O(gen[4175]),
			.E(gen[4177]),

			.SO(gen[4270]),
			.S(gen[4271]),
			.SE(gen[4272]),

			.SELF(gen[4176]),
			.cell_state(gen[4176])
		); 

/******************* CELL 4177 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4177 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4081]),
			.N(gen[4082]),
			.NE(gen[4083]),

			.O(gen[4176]),
			.E(gen[4178]),

			.SO(gen[4271]),
			.S(gen[4272]),
			.SE(gen[4273]),

			.SELF(gen[4177]),
			.cell_state(gen[4177])
		); 

/******************* CELL 4178 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4178 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4082]),
			.N(gen[4083]),
			.NE(gen[4084]),

			.O(gen[4177]),
			.E(gen[4179]),

			.SO(gen[4272]),
			.S(gen[4273]),
			.SE(gen[4274]),

			.SELF(gen[4178]),
			.cell_state(gen[4178])
		); 

/******************* CELL 4179 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4179 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4083]),
			.N(gen[4084]),
			.NE(gen[4083]),

			.O(gen[4178]),
			.E(gen[4178]),

			.SO(gen[4273]),
			.S(gen[4274]),
			.SE(gen[4273]),

			.SELF(gen[4179]),
			.cell_state(gen[4179])
		); 

/******************* CELL 4180 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4180 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4086]),
			.N(gen[4085]),
			.NE(gen[4086]),

			.O(gen[4181]),
			.E(gen[4181]),

			.SO(gen[4276]),
			.S(gen[4275]),
			.SE(gen[4276]),

			.SELF(gen[4180]),
			.cell_state(gen[4180])
		); 

/******************* CELL 4181 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4181 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4085]),
			.N(gen[4086]),
			.NE(gen[4087]),

			.O(gen[4180]),
			.E(gen[4182]),

			.SO(gen[4275]),
			.S(gen[4276]),
			.SE(gen[4277]),

			.SELF(gen[4181]),
			.cell_state(gen[4181])
		); 

/******************* CELL 4182 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4182 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4086]),
			.N(gen[4087]),
			.NE(gen[4088]),

			.O(gen[4181]),
			.E(gen[4183]),

			.SO(gen[4276]),
			.S(gen[4277]),
			.SE(gen[4278]),

			.SELF(gen[4182]),
			.cell_state(gen[4182])
		); 

/******************* CELL 4183 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4183 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4087]),
			.N(gen[4088]),
			.NE(gen[4089]),

			.O(gen[4182]),
			.E(gen[4184]),

			.SO(gen[4277]),
			.S(gen[4278]),
			.SE(gen[4279]),

			.SELF(gen[4183]),
			.cell_state(gen[4183])
		); 

/******************* CELL 4184 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4184 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4088]),
			.N(gen[4089]),
			.NE(gen[4090]),

			.O(gen[4183]),
			.E(gen[4185]),

			.SO(gen[4278]),
			.S(gen[4279]),
			.SE(gen[4280]),

			.SELF(gen[4184]),
			.cell_state(gen[4184])
		); 

/******************* CELL 4185 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4185 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4089]),
			.N(gen[4090]),
			.NE(gen[4091]),

			.O(gen[4184]),
			.E(gen[4186]),

			.SO(gen[4279]),
			.S(gen[4280]),
			.SE(gen[4281]),

			.SELF(gen[4185]),
			.cell_state(gen[4185])
		); 

/******************* CELL 4186 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4186 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4090]),
			.N(gen[4091]),
			.NE(gen[4092]),

			.O(gen[4185]),
			.E(gen[4187]),

			.SO(gen[4280]),
			.S(gen[4281]),
			.SE(gen[4282]),

			.SELF(gen[4186]),
			.cell_state(gen[4186])
		); 

/******************* CELL 4187 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4187 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4091]),
			.N(gen[4092]),
			.NE(gen[4093]),

			.O(gen[4186]),
			.E(gen[4188]),

			.SO(gen[4281]),
			.S(gen[4282]),
			.SE(gen[4283]),

			.SELF(gen[4187]),
			.cell_state(gen[4187])
		); 

/******************* CELL 4188 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4188 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4092]),
			.N(gen[4093]),
			.NE(gen[4094]),

			.O(gen[4187]),
			.E(gen[4189]),

			.SO(gen[4282]),
			.S(gen[4283]),
			.SE(gen[4284]),

			.SELF(gen[4188]),
			.cell_state(gen[4188])
		); 

/******************* CELL 4189 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4189 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4093]),
			.N(gen[4094]),
			.NE(gen[4095]),

			.O(gen[4188]),
			.E(gen[4190]),

			.SO(gen[4283]),
			.S(gen[4284]),
			.SE(gen[4285]),

			.SELF(gen[4189]),
			.cell_state(gen[4189])
		); 

/******************* CELL 4190 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4190 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4094]),
			.N(gen[4095]),
			.NE(gen[4096]),

			.O(gen[4189]),
			.E(gen[4191]),

			.SO(gen[4284]),
			.S(gen[4285]),
			.SE(gen[4286]),

			.SELF(gen[4190]),
			.cell_state(gen[4190])
		); 

/******************* CELL 4191 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4191 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4095]),
			.N(gen[4096]),
			.NE(gen[4097]),

			.O(gen[4190]),
			.E(gen[4192]),

			.SO(gen[4285]),
			.S(gen[4286]),
			.SE(gen[4287]),

			.SELF(gen[4191]),
			.cell_state(gen[4191])
		); 

/******************* CELL 4192 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4192 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4096]),
			.N(gen[4097]),
			.NE(gen[4098]),

			.O(gen[4191]),
			.E(gen[4193]),

			.SO(gen[4286]),
			.S(gen[4287]),
			.SE(gen[4288]),

			.SELF(gen[4192]),
			.cell_state(gen[4192])
		); 

/******************* CELL 4193 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4193 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4097]),
			.N(gen[4098]),
			.NE(gen[4099]),

			.O(gen[4192]),
			.E(gen[4194]),

			.SO(gen[4287]),
			.S(gen[4288]),
			.SE(gen[4289]),

			.SELF(gen[4193]),
			.cell_state(gen[4193])
		); 

/******************* CELL 4194 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4194 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4098]),
			.N(gen[4099]),
			.NE(gen[4100]),

			.O(gen[4193]),
			.E(gen[4195]),

			.SO(gen[4288]),
			.S(gen[4289]),
			.SE(gen[4290]),

			.SELF(gen[4194]),
			.cell_state(gen[4194])
		); 

/******************* CELL 4195 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4195 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4099]),
			.N(gen[4100]),
			.NE(gen[4101]),

			.O(gen[4194]),
			.E(gen[4196]),

			.SO(gen[4289]),
			.S(gen[4290]),
			.SE(gen[4291]),

			.SELF(gen[4195]),
			.cell_state(gen[4195])
		); 

/******************* CELL 4196 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4196 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4100]),
			.N(gen[4101]),
			.NE(gen[4102]),

			.O(gen[4195]),
			.E(gen[4197]),

			.SO(gen[4290]),
			.S(gen[4291]),
			.SE(gen[4292]),

			.SELF(gen[4196]),
			.cell_state(gen[4196])
		); 

/******************* CELL 4197 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4197 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4101]),
			.N(gen[4102]),
			.NE(gen[4103]),

			.O(gen[4196]),
			.E(gen[4198]),

			.SO(gen[4291]),
			.S(gen[4292]),
			.SE(gen[4293]),

			.SELF(gen[4197]),
			.cell_state(gen[4197])
		); 

/******************* CELL 4198 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4198 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4102]),
			.N(gen[4103]),
			.NE(gen[4104]),

			.O(gen[4197]),
			.E(gen[4199]),

			.SO(gen[4292]),
			.S(gen[4293]),
			.SE(gen[4294]),

			.SELF(gen[4198]),
			.cell_state(gen[4198])
		); 

/******************* CELL 4199 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4199 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4103]),
			.N(gen[4104]),
			.NE(gen[4105]),

			.O(gen[4198]),
			.E(gen[4200]),

			.SO(gen[4293]),
			.S(gen[4294]),
			.SE(gen[4295]),

			.SELF(gen[4199]),
			.cell_state(gen[4199])
		); 

/******************* CELL 4200 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4200 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4104]),
			.N(gen[4105]),
			.NE(gen[4106]),

			.O(gen[4199]),
			.E(gen[4201]),

			.SO(gen[4294]),
			.S(gen[4295]),
			.SE(gen[4296]),

			.SELF(gen[4200]),
			.cell_state(gen[4200])
		); 

/******************* CELL 4201 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4201 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4105]),
			.N(gen[4106]),
			.NE(gen[4107]),

			.O(gen[4200]),
			.E(gen[4202]),

			.SO(gen[4295]),
			.S(gen[4296]),
			.SE(gen[4297]),

			.SELF(gen[4201]),
			.cell_state(gen[4201])
		); 

/******************* CELL 4202 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4202 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4106]),
			.N(gen[4107]),
			.NE(gen[4108]),

			.O(gen[4201]),
			.E(gen[4203]),

			.SO(gen[4296]),
			.S(gen[4297]),
			.SE(gen[4298]),

			.SELF(gen[4202]),
			.cell_state(gen[4202])
		); 

/******************* CELL 4203 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4203 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4107]),
			.N(gen[4108]),
			.NE(gen[4109]),

			.O(gen[4202]),
			.E(gen[4204]),

			.SO(gen[4297]),
			.S(gen[4298]),
			.SE(gen[4299]),

			.SELF(gen[4203]),
			.cell_state(gen[4203])
		); 

/******************* CELL 4204 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4204 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4108]),
			.N(gen[4109]),
			.NE(gen[4110]),

			.O(gen[4203]),
			.E(gen[4205]),

			.SO(gen[4298]),
			.S(gen[4299]),
			.SE(gen[4300]),

			.SELF(gen[4204]),
			.cell_state(gen[4204])
		); 

/******************* CELL 4205 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4205 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4109]),
			.N(gen[4110]),
			.NE(gen[4111]),

			.O(gen[4204]),
			.E(gen[4206]),

			.SO(gen[4299]),
			.S(gen[4300]),
			.SE(gen[4301]),

			.SELF(gen[4205]),
			.cell_state(gen[4205])
		); 

/******************* CELL 4206 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4206 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4110]),
			.N(gen[4111]),
			.NE(gen[4112]),

			.O(gen[4205]),
			.E(gen[4207]),

			.SO(gen[4300]),
			.S(gen[4301]),
			.SE(gen[4302]),

			.SELF(gen[4206]),
			.cell_state(gen[4206])
		); 

/******************* CELL 4207 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4207 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4111]),
			.N(gen[4112]),
			.NE(gen[4113]),

			.O(gen[4206]),
			.E(gen[4208]),

			.SO(gen[4301]),
			.S(gen[4302]),
			.SE(gen[4303]),

			.SELF(gen[4207]),
			.cell_state(gen[4207])
		); 

/******************* CELL 4208 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4208 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4112]),
			.N(gen[4113]),
			.NE(gen[4114]),

			.O(gen[4207]),
			.E(gen[4209]),

			.SO(gen[4302]),
			.S(gen[4303]),
			.SE(gen[4304]),

			.SELF(gen[4208]),
			.cell_state(gen[4208])
		); 

/******************* CELL 4209 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4209 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4113]),
			.N(gen[4114]),
			.NE(gen[4115]),

			.O(gen[4208]),
			.E(gen[4210]),

			.SO(gen[4303]),
			.S(gen[4304]),
			.SE(gen[4305]),

			.SELF(gen[4209]),
			.cell_state(gen[4209])
		); 

/******************* CELL 4210 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4210 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4114]),
			.N(gen[4115]),
			.NE(gen[4116]),

			.O(gen[4209]),
			.E(gen[4211]),

			.SO(gen[4304]),
			.S(gen[4305]),
			.SE(gen[4306]),

			.SELF(gen[4210]),
			.cell_state(gen[4210])
		); 

/******************* CELL 4211 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4211 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4115]),
			.N(gen[4116]),
			.NE(gen[4117]),

			.O(gen[4210]),
			.E(gen[4212]),

			.SO(gen[4305]),
			.S(gen[4306]),
			.SE(gen[4307]),

			.SELF(gen[4211]),
			.cell_state(gen[4211])
		); 

/******************* CELL 4212 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4212 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4116]),
			.N(gen[4117]),
			.NE(gen[4118]),

			.O(gen[4211]),
			.E(gen[4213]),

			.SO(gen[4306]),
			.S(gen[4307]),
			.SE(gen[4308]),

			.SELF(gen[4212]),
			.cell_state(gen[4212])
		); 

/******************* CELL 4213 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4213 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4117]),
			.N(gen[4118]),
			.NE(gen[4119]),

			.O(gen[4212]),
			.E(gen[4214]),

			.SO(gen[4307]),
			.S(gen[4308]),
			.SE(gen[4309]),

			.SELF(gen[4213]),
			.cell_state(gen[4213])
		); 

/******************* CELL 4214 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4214 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4118]),
			.N(gen[4119]),
			.NE(gen[4120]),

			.O(gen[4213]),
			.E(gen[4215]),

			.SO(gen[4308]),
			.S(gen[4309]),
			.SE(gen[4310]),

			.SELF(gen[4214]),
			.cell_state(gen[4214])
		); 

/******************* CELL 4215 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4215 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4119]),
			.N(gen[4120]),
			.NE(gen[4121]),

			.O(gen[4214]),
			.E(gen[4216]),

			.SO(gen[4309]),
			.S(gen[4310]),
			.SE(gen[4311]),

			.SELF(gen[4215]),
			.cell_state(gen[4215])
		); 

/******************* CELL 4216 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4216 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4120]),
			.N(gen[4121]),
			.NE(gen[4122]),

			.O(gen[4215]),
			.E(gen[4217]),

			.SO(gen[4310]),
			.S(gen[4311]),
			.SE(gen[4312]),

			.SELF(gen[4216]),
			.cell_state(gen[4216])
		); 

/******************* CELL 4217 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4217 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4121]),
			.N(gen[4122]),
			.NE(gen[4123]),

			.O(gen[4216]),
			.E(gen[4218]),

			.SO(gen[4311]),
			.S(gen[4312]),
			.SE(gen[4313]),

			.SELF(gen[4217]),
			.cell_state(gen[4217])
		); 

/******************* CELL 4218 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4218 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4122]),
			.N(gen[4123]),
			.NE(gen[4124]),

			.O(gen[4217]),
			.E(gen[4219]),

			.SO(gen[4312]),
			.S(gen[4313]),
			.SE(gen[4314]),

			.SELF(gen[4218]),
			.cell_state(gen[4218])
		); 

/******************* CELL 4219 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4219 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4123]),
			.N(gen[4124]),
			.NE(gen[4125]),

			.O(gen[4218]),
			.E(gen[4220]),

			.SO(gen[4313]),
			.S(gen[4314]),
			.SE(gen[4315]),

			.SELF(gen[4219]),
			.cell_state(gen[4219])
		); 

/******************* CELL 4220 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4220 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4124]),
			.N(gen[4125]),
			.NE(gen[4126]),

			.O(gen[4219]),
			.E(gen[4221]),

			.SO(gen[4314]),
			.S(gen[4315]),
			.SE(gen[4316]),

			.SELF(gen[4220]),
			.cell_state(gen[4220])
		); 

/******************* CELL 4221 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4221 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4125]),
			.N(gen[4126]),
			.NE(gen[4127]),

			.O(gen[4220]),
			.E(gen[4222]),

			.SO(gen[4315]),
			.S(gen[4316]),
			.SE(gen[4317]),

			.SELF(gen[4221]),
			.cell_state(gen[4221])
		); 

/******************* CELL 4222 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4222 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4126]),
			.N(gen[4127]),
			.NE(gen[4128]),

			.O(gen[4221]),
			.E(gen[4223]),

			.SO(gen[4316]),
			.S(gen[4317]),
			.SE(gen[4318]),

			.SELF(gen[4222]),
			.cell_state(gen[4222])
		); 

/******************* CELL 4223 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4223 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4127]),
			.N(gen[4128]),
			.NE(gen[4129]),

			.O(gen[4222]),
			.E(gen[4224]),

			.SO(gen[4317]),
			.S(gen[4318]),
			.SE(gen[4319]),

			.SELF(gen[4223]),
			.cell_state(gen[4223])
		); 

/******************* CELL 4224 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4224 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4128]),
			.N(gen[4129]),
			.NE(gen[4130]),

			.O(gen[4223]),
			.E(gen[4225]),

			.SO(gen[4318]),
			.S(gen[4319]),
			.SE(gen[4320]),

			.SELF(gen[4224]),
			.cell_state(gen[4224])
		); 

/******************* CELL 4225 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4225 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4129]),
			.N(gen[4130]),
			.NE(gen[4131]),

			.O(gen[4224]),
			.E(gen[4226]),

			.SO(gen[4319]),
			.S(gen[4320]),
			.SE(gen[4321]),

			.SELF(gen[4225]),
			.cell_state(gen[4225])
		); 

/******************* CELL 4226 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4226 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4130]),
			.N(gen[4131]),
			.NE(gen[4132]),

			.O(gen[4225]),
			.E(gen[4227]),

			.SO(gen[4320]),
			.S(gen[4321]),
			.SE(gen[4322]),

			.SELF(gen[4226]),
			.cell_state(gen[4226])
		); 

/******************* CELL 4227 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4227 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4131]),
			.N(gen[4132]),
			.NE(gen[4133]),

			.O(gen[4226]),
			.E(gen[4228]),

			.SO(gen[4321]),
			.S(gen[4322]),
			.SE(gen[4323]),

			.SELF(gen[4227]),
			.cell_state(gen[4227])
		); 

/******************* CELL 4228 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4228 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4132]),
			.N(gen[4133]),
			.NE(gen[4134]),

			.O(gen[4227]),
			.E(gen[4229]),

			.SO(gen[4322]),
			.S(gen[4323]),
			.SE(gen[4324]),

			.SELF(gen[4228]),
			.cell_state(gen[4228])
		); 

/******************* CELL 4229 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4229 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4133]),
			.N(gen[4134]),
			.NE(gen[4135]),

			.O(gen[4228]),
			.E(gen[4230]),

			.SO(gen[4323]),
			.S(gen[4324]),
			.SE(gen[4325]),

			.SELF(gen[4229]),
			.cell_state(gen[4229])
		); 

/******************* CELL 4230 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4230 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4134]),
			.N(gen[4135]),
			.NE(gen[4136]),

			.O(gen[4229]),
			.E(gen[4231]),

			.SO(gen[4324]),
			.S(gen[4325]),
			.SE(gen[4326]),

			.SELF(gen[4230]),
			.cell_state(gen[4230])
		); 

/******************* CELL 4231 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4231 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4135]),
			.N(gen[4136]),
			.NE(gen[4137]),

			.O(gen[4230]),
			.E(gen[4232]),

			.SO(gen[4325]),
			.S(gen[4326]),
			.SE(gen[4327]),

			.SELF(gen[4231]),
			.cell_state(gen[4231])
		); 

/******************* CELL 4232 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4232 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4136]),
			.N(gen[4137]),
			.NE(gen[4138]),

			.O(gen[4231]),
			.E(gen[4233]),

			.SO(gen[4326]),
			.S(gen[4327]),
			.SE(gen[4328]),

			.SELF(gen[4232]),
			.cell_state(gen[4232])
		); 

/******************* CELL 4233 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4233 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4137]),
			.N(gen[4138]),
			.NE(gen[4139]),

			.O(gen[4232]),
			.E(gen[4234]),

			.SO(gen[4327]),
			.S(gen[4328]),
			.SE(gen[4329]),

			.SELF(gen[4233]),
			.cell_state(gen[4233])
		); 

/******************* CELL 4234 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4234 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4138]),
			.N(gen[4139]),
			.NE(gen[4140]),

			.O(gen[4233]),
			.E(gen[4235]),

			.SO(gen[4328]),
			.S(gen[4329]),
			.SE(gen[4330]),

			.SELF(gen[4234]),
			.cell_state(gen[4234])
		); 

/******************* CELL 4235 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4235 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4139]),
			.N(gen[4140]),
			.NE(gen[4141]),

			.O(gen[4234]),
			.E(gen[4236]),

			.SO(gen[4329]),
			.S(gen[4330]),
			.SE(gen[4331]),

			.SELF(gen[4235]),
			.cell_state(gen[4235])
		); 

/******************* CELL 4236 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4236 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4140]),
			.N(gen[4141]),
			.NE(gen[4142]),

			.O(gen[4235]),
			.E(gen[4237]),

			.SO(gen[4330]),
			.S(gen[4331]),
			.SE(gen[4332]),

			.SELF(gen[4236]),
			.cell_state(gen[4236])
		); 

/******************* CELL 4237 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4237 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4141]),
			.N(gen[4142]),
			.NE(gen[4143]),

			.O(gen[4236]),
			.E(gen[4238]),

			.SO(gen[4331]),
			.S(gen[4332]),
			.SE(gen[4333]),

			.SELF(gen[4237]),
			.cell_state(gen[4237])
		); 

/******************* CELL 4238 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4238 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4142]),
			.N(gen[4143]),
			.NE(gen[4144]),

			.O(gen[4237]),
			.E(gen[4239]),

			.SO(gen[4332]),
			.S(gen[4333]),
			.SE(gen[4334]),

			.SELF(gen[4238]),
			.cell_state(gen[4238])
		); 

/******************* CELL 4239 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4239 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4143]),
			.N(gen[4144]),
			.NE(gen[4145]),

			.O(gen[4238]),
			.E(gen[4240]),

			.SO(gen[4333]),
			.S(gen[4334]),
			.SE(gen[4335]),

			.SELF(gen[4239]),
			.cell_state(gen[4239])
		); 

/******************* CELL 4240 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4240 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4144]),
			.N(gen[4145]),
			.NE(gen[4146]),

			.O(gen[4239]),
			.E(gen[4241]),

			.SO(gen[4334]),
			.S(gen[4335]),
			.SE(gen[4336]),

			.SELF(gen[4240]),
			.cell_state(gen[4240])
		); 

/******************* CELL 4241 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4241 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4145]),
			.N(gen[4146]),
			.NE(gen[4147]),

			.O(gen[4240]),
			.E(gen[4242]),

			.SO(gen[4335]),
			.S(gen[4336]),
			.SE(gen[4337]),

			.SELF(gen[4241]),
			.cell_state(gen[4241])
		); 

/******************* CELL 4242 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4242 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4146]),
			.N(gen[4147]),
			.NE(gen[4148]),

			.O(gen[4241]),
			.E(gen[4243]),

			.SO(gen[4336]),
			.S(gen[4337]),
			.SE(gen[4338]),

			.SELF(gen[4242]),
			.cell_state(gen[4242])
		); 

/******************* CELL 4243 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4243 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4147]),
			.N(gen[4148]),
			.NE(gen[4149]),

			.O(gen[4242]),
			.E(gen[4244]),

			.SO(gen[4337]),
			.S(gen[4338]),
			.SE(gen[4339]),

			.SELF(gen[4243]),
			.cell_state(gen[4243])
		); 

/******************* CELL 4244 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4244 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4148]),
			.N(gen[4149]),
			.NE(gen[4150]),

			.O(gen[4243]),
			.E(gen[4245]),

			.SO(gen[4338]),
			.S(gen[4339]),
			.SE(gen[4340]),

			.SELF(gen[4244]),
			.cell_state(gen[4244])
		); 

/******************* CELL 4245 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4245 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4149]),
			.N(gen[4150]),
			.NE(gen[4151]),

			.O(gen[4244]),
			.E(gen[4246]),

			.SO(gen[4339]),
			.S(gen[4340]),
			.SE(gen[4341]),

			.SELF(gen[4245]),
			.cell_state(gen[4245])
		); 

/******************* CELL 4246 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4246 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4150]),
			.N(gen[4151]),
			.NE(gen[4152]),

			.O(gen[4245]),
			.E(gen[4247]),

			.SO(gen[4340]),
			.S(gen[4341]),
			.SE(gen[4342]),

			.SELF(gen[4246]),
			.cell_state(gen[4246])
		); 

/******************* CELL 4247 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4247 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4151]),
			.N(gen[4152]),
			.NE(gen[4153]),

			.O(gen[4246]),
			.E(gen[4248]),

			.SO(gen[4341]),
			.S(gen[4342]),
			.SE(gen[4343]),

			.SELF(gen[4247]),
			.cell_state(gen[4247])
		); 

/******************* CELL 4248 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4248 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4152]),
			.N(gen[4153]),
			.NE(gen[4154]),

			.O(gen[4247]),
			.E(gen[4249]),

			.SO(gen[4342]),
			.S(gen[4343]),
			.SE(gen[4344]),

			.SELF(gen[4248]),
			.cell_state(gen[4248])
		); 

/******************* CELL 4249 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4249 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4153]),
			.N(gen[4154]),
			.NE(gen[4155]),

			.O(gen[4248]),
			.E(gen[4250]),

			.SO(gen[4343]),
			.S(gen[4344]),
			.SE(gen[4345]),

			.SELF(gen[4249]),
			.cell_state(gen[4249])
		); 

/******************* CELL 4250 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4250 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4154]),
			.N(gen[4155]),
			.NE(gen[4156]),

			.O(gen[4249]),
			.E(gen[4251]),

			.SO(gen[4344]),
			.S(gen[4345]),
			.SE(gen[4346]),

			.SELF(gen[4250]),
			.cell_state(gen[4250])
		); 

/******************* CELL 4251 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4251 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4155]),
			.N(gen[4156]),
			.NE(gen[4157]),

			.O(gen[4250]),
			.E(gen[4252]),

			.SO(gen[4345]),
			.S(gen[4346]),
			.SE(gen[4347]),

			.SELF(gen[4251]),
			.cell_state(gen[4251])
		); 

/******************* CELL 4252 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4252 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4156]),
			.N(gen[4157]),
			.NE(gen[4158]),

			.O(gen[4251]),
			.E(gen[4253]),

			.SO(gen[4346]),
			.S(gen[4347]),
			.SE(gen[4348]),

			.SELF(gen[4252]),
			.cell_state(gen[4252])
		); 

/******************* CELL 4253 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4253 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4157]),
			.N(gen[4158]),
			.NE(gen[4159]),

			.O(gen[4252]),
			.E(gen[4254]),

			.SO(gen[4347]),
			.S(gen[4348]),
			.SE(gen[4349]),

			.SELF(gen[4253]),
			.cell_state(gen[4253])
		); 

/******************* CELL 4254 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4254 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4158]),
			.N(gen[4159]),
			.NE(gen[4160]),

			.O(gen[4253]),
			.E(gen[4255]),

			.SO(gen[4348]),
			.S(gen[4349]),
			.SE(gen[4350]),

			.SELF(gen[4254]),
			.cell_state(gen[4254])
		); 

/******************* CELL 4255 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4255 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4159]),
			.N(gen[4160]),
			.NE(gen[4161]),

			.O(gen[4254]),
			.E(gen[4256]),

			.SO(gen[4349]),
			.S(gen[4350]),
			.SE(gen[4351]),

			.SELF(gen[4255]),
			.cell_state(gen[4255])
		); 

/******************* CELL 4256 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4256 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4160]),
			.N(gen[4161]),
			.NE(gen[4162]),

			.O(gen[4255]),
			.E(gen[4257]),

			.SO(gen[4350]),
			.S(gen[4351]),
			.SE(gen[4352]),

			.SELF(gen[4256]),
			.cell_state(gen[4256])
		); 

/******************* CELL 4257 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4257 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4161]),
			.N(gen[4162]),
			.NE(gen[4163]),

			.O(gen[4256]),
			.E(gen[4258]),

			.SO(gen[4351]),
			.S(gen[4352]),
			.SE(gen[4353]),

			.SELF(gen[4257]),
			.cell_state(gen[4257])
		); 

/******************* CELL 4258 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4258 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4162]),
			.N(gen[4163]),
			.NE(gen[4164]),

			.O(gen[4257]),
			.E(gen[4259]),

			.SO(gen[4352]),
			.S(gen[4353]),
			.SE(gen[4354]),

			.SELF(gen[4258]),
			.cell_state(gen[4258])
		); 

/******************* CELL 4259 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4259 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4163]),
			.N(gen[4164]),
			.NE(gen[4165]),

			.O(gen[4258]),
			.E(gen[4260]),

			.SO(gen[4353]),
			.S(gen[4354]),
			.SE(gen[4355]),

			.SELF(gen[4259]),
			.cell_state(gen[4259])
		); 

/******************* CELL 4260 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4260 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4164]),
			.N(gen[4165]),
			.NE(gen[4166]),

			.O(gen[4259]),
			.E(gen[4261]),

			.SO(gen[4354]),
			.S(gen[4355]),
			.SE(gen[4356]),

			.SELF(gen[4260]),
			.cell_state(gen[4260])
		); 

/******************* CELL 4261 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4261 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4165]),
			.N(gen[4166]),
			.NE(gen[4167]),

			.O(gen[4260]),
			.E(gen[4262]),

			.SO(gen[4355]),
			.S(gen[4356]),
			.SE(gen[4357]),

			.SELF(gen[4261]),
			.cell_state(gen[4261])
		); 

/******************* CELL 4262 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4262 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4166]),
			.N(gen[4167]),
			.NE(gen[4168]),

			.O(gen[4261]),
			.E(gen[4263]),

			.SO(gen[4356]),
			.S(gen[4357]),
			.SE(gen[4358]),

			.SELF(gen[4262]),
			.cell_state(gen[4262])
		); 

/******************* CELL 4263 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4263 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4167]),
			.N(gen[4168]),
			.NE(gen[4169]),

			.O(gen[4262]),
			.E(gen[4264]),

			.SO(gen[4357]),
			.S(gen[4358]),
			.SE(gen[4359]),

			.SELF(gen[4263]),
			.cell_state(gen[4263])
		); 

/******************* CELL 4264 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4264 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4168]),
			.N(gen[4169]),
			.NE(gen[4170]),

			.O(gen[4263]),
			.E(gen[4265]),

			.SO(gen[4358]),
			.S(gen[4359]),
			.SE(gen[4360]),

			.SELF(gen[4264]),
			.cell_state(gen[4264])
		); 

/******************* CELL 4265 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4265 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4169]),
			.N(gen[4170]),
			.NE(gen[4171]),

			.O(gen[4264]),
			.E(gen[4266]),

			.SO(gen[4359]),
			.S(gen[4360]),
			.SE(gen[4361]),

			.SELF(gen[4265]),
			.cell_state(gen[4265])
		); 

/******************* CELL 4266 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4266 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4170]),
			.N(gen[4171]),
			.NE(gen[4172]),

			.O(gen[4265]),
			.E(gen[4267]),

			.SO(gen[4360]),
			.S(gen[4361]),
			.SE(gen[4362]),

			.SELF(gen[4266]),
			.cell_state(gen[4266])
		); 

/******************* CELL 4267 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4267 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4171]),
			.N(gen[4172]),
			.NE(gen[4173]),

			.O(gen[4266]),
			.E(gen[4268]),

			.SO(gen[4361]),
			.S(gen[4362]),
			.SE(gen[4363]),

			.SELF(gen[4267]),
			.cell_state(gen[4267])
		); 

/******************* CELL 4268 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4268 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4172]),
			.N(gen[4173]),
			.NE(gen[4174]),

			.O(gen[4267]),
			.E(gen[4269]),

			.SO(gen[4362]),
			.S(gen[4363]),
			.SE(gen[4364]),

			.SELF(gen[4268]),
			.cell_state(gen[4268])
		); 

/******************* CELL 4269 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4269 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4173]),
			.N(gen[4174]),
			.NE(gen[4175]),

			.O(gen[4268]),
			.E(gen[4270]),

			.SO(gen[4363]),
			.S(gen[4364]),
			.SE(gen[4365]),

			.SELF(gen[4269]),
			.cell_state(gen[4269])
		); 

/******************* CELL 4270 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4270 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4174]),
			.N(gen[4175]),
			.NE(gen[4176]),

			.O(gen[4269]),
			.E(gen[4271]),

			.SO(gen[4364]),
			.S(gen[4365]),
			.SE(gen[4366]),

			.SELF(gen[4270]),
			.cell_state(gen[4270])
		); 

/******************* CELL 4271 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4271 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4175]),
			.N(gen[4176]),
			.NE(gen[4177]),

			.O(gen[4270]),
			.E(gen[4272]),

			.SO(gen[4365]),
			.S(gen[4366]),
			.SE(gen[4367]),

			.SELF(gen[4271]),
			.cell_state(gen[4271])
		); 

/******************* CELL 4272 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4272 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4176]),
			.N(gen[4177]),
			.NE(gen[4178]),

			.O(gen[4271]),
			.E(gen[4273]),

			.SO(gen[4366]),
			.S(gen[4367]),
			.SE(gen[4368]),

			.SELF(gen[4272]),
			.cell_state(gen[4272])
		); 

/******************* CELL 4273 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4273 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4177]),
			.N(gen[4178]),
			.NE(gen[4179]),

			.O(gen[4272]),
			.E(gen[4274]),

			.SO(gen[4367]),
			.S(gen[4368]),
			.SE(gen[4369]),

			.SELF(gen[4273]),
			.cell_state(gen[4273])
		); 

/******************* CELL 4274 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4274 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4178]),
			.N(gen[4179]),
			.NE(gen[4178]),

			.O(gen[4273]),
			.E(gen[4273]),

			.SO(gen[4368]),
			.S(gen[4369]),
			.SE(gen[4368]),

			.SELF(gen[4274]),
			.cell_state(gen[4274])
		); 

/******************* CELL 4275 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4275 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4181]),
			.N(gen[4180]),
			.NE(gen[4181]),

			.O(gen[4276]),
			.E(gen[4276]),

			.SO(gen[4371]),
			.S(gen[4370]),
			.SE(gen[4371]),

			.SELF(gen[4275]),
			.cell_state(gen[4275])
		); 

/******************* CELL 4276 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4276 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4180]),
			.N(gen[4181]),
			.NE(gen[4182]),

			.O(gen[4275]),
			.E(gen[4277]),

			.SO(gen[4370]),
			.S(gen[4371]),
			.SE(gen[4372]),

			.SELF(gen[4276]),
			.cell_state(gen[4276])
		); 

/******************* CELL 4277 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4277 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4181]),
			.N(gen[4182]),
			.NE(gen[4183]),

			.O(gen[4276]),
			.E(gen[4278]),

			.SO(gen[4371]),
			.S(gen[4372]),
			.SE(gen[4373]),

			.SELF(gen[4277]),
			.cell_state(gen[4277])
		); 

/******************* CELL 4278 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4278 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4182]),
			.N(gen[4183]),
			.NE(gen[4184]),

			.O(gen[4277]),
			.E(gen[4279]),

			.SO(gen[4372]),
			.S(gen[4373]),
			.SE(gen[4374]),

			.SELF(gen[4278]),
			.cell_state(gen[4278])
		); 

/******************* CELL 4279 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4279 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4183]),
			.N(gen[4184]),
			.NE(gen[4185]),

			.O(gen[4278]),
			.E(gen[4280]),

			.SO(gen[4373]),
			.S(gen[4374]),
			.SE(gen[4375]),

			.SELF(gen[4279]),
			.cell_state(gen[4279])
		); 

/******************* CELL 4280 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4280 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4184]),
			.N(gen[4185]),
			.NE(gen[4186]),

			.O(gen[4279]),
			.E(gen[4281]),

			.SO(gen[4374]),
			.S(gen[4375]),
			.SE(gen[4376]),

			.SELF(gen[4280]),
			.cell_state(gen[4280])
		); 

/******************* CELL 4281 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4281 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4185]),
			.N(gen[4186]),
			.NE(gen[4187]),

			.O(gen[4280]),
			.E(gen[4282]),

			.SO(gen[4375]),
			.S(gen[4376]),
			.SE(gen[4377]),

			.SELF(gen[4281]),
			.cell_state(gen[4281])
		); 

/******************* CELL 4282 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4282 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4186]),
			.N(gen[4187]),
			.NE(gen[4188]),

			.O(gen[4281]),
			.E(gen[4283]),

			.SO(gen[4376]),
			.S(gen[4377]),
			.SE(gen[4378]),

			.SELF(gen[4282]),
			.cell_state(gen[4282])
		); 

/******************* CELL 4283 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4283 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4187]),
			.N(gen[4188]),
			.NE(gen[4189]),

			.O(gen[4282]),
			.E(gen[4284]),

			.SO(gen[4377]),
			.S(gen[4378]),
			.SE(gen[4379]),

			.SELF(gen[4283]),
			.cell_state(gen[4283])
		); 

/******************* CELL 4284 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4284 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4188]),
			.N(gen[4189]),
			.NE(gen[4190]),

			.O(gen[4283]),
			.E(gen[4285]),

			.SO(gen[4378]),
			.S(gen[4379]),
			.SE(gen[4380]),

			.SELF(gen[4284]),
			.cell_state(gen[4284])
		); 

/******************* CELL 4285 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4285 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4189]),
			.N(gen[4190]),
			.NE(gen[4191]),

			.O(gen[4284]),
			.E(gen[4286]),

			.SO(gen[4379]),
			.S(gen[4380]),
			.SE(gen[4381]),

			.SELF(gen[4285]),
			.cell_state(gen[4285])
		); 

/******************* CELL 4286 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4286 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4190]),
			.N(gen[4191]),
			.NE(gen[4192]),

			.O(gen[4285]),
			.E(gen[4287]),

			.SO(gen[4380]),
			.S(gen[4381]),
			.SE(gen[4382]),

			.SELF(gen[4286]),
			.cell_state(gen[4286])
		); 

/******************* CELL 4287 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4287 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4191]),
			.N(gen[4192]),
			.NE(gen[4193]),

			.O(gen[4286]),
			.E(gen[4288]),

			.SO(gen[4381]),
			.S(gen[4382]),
			.SE(gen[4383]),

			.SELF(gen[4287]),
			.cell_state(gen[4287])
		); 

/******************* CELL 4288 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4288 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4192]),
			.N(gen[4193]),
			.NE(gen[4194]),

			.O(gen[4287]),
			.E(gen[4289]),

			.SO(gen[4382]),
			.S(gen[4383]),
			.SE(gen[4384]),

			.SELF(gen[4288]),
			.cell_state(gen[4288])
		); 

/******************* CELL 4289 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4289 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4193]),
			.N(gen[4194]),
			.NE(gen[4195]),

			.O(gen[4288]),
			.E(gen[4290]),

			.SO(gen[4383]),
			.S(gen[4384]),
			.SE(gen[4385]),

			.SELF(gen[4289]),
			.cell_state(gen[4289])
		); 

/******************* CELL 4290 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4290 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4194]),
			.N(gen[4195]),
			.NE(gen[4196]),

			.O(gen[4289]),
			.E(gen[4291]),

			.SO(gen[4384]),
			.S(gen[4385]),
			.SE(gen[4386]),

			.SELF(gen[4290]),
			.cell_state(gen[4290])
		); 

/******************* CELL 4291 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4291 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4195]),
			.N(gen[4196]),
			.NE(gen[4197]),

			.O(gen[4290]),
			.E(gen[4292]),

			.SO(gen[4385]),
			.S(gen[4386]),
			.SE(gen[4387]),

			.SELF(gen[4291]),
			.cell_state(gen[4291])
		); 

/******************* CELL 4292 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4292 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4196]),
			.N(gen[4197]),
			.NE(gen[4198]),

			.O(gen[4291]),
			.E(gen[4293]),

			.SO(gen[4386]),
			.S(gen[4387]),
			.SE(gen[4388]),

			.SELF(gen[4292]),
			.cell_state(gen[4292])
		); 

/******************* CELL 4293 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4293 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4197]),
			.N(gen[4198]),
			.NE(gen[4199]),

			.O(gen[4292]),
			.E(gen[4294]),

			.SO(gen[4387]),
			.S(gen[4388]),
			.SE(gen[4389]),

			.SELF(gen[4293]),
			.cell_state(gen[4293])
		); 

/******************* CELL 4294 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4294 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4198]),
			.N(gen[4199]),
			.NE(gen[4200]),

			.O(gen[4293]),
			.E(gen[4295]),

			.SO(gen[4388]),
			.S(gen[4389]),
			.SE(gen[4390]),

			.SELF(gen[4294]),
			.cell_state(gen[4294])
		); 

/******************* CELL 4295 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4295 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4199]),
			.N(gen[4200]),
			.NE(gen[4201]),

			.O(gen[4294]),
			.E(gen[4296]),

			.SO(gen[4389]),
			.S(gen[4390]),
			.SE(gen[4391]),

			.SELF(gen[4295]),
			.cell_state(gen[4295])
		); 

/******************* CELL 4296 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4296 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4200]),
			.N(gen[4201]),
			.NE(gen[4202]),

			.O(gen[4295]),
			.E(gen[4297]),

			.SO(gen[4390]),
			.S(gen[4391]),
			.SE(gen[4392]),

			.SELF(gen[4296]),
			.cell_state(gen[4296])
		); 

/******************* CELL 4297 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4297 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4201]),
			.N(gen[4202]),
			.NE(gen[4203]),

			.O(gen[4296]),
			.E(gen[4298]),

			.SO(gen[4391]),
			.S(gen[4392]),
			.SE(gen[4393]),

			.SELF(gen[4297]),
			.cell_state(gen[4297])
		); 

/******************* CELL 4298 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4298 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4202]),
			.N(gen[4203]),
			.NE(gen[4204]),

			.O(gen[4297]),
			.E(gen[4299]),

			.SO(gen[4392]),
			.S(gen[4393]),
			.SE(gen[4394]),

			.SELF(gen[4298]),
			.cell_state(gen[4298])
		); 

/******************* CELL 4299 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4299 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4203]),
			.N(gen[4204]),
			.NE(gen[4205]),

			.O(gen[4298]),
			.E(gen[4300]),

			.SO(gen[4393]),
			.S(gen[4394]),
			.SE(gen[4395]),

			.SELF(gen[4299]),
			.cell_state(gen[4299])
		); 

/******************* CELL 4300 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4300 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4204]),
			.N(gen[4205]),
			.NE(gen[4206]),

			.O(gen[4299]),
			.E(gen[4301]),

			.SO(gen[4394]),
			.S(gen[4395]),
			.SE(gen[4396]),

			.SELF(gen[4300]),
			.cell_state(gen[4300])
		); 

/******************* CELL 4301 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4301 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4205]),
			.N(gen[4206]),
			.NE(gen[4207]),

			.O(gen[4300]),
			.E(gen[4302]),

			.SO(gen[4395]),
			.S(gen[4396]),
			.SE(gen[4397]),

			.SELF(gen[4301]),
			.cell_state(gen[4301])
		); 

/******************* CELL 4302 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4302 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4206]),
			.N(gen[4207]),
			.NE(gen[4208]),

			.O(gen[4301]),
			.E(gen[4303]),

			.SO(gen[4396]),
			.S(gen[4397]),
			.SE(gen[4398]),

			.SELF(gen[4302]),
			.cell_state(gen[4302])
		); 

/******************* CELL 4303 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4303 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4207]),
			.N(gen[4208]),
			.NE(gen[4209]),

			.O(gen[4302]),
			.E(gen[4304]),

			.SO(gen[4397]),
			.S(gen[4398]),
			.SE(gen[4399]),

			.SELF(gen[4303]),
			.cell_state(gen[4303])
		); 

/******************* CELL 4304 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4304 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4208]),
			.N(gen[4209]),
			.NE(gen[4210]),

			.O(gen[4303]),
			.E(gen[4305]),

			.SO(gen[4398]),
			.S(gen[4399]),
			.SE(gen[4400]),

			.SELF(gen[4304]),
			.cell_state(gen[4304])
		); 

/******************* CELL 4305 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4305 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4209]),
			.N(gen[4210]),
			.NE(gen[4211]),

			.O(gen[4304]),
			.E(gen[4306]),

			.SO(gen[4399]),
			.S(gen[4400]),
			.SE(gen[4401]),

			.SELF(gen[4305]),
			.cell_state(gen[4305])
		); 

/******************* CELL 4306 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4306 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4210]),
			.N(gen[4211]),
			.NE(gen[4212]),

			.O(gen[4305]),
			.E(gen[4307]),

			.SO(gen[4400]),
			.S(gen[4401]),
			.SE(gen[4402]),

			.SELF(gen[4306]),
			.cell_state(gen[4306])
		); 

/******************* CELL 4307 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4307 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4211]),
			.N(gen[4212]),
			.NE(gen[4213]),

			.O(gen[4306]),
			.E(gen[4308]),

			.SO(gen[4401]),
			.S(gen[4402]),
			.SE(gen[4403]),

			.SELF(gen[4307]),
			.cell_state(gen[4307])
		); 

/******************* CELL 4308 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4308 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4212]),
			.N(gen[4213]),
			.NE(gen[4214]),

			.O(gen[4307]),
			.E(gen[4309]),

			.SO(gen[4402]),
			.S(gen[4403]),
			.SE(gen[4404]),

			.SELF(gen[4308]),
			.cell_state(gen[4308])
		); 

/******************* CELL 4309 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4309 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4213]),
			.N(gen[4214]),
			.NE(gen[4215]),

			.O(gen[4308]),
			.E(gen[4310]),

			.SO(gen[4403]),
			.S(gen[4404]),
			.SE(gen[4405]),

			.SELF(gen[4309]),
			.cell_state(gen[4309])
		); 

/******************* CELL 4310 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4310 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4214]),
			.N(gen[4215]),
			.NE(gen[4216]),

			.O(gen[4309]),
			.E(gen[4311]),

			.SO(gen[4404]),
			.S(gen[4405]),
			.SE(gen[4406]),

			.SELF(gen[4310]),
			.cell_state(gen[4310])
		); 

/******************* CELL 4311 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4311 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4215]),
			.N(gen[4216]),
			.NE(gen[4217]),

			.O(gen[4310]),
			.E(gen[4312]),

			.SO(gen[4405]),
			.S(gen[4406]),
			.SE(gen[4407]),

			.SELF(gen[4311]),
			.cell_state(gen[4311])
		); 

/******************* CELL 4312 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4312 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4216]),
			.N(gen[4217]),
			.NE(gen[4218]),

			.O(gen[4311]),
			.E(gen[4313]),

			.SO(gen[4406]),
			.S(gen[4407]),
			.SE(gen[4408]),

			.SELF(gen[4312]),
			.cell_state(gen[4312])
		); 

/******************* CELL 4313 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4313 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4217]),
			.N(gen[4218]),
			.NE(gen[4219]),

			.O(gen[4312]),
			.E(gen[4314]),

			.SO(gen[4407]),
			.S(gen[4408]),
			.SE(gen[4409]),

			.SELF(gen[4313]),
			.cell_state(gen[4313])
		); 

/******************* CELL 4314 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4314 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4218]),
			.N(gen[4219]),
			.NE(gen[4220]),

			.O(gen[4313]),
			.E(gen[4315]),

			.SO(gen[4408]),
			.S(gen[4409]),
			.SE(gen[4410]),

			.SELF(gen[4314]),
			.cell_state(gen[4314])
		); 

/******************* CELL 4315 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4315 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4219]),
			.N(gen[4220]),
			.NE(gen[4221]),

			.O(gen[4314]),
			.E(gen[4316]),

			.SO(gen[4409]),
			.S(gen[4410]),
			.SE(gen[4411]),

			.SELF(gen[4315]),
			.cell_state(gen[4315])
		); 

/******************* CELL 4316 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4316 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4220]),
			.N(gen[4221]),
			.NE(gen[4222]),

			.O(gen[4315]),
			.E(gen[4317]),

			.SO(gen[4410]),
			.S(gen[4411]),
			.SE(gen[4412]),

			.SELF(gen[4316]),
			.cell_state(gen[4316])
		); 

/******************* CELL 4317 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4317 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4221]),
			.N(gen[4222]),
			.NE(gen[4223]),

			.O(gen[4316]),
			.E(gen[4318]),

			.SO(gen[4411]),
			.S(gen[4412]),
			.SE(gen[4413]),

			.SELF(gen[4317]),
			.cell_state(gen[4317])
		); 

/******************* CELL 4318 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4318 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4222]),
			.N(gen[4223]),
			.NE(gen[4224]),

			.O(gen[4317]),
			.E(gen[4319]),

			.SO(gen[4412]),
			.S(gen[4413]),
			.SE(gen[4414]),

			.SELF(gen[4318]),
			.cell_state(gen[4318])
		); 

/******************* CELL 4319 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4319 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4223]),
			.N(gen[4224]),
			.NE(gen[4225]),

			.O(gen[4318]),
			.E(gen[4320]),

			.SO(gen[4413]),
			.S(gen[4414]),
			.SE(gen[4415]),

			.SELF(gen[4319]),
			.cell_state(gen[4319])
		); 

/******************* CELL 4320 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4320 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4224]),
			.N(gen[4225]),
			.NE(gen[4226]),

			.O(gen[4319]),
			.E(gen[4321]),

			.SO(gen[4414]),
			.S(gen[4415]),
			.SE(gen[4416]),

			.SELF(gen[4320]),
			.cell_state(gen[4320])
		); 

/******************* CELL 4321 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4321 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4225]),
			.N(gen[4226]),
			.NE(gen[4227]),

			.O(gen[4320]),
			.E(gen[4322]),

			.SO(gen[4415]),
			.S(gen[4416]),
			.SE(gen[4417]),

			.SELF(gen[4321]),
			.cell_state(gen[4321])
		); 

/******************* CELL 4322 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4322 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4226]),
			.N(gen[4227]),
			.NE(gen[4228]),

			.O(gen[4321]),
			.E(gen[4323]),

			.SO(gen[4416]),
			.S(gen[4417]),
			.SE(gen[4418]),

			.SELF(gen[4322]),
			.cell_state(gen[4322])
		); 

/******************* CELL 4323 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4323 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4227]),
			.N(gen[4228]),
			.NE(gen[4229]),

			.O(gen[4322]),
			.E(gen[4324]),

			.SO(gen[4417]),
			.S(gen[4418]),
			.SE(gen[4419]),

			.SELF(gen[4323]),
			.cell_state(gen[4323])
		); 

/******************* CELL 4324 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4324 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4228]),
			.N(gen[4229]),
			.NE(gen[4230]),

			.O(gen[4323]),
			.E(gen[4325]),

			.SO(gen[4418]),
			.S(gen[4419]),
			.SE(gen[4420]),

			.SELF(gen[4324]),
			.cell_state(gen[4324])
		); 

/******************* CELL 4325 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4325 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4229]),
			.N(gen[4230]),
			.NE(gen[4231]),

			.O(gen[4324]),
			.E(gen[4326]),

			.SO(gen[4419]),
			.S(gen[4420]),
			.SE(gen[4421]),

			.SELF(gen[4325]),
			.cell_state(gen[4325])
		); 

/******************* CELL 4326 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4326 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4230]),
			.N(gen[4231]),
			.NE(gen[4232]),

			.O(gen[4325]),
			.E(gen[4327]),

			.SO(gen[4420]),
			.S(gen[4421]),
			.SE(gen[4422]),

			.SELF(gen[4326]),
			.cell_state(gen[4326])
		); 

/******************* CELL 4327 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4327 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4231]),
			.N(gen[4232]),
			.NE(gen[4233]),

			.O(gen[4326]),
			.E(gen[4328]),

			.SO(gen[4421]),
			.S(gen[4422]),
			.SE(gen[4423]),

			.SELF(gen[4327]),
			.cell_state(gen[4327])
		); 

/******************* CELL 4328 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4328 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4232]),
			.N(gen[4233]),
			.NE(gen[4234]),

			.O(gen[4327]),
			.E(gen[4329]),

			.SO(gen[4422]),
			.S(gen[4423]),
			.SE(gen[4424]),

			.SELF(gen[4328]),
			.cell_state(gen[4328])
		); 

/******************* CELL 4329 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4329 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4233]),
			.N(gen[4234]),
			.NE(gen[4235]),

			.O(gen[4328]),
			.E(gen[4330]),

			.SO(gen[4423]),
			.S(gen[4424]),
			.SE(gen[4425]),

			.SELF(gen[4329]),
			.cell_state(gen[4329])
		); 

/******************* CELL 4330 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4330 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4234]),
			.N(gen[4235]),
			.NE(gen[4236]),

			.O(gen[4329]),
			.E(gen[4331]),

			.SO(gen[4424]),
			.S(gen[4425]),
			.SE(gen[4426]),

			.SELF(gen[4330]),
			.cell_state(gen[4330])
		); 

/******************* CELL 4331 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4331 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4235]),
			.N(gen[4236]),
			.NE(gen[4237]),

			.O(gen[4330]),
			.E(gen[4332]),

			.SO(gen[4425]),
			.S(gen[4426]),
			.SE(gen[4427]),

			.SELF(gen[4331]),
			.cell_state(gen[4331])
		); 

/******************* CELL 4332 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4332 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4236]),
			.N(gen[4237]),
			.NE(gen[4238]),

			.O(gen[4331]),
			.E(gen[4333]),

			.SO(gen[4426]),
			.S(gen[4427]),
			.SE(gen[4428]),

			.SELF(gen[4332]),
			.cell_state(gen[4332])
		); 

/******************* CELL 4333 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4333 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4237]),
			.N(gen[4238]),
			.NE(gen[4239]),

			.O(gen[4332]),
			.E(gen[4334]),

			.SO(gen[4427]),
			.S(gen[4428]),
			.SE(gen[4429]),

			.SELF(gen[4333]),
			.cell_state(gen[4333])
		); 

/******************* CELL 4334 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4334 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4238]),
			.N(gen[4239]),
			.NE(gen[4240]),

			.O(gen[4333]),
			.E(gen[4335]),

			.SO(gen[4428]),
			.S(gen[4429]),
			.SE(gen[4430]),

			.SELF(gen[4334]),
			.cell_state(gen[4334])
		); 

/******************* CELL 4335 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4335 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4239]),
			.N(gen[4240]),
			.NE(gen[4241]),

			.O(gen[4334]),
			.E(gen[4336]),

			.SO(gen[4429]),
			.S(gen[4430]),
			.SE(gen[4431]),

			.SELF(gen[4335]),
			.cell_state(gen[4335])
		); 

/******************* CELL 4336 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4336 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4240]),
			.N(gen[4241]),
			.NE(gen[4242]),

			.O(gen[4335]),
			.E(gen[4337]),

			.SO(gen[4430]),
			.S(gen[4431]),
			.SE(gen[4432]),

			.SELF(gen[4336]),
			.cell_state(gen[4336])
		); 

/******************* CELL 4337 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4337 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4241]),
			.N(gen[4242]),
			.NE(gen[4243]),

			.O(gen[4336]),
			.E(gen[4338]),

			.SO(gen[4431]),
			.S(gen[4432]),
			.SE(gen[4433]),

			.SELF(gen[4337]),
			.cell_state(gen[4337])
		); 

/******************* CELL 4338 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4338 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4242]),
			.N(gen[4243]),
			.NE(gen[4244]),

			.O(gen[4337]),
			.E(gen[4339]),

			.SO(gen[4432]),
			.S(gen[4433]),
			.SE(gen[4434]),

			.SELF(gen[4338]),
			.cell_state(gen[4338])
		); 

/******************* CELL 4339 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4339 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4243]),
			.N(gen[4244]),
			.NE(gen[4245]),

			.O(gen[4338]),
			.E(gen[4340]),

			.SO(gen[4433]),
			.S(gen[4434]),
			.SE(gen[4435]),

			.SELF(gen[4339]),
			.cell_state(gen[4339])
		); 

/******************* CELL 4340 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4340 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4244]),
			.N(gen[4245]),
			.NE(gen[4246]),

			.O(gen[4339]),
			.E(gen[4341]),

			.SO(gen[4434]),
			.S(gen[4435]),
			.SE(gen[4436]),

			.SELF(gen[4340]),
			.cell_state(gen[4340])
		); 

/******************* CELL 4341 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4341 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4245]),
			.N(gen[4246]),
			.NE(gen[4247]),

			.O(gen[4340]),
			.E(gen[4342]),

			.SO(gen[4435]),
			.S(gen[4436]),
			.SE(gen[4437]),

			.SELF(gen[4341]),
			.cell_state(gen[4341])
		); 

/******************* CELL 4342 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4342 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4246]),
			.N(gen[4247]),
			.NE(gen[4248]),

			.O(gen[4341]),
			.E(gen[4343]),

			.SO(gen[4436]),
			.S(gen[4437]),
			.SE(gen[4438]),

			.SELF(gen[4342]),
			.cell_state(gen[4342])
		); 

/******************* CELL 4343 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4343 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4247]),
			.N(gen[4248]),
			.NE(gen[4249]),

			.O(gen[4342]),
			.E(gen[4344]),

			.SO(gen[4437]),
			.S(gen[4438]),
			.SE(gen[4439]),

			.SELF(gen[4343]),
			.cell_state(gen[4343])
		); 

/******************* CELL 4344 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4344 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4248]),
			.N(gen[4249]),
			.NE(gen[4250]),

			.O(gen[4343]),
			.E(gen[4345]),

			.SO(gen[4438]),
			.S(gen[4439]),
			.SE(gen[4440]),

			.SELF(gen[4344]),
			.cell_state(gen[4344])
		); 

/******************* CELL 4345 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4345 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4249]),
			.N(gen[4250]),
			.NE(gen[4251]),

			.O(gen[4344]),
			.E(gen[4346]),

			.SO(gen[4439]),
			.S(gen[4440]),
			.SE(gen[4441]),

			.SELF(gen[4345]),
			.cell_state(gen[4345])
		); 

/******************* CELL 4346 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4346 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4250]),
			.N(gen[4251]),
			.NE(gen[4252]),

			.O(gen[4345]),
			.E(gen[4347]),

			.SO(gen[4440]),
			.S(gen[4441]),
			.SE(gen[4442]),

			.SELF(gen[4346]),
			.cell_state(gen[4346])
		); 

/******************* CELL 4347 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4347 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4251]),
			.N(gen[4252]),
			.NE(gen[4253]),

			.O(gen[4346]),
			.E(gen[4348]),

			.SO(gen[4441]),
			.S(gen[4442]),
			.SE(gen[4443]),

			.SELF(gen[4347]),
			.cell_state(gen[4347])
		); 

/******************* CELL 4348 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4348 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4252]),
			.N(gen[4253]),
			.NE(gen[4254]),

			.O(gen[4347]),
			.E(gen[4349]),

			.SO(gen[4442]),
			.S(gen[4443]),
			.SE(gen[4444]),

			.SELF(gen[4348]),
			.cell_state(gen[4348])
		); 

/******************* CELL 4349 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4349 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4253]),
			.N(gen[4254]),
			.NE(gen[4255]),

			.O(gen[4348]),
			.E(gen[4350]),

			.SO(gen[4443]),
			.S(gen[4444]),
			.SE(gen[4445]),

			.SELF(gen[4349]),
			.cell_state(gen[4349])
		); 

/******************* CELL 4350 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4350 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4254]),
			.N(gen[4255]),
			.NE(gen[4256]),

			.O(gen[4349]),
			.E(gen[4351]),

			.SO(gen[4444]),
			.S(gen[4445]),
			.SE(gen[4446]),

			.SELF(gen[4350]),
			.cell_state(gen[4350])
		); 

/******************* CELL 4351 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4351 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4255]),
			.N(gen[4256]),
			.NE(gen[4257]),

			.O(gen[4350]),
			.E(gen[4352]),

			.SO(gen[4445]),
			.S(gen[4446]),
			.SE(gen[4447]),

			.SELF(gen[4351]),
			.cell_state(gen[4351])
		); 

/******************* CELL 4352 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4352 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4256]),
			.N(gen[4257]),
			.NE(gen[4258]),

			.O(gen[4351]),
			.E(gen[4353]),

			.SO(gen[4446]),
			.S(gen[4447]),
			.SE(gen[4448]),

			.SELF(gen[4352]),
			.cell_state(gen[4352])
		); 

/******************* CELL 4353 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4353 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4257]),
			.N(gen[4258]),
			.NE(gen[4259]),

			.O(gen[4352]),
			.E(gen[4354]),

			.SO(gen[4447]),
			.S(gen[4448]),
			.SE(gen[4449]),

			.SELF(gen[4353]),
			.cell_state(gen[4353])
		); 

/******************* CELL 4354 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4354 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4258]),
			.N(gen[4259]),
			.NE(gen[4260]),

			.O(gen[4353]),
			.E(gen[4355]),

			.SO(gen[4448]),
			.S(gen[4449]),
			.SE(gen[4450]),

			.SELF(gen[4354]),
			.cell_state(gen[4354])
		); 

/******************* CELL 4355 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4355 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4259]),
			.N(gen[4260]),
			.NE(gen[4261]),

			.O(gen[4354]),
			.E(gen[4356]),

			.SO(gen[4449]),
			.S(gen[4450]),
			.SE(gen[4451]),

			.SELF(gen[4355]),
			.cell_state(gen[4355])
		); 

/******************* CELL 4356 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4356 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4260]),
			.N(gen[4261]),
			.NE(gen[4262]),

			.O(gen[4355]),
			.E(gen[4357]),

			.SO(gen[4450]),
			.S(gen[4451]),
			.SE(gen[4452]),

			.SELF(gen[4356]),
			.cell_state(gen[4356])
		); 

/******************* CELL 4357 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4357 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4261]),
			.N(gen[4262]),
			.NE(gen[4263]),

			.O(gen[4356]),
			.E(gen[4358]),

			.SO(gen[4451]),
			.S(gen[4452]),
			.SE(gen[4453]),

			.SELF(gen[4357]),
			.cell_state(gen[4357])
		); 

/******************* CELL 4358 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4358 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4262]),
			.N(gen[4263]),
			.NE(gen[4264]),

			.O(gen[4357]),
			.E(gen[4359]),

			.SO(gen[4452]),
			.S(gen[4453]),
			.SE(gen[4454]),

			.SELF(gen[4358]),
			.cell_state(gen[4358])
		); 

/******************* CELL 4359 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4359 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4263]),
			.N(gen[4264]),
			.NE(gen[4265]),

			.O(gen[4358]),
			.E(gen[4360]),

			.SO(gen[4453]),
			.S(gen[4454]),
			.SE(gen[4455]),

			.SELF(gen[4359]),
			.cell_state(gen[4359])
		); 

/******************* CELL 4360 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4360 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4264]),
			.N(gen[4265]),
			.NE(gen[4266]),

			.O(gen[4359]),
			.E(gen[4361]),

			.SO(gen[4454]),
			.S(gen[4455]),
			.SE(gen[4456]),

			.SELF(gen[4360]),
			.cell_state(gen[4360])
		); 

/******************* CELL 4361 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4361 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4265]),
			.N(gen[4266]),
			.NE(gen[4267]),

			.O(gen[4360]),
			.E(gen[4362]),

			.SO(gen[4455]),
			.S(gen[4456]),
			.SE(gen[4457]),

			.SELF(gen[4361]),
			.cell_state(gen[4361])
		); 

/******************* CELL 4362 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4362 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4266]),
			.N(gen[4267]),
			.NE(gen[4268]),

			.O(gen[4361]),
			.E(gen[4363]),

			.SO(gen[4456]),
			.S(gen[4457]),
			.SE(gen[4458]),

			.SELF(gen[4362]),
			.cell_state(gen[4362])
		); 

/******************* CELL 4363 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4363 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4267]),
			.N(gen[4268]),
			.NE(gen[4269]),

			.O(gen[4362]),
			.E(gen[4364]),

			.SO(gen[4457]),
			.S(gen[4458]),
			.SE(gen[4459]),

			.SELF(gen[4363]),
			.cell_state(gen[4363])
		); 

/******************* CELL 4364 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4364 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4268]),
			.N(gen[4269]),
			.NE(gen[4270]),

			.O(gen[4363]),
			.E(gen[4365]),

			.SO(gen[4458]),
			.S(gen[4459]),
			.SE(gen[4460]),

			.SELF(gen[4364]),
			.cell_state(gen[4364])
		); 

/******************* CELL 4365 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4365 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4269]),
			.N(gen[4270]),
			.NE(gen[4271]),

			.O(gen[4364]),
			.E(gen[4366]),

			.SO(gen[4459]),
			.S(gen[4460]),
			.SE(gen[4461]),

			.SELF(gen[4365]),
			.cell_state(gen[4365])
		); 

/******************* CELL 4366 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4366 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4270]),
			.N(gen[4271]),
			.NE(gen[4272]),

			.O(gen[4365]),
			.E(gen[4367]),

			.SO(gen[4460]),
			.S(gen[4461]),
			.SE(gen[4462]),

			.SELF(gen[4366]),
			.cell_state(gen[4366])
		); 

/******************* CELL 4367 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4367 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4271]),
			.N(gen[4272]),
			.NE(gen[4273]),

			.O(gen[4366]),
			.E(gen[4368]),

			.SO(gen[4461]),
			.S(gen[4462]),
			.SE(gen[4463]),

			.SELF(gen[4367]),
			.cell_state(gen[4367])
		); 

/******************* CELL 4368 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4368 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4272]),
			.N(gen[4273]),
			.NE(gen[4274]),

			.O(gen[4367]),
			.E(gen[4369]),

			.SO(gen[4462]),
			.S(gen[4463]),
			.SE(gen[4464]),

			.SELF(gen[4368]),
			.cell_state(gen[4368])
		); 

/******************* CELL 4369 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4369 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4273]),
			.N(gen[4274]),
			.NE(gen[4273]),

			.O(gen[4368]),
			.E(gen[4368]),

			.SO(gen[4463]),
			.S(gen[4464]),
			.SE(gen[4463]),

			.SELF(gen[4369]),
			.cell_state(gen[4369])
		); 

/******************* CELL 4370 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4370 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4276]),
			.N(gen[4275]),
			.NE(gen[4276]),

			.O(gen[4371]),
			.E(gen[4371]),

			.SO(gen[4466]),
			.S(gen[4465]),
			.SE(gen[4466]),

			.SELF(gen[4370]),
			.cell_state(gen[4370])
		); 

/******************* CELL 4371 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4371 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4275]),
			.N(gen[4276]),
			.NE(gen[4277]),

			.O(gen[4370]),
			.E(gen[4372]),

			.SO(gen[4465]),
			.S(gen[4466]),
			.SE(gen[4467]),

			.SELF(gen[4371]),
			.cell_state(gen[4371])
		); 

/******************* CELL 4372 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4372 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4276]),
			.N(gen[4277]),
			.NE(gen[4278]),

			.O(gen[4371]),
			.E(gen[4373]),

			.SO(gen[4466]),
			.S(gen[4467]),
			.SE(gen[4468]),

			.SELF(gen[4372]),
			.cell_state(gen[4372])
		); 

/******************* CELL 4373 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4373 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4277]),
			.N(gen[4278]),
			.NE(gen[4279]),

			.O(gen[4372]),
			.E(gen[4374]),

			.SO(gen[4467]),
			.S(gen[4468]),
			.SE(gen[4469]),

			.SELF(gen[4373]),
			.cell_state(gen[4373])
		); 

/******************* CELL 4374 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4374 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4278]),
			.N(gen[4279]),
			.NE(gen[4280]),

			.O(gen[4373]),
			.E(gen[4375]),

			.SO(gen[4468]),
			.S(gen[4469]),
			.SE(gen[4470]),

			.SELF(gen[4374]),
			.cell_state(gen[4374])
		); 

/******************* CELL 4375 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4375 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4279]),
			.N(gen[4280]),
			.NE(gen[4281]),

			.O(gen[4374]),
			.E(gen[4376]),

			.SO(gen[4469]),
			.S(gen[4470]),
			.SE(gen[4471]),

			.SELF(gen[4375]),
			.cell_state(gen[4375])
		); 

/******************* CELL 4376 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4376 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4280]),
			.N(gen[4281]),
			.NE(gen[4282]),

			.O(gen[4375]),
			.E(gen[4377]),

			.SO(gen[4470]),
			.S(gen[4471]),
			.SE(gen[4472]),

			.SELF(gen[4376]),
			.cell_state(gen[4376])
		); 

/******************* CELL 4377 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4377 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4281]),
			.N(gen[4282]),
			.NE(gen[4283]),

			.O(gen[4376]),
			.E(gen[4378]),

			.SO(gen[4471]),
			.S(gen[4472]),
			.SE(gen[4473]),

			.SELF(gen[4377]),
			.cell_state(gen[4377])
		); 

/******************* CELL 4378 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4378 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4282]),
			.N(gen[4283]),
			.NE(gen[4284]),

			.O(gen[4377]),
			.E(gen[4379]),

			.SO(gen[4472]),
			.S(gen[4473]),
			.SE(gen[4474]),

			.SELF(gen[4378]),
			.cell_state(gen[4378])
		); 

/******************* CELL 4379 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4379 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4283]),
			.N(gen[4284]),
			.NE(gen[4285]),

			.O(gen[4378]),
			.E(gen[4380]),

			.SO(gen[4473]),
			.S(gen[4474]),
			.SE(gen[4475]),

			.SELF(gen[4379]),
			.cell_state(gen[4379])
		); 

/******************* CELL 4380 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4380 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4284]),
			.N(gen[4285]),
			.NE(gen[4286]),

			.O(gen[4379]),
			.E(gen[4381]),

			.SO(gen[4474]),
			.S(gen[4475]),
			.SE(gen[4476]),

			.SELF(gen[4380]),
			.cell_state(gen[4380])
		); 

/******************* CELL 4381 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4381 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4285]),
			.N(gen[4286]),
			.NE(gen[4287]),

			.O(gen[4380]),
			.E(gen[4382]),

			.SO(gen[4475]),
			.S(gen[4476]),
			.SE(gen[4477]),

			.SELF(gen[4381]),
			.cell_state(gen[4381])
		); 

/******************* CELL 4382 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4382 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4286]),
			.N(gen[4287]),
			.NE(gen[4288]),

			.O(gen[4381]),
			.E(gen[4383]),

			.SO(gen[4476]),
			.S(gen[4477]),
			.SE(gen[4478]),

			.SELF(gen[4382]),
			.cell_state(gen[4382])
		); 

/******************* CELL 4383 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4383 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4287]),
			.N(gen[4288]),
			.NE(gen[4289]),

			.O(gen[4382]),
			.E(gen[4384]),

			.SO(gen[4477]),
			.S(gen[4478]),
			.SE(gen[4479]),

			.SELF(gen[4383]),
			.cell_state(gen[4383])
		); 

/******************* CELL 4384 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4384 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4288]),
			.N(gen[4289]),
			.NE(gen[4290]),

			.O(gen[4383]),
			.E(gen[4385]),

			.SO(gen[4478]),
			.S(gen[4479]),
			.SE(gen[4480]),

			.SELF(gen[4384]),
			.cell_state(gen[4384])
		); 

/******************* CELL 4385 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4385 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4289]),
			.N(gen[4290]),
			.NE(gen[4291]),

			.O(gen[4384]),
			.E(gen[4386]),

			.SO(gen[4479]),
			.S(gen[4480]),
			.SE(gen[4481]),

			.SELF(gen[4385]),
			.cell_state(gen[4385])
		); 

/******************* CELL 4386 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4386 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4290]),
			.N(gen[4291]),
			.NE(gen[4292]),

			.O(gen[4385]),
			.E(gen[4387]),

			.SO(gen[4480]),
			.S(gen[4481]),
			.SE(gen[4482]),

			.SELF(gen[4386]),
			.cell_state(gen[4386])
		); 

/******************* CELL 4387 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4387 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4291]),
			.N(gen[4292]),
			.NE(gen[4293]),

			.O(gen[4386]),
			.E(gen[4388]),

			.SO(gen[4481]),
			.S(gen[4482]),
			.SE(gen[4483]),

			.SELF(gen[4387]),
			.cell_state(gen[4387])
		); 

/******************* CELL 4388 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4388 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4292]),
			.N(gen[4293]),
			.NE(gen[4294]),

			.O(gen[4387]),
			.E(gen[4389]),

			.SO(gen[4482]),
			.S(gen[4483]),
			.SE(gen[4484]),

			.SELF(gen[4388]),
			.cell_state(gen[4388])
		); 

/******************* CELL 4389 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4389 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4293]),
			.N(gen[4294]),
			.NE(gen[4295]),

			.O(gen[4388]),
			.E(gen[4390]),

			.SO(gen[4483]),
			.S(gen[4484]),
			.SE(gen[4485]),

			.SELF(gen[4389]),
			.cell_state(gen[4389])
		); 

/******************* CELL 4390 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4390 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4294]),
			.N(gen[4295]),
			.NE(gen[4296]),

			.O(gen[4389]),
			.E(gen[4391]),

			.SO(gen[4484]),
			.S(gen[4485]),
			.SE(gen[4486]),

			.SELF(gen[4390]),
			.cell_state(gen[4390])
		); 

/******************* CELL 4391 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4391 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4295]),
			.N(gen[4296]),
			.NE(gen[4297]),

			.O(gen[4390]),
			.E(gen[4392]),

			.SO(gen[4485]),
			.S(gen[4486]),
			.SE(gen[4487]),

			.SELF(gen[4391]),
			.cell_state(gen[4391])
		); 

/******************* CELL 4392 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4392 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4296]),
			.N(gen[4297]),
			.NE(gen[4298]),

			.O(gen[4391]),
			.E(gen[4393]),

			.SO(gen[4486]),
			.S(gen[4487]),
			.SE(gen[4488]),

			.SELF(gen[4392]),
			.cell_state(gen[4392])
		); 

/******************* CELL 4393 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4393 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4297]),
			.N(gen[4298]),
			.NE(gen[4299]),

			.O(gen[4392]),
			.E(gen[4394]),

			.SO(gen[4487]),
			.S(gen[4488]),
			.SE(gen[4489]),

			.SELF(gen[4393]),
			.cell_state(gen[4393])
		); 

/******************* CELL 4394 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4394 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4298]),
			.N(gen[4299]),
			.NE(gen[4300]),

			.O(gen[4393]),
			.E(gen[4395]),

			.SO(gen[4488]),
			.S(gen[4489]),
			.SE(gen[4490]),

			.SELF(gen[4394]),
			.cell_state(gen[4394])
		); 

/******************* CELL 4395 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4395 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4299]),
			.N(gen[4300]),
			.NE(gen[4301]),

			.O(gen[4394]),
			.E(gen[4396]),

			.SO(gen[4489]),
			.S(gen[4490]),
			.SE(gen[4491]),

			.SELF(gen[4395]),
			.cell_state(gen[4395])
		); 

/******************* CELL 4396 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4396 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4300]),
			.N(gen[4301]),
			.NE(gen[4302]),

			.O(gen[4395]),
			.E(gen[4397]),

			.SO(gen[4490]),
			.S(gen[4491]),
			.SE(gen[4492]),

			.SELF(gen[4396]),
			.cell_state(gen[4396])
		); 

/******************* CELL 4397 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4397 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4301]),
			.N(gen[4302]),
			.NE(gen[4303]),

			.O(gen[4396]),
			.E(gen[4398]),

			.SO(gen[4491]),
			.S(gen[4492]),
			.SE(gen[4493]),

			.SELF(gen[4397]),
			.cell_state(gen[4397])
		); 

/******************* CELL 4398 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4398 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4302]),
			.N(gen[4303]),
			.NE(gen[4304]),

			.O(gen[4397]),
			.E(gen[4399]),

			.SO(gen[4492]),
			.S(gen[4493]),
			.SE(gen[4494]),

			.SELF(gen[4398]),
			.cell_state(gen[4398])
		); 

/******************* CELL 4399 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4399 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4303]),
			.N(gen[4304]),
			.NE(gen[4305]),

			.O(gen[4398]),
			.E(gen[4400]),

			.SO(gen[4493]),
			.S(gen[4494]),
			.SE(gen[4495]),

			.SELF(gen[4399]),
			.cell_state(gen[4399])
		); 

/******************* CELL 4400 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4400 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4304]),
			.N(gen[4305]),
			.NE(gen[4306]),

			.O(gen[4399]),
			.E(gen[4401]),

			.SO(gen[4494]),
			.S(gen[4495]),
			.SE(gen[4496]),

			.SELF(gen[4400]),
			.cell_state(gen[4400])
		); 

/******************* CELL 4401 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4401 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4305]),
			.N(gen[4306]),
			.NE(gen[4307]),

			.O(gen[4400]),
			.E(gen[4402]),

			.SO(gen[4495]),
			.S(gen[4496]),
			.SE(gen[4497]),

			.SELF(gen[4401]),
			.cell_state(gen[4401])
		); 

/******************* CELL 4402 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4402 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4306]),
			.N(gen[4307]),
			.NE(gen[4308]),

			.O(gen[4401]),
			.E(gen[4403]),

			.SO(gen[4496]),
			.S(gen[4497]),
			.SE(gen[4498]),

			.SELF(gen[4402]),
			.cell_state(gen[4402])
		); 

/******************* CELL 4403 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4403 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4307]),
			.N(gen[4308]),
			.NE(gen[4309]),

			.O(gen[4402]),
			.E(gen[4404]),

			.SO(gen[4497]),
			.S(gen[4498]),
			.SE(gen[4499]),

			.SELF(gen[4403]),
			.cell_state(gen[4403])
		); 

/******************* CELL 4404 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4404 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4308]),
			.N(gen[4309]),
			.NE(gen[4310]),

			.O(gen[4403]),
			.E(gen[4405]),

			.SO(gen[4498]),
			.S(gen[4499]),
			.SE(gen[4500]),

			.SELF(gen[4404]),
			.cell_state(gen[4404])
		); 

/******************* CELL 4405 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4405 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4309]),
			.N(gen[4310]),
			.NE(gen[4311]),

			.O(gen[4404]),
			.E(gen[4406]),

			.SO(gen[4499]),
			.S(gen[4500]),
			.SE(gen[4501]),

			.SELF(gen[4405]),
			.cell_state(gen[4405])
		); 

/******************* CELL 4406 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4406 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4310]),
			.N(gen[4311]),
			.NE(gen[4312]),

			.O(gen[4405]),
			.E(gen[4407]),

			.SO(gen[4500]),
			.S(gen[4501]),
			.SE(gen[4502]),

			.SELF(gen[4406]),
			.cell_state(gen[4406])
		); 

/******************* CELL 4407 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4407 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4311]),
			.N(gen[4312]),
			.NE(gen[4313]),

			.O(gen[4406]),
			.E(gen[4408]),

			.SO(gen[4501]),
			.S(gen[4502]),
			.SE(gen[4503]),

			.SELF(gen[4407]),
			.cell_state(gen[4407])
		); 

/******************* CELL 4408 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4408 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4312]),
			.N(gen[4313]),
			.NE(gen[4314]),

			.O(gen[4407]),
			.E(gen[4409]),

			.SO(gen[4502]),
			.S(gen[4503]),
			.SE(gen[4504]),

			.SELF(gen[4408]),
			.cell_state(gen[4408])
		); 

/******************* CELL 4409 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4409 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4313]),
			.N(gen[4314]),
			.NE(gen[4315]),

			.O(gen[4408]),
			.E(gen[4410]),

			.SO(gen[4503]),
			.S(gen[4504]),
			.SE(gen[4505]),

			.SELF(gen[4409]),
			.cell_state(gen[4409])
		); 

/******************* CELL 4410 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4410 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4314]),
			.N(gen[4315]),
			.NE(gen[4316]),

			.O(gen[4409]),
			.E(gen[4411]),

			.SO(gen[4504]),
			.S(gen[4505]),
			.SE(gen[4506]),

			.SELF(gen[4410]),
			.cell_state(gen[4410])
		); 

/******************* CELL 4411 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4411 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4315]),
			.N(gen[4316]),
			.NE(gen[4317]),

			.O(gen[4410]),
			.E(gen[4412]),

			.SO(gen[4505]),
			.S(gen[4506]),
			.SE(gen[4507]),

			.SELF(gen[4411]),
			.cell_state(gen[4411])
		); 

/******************* CELL 4412 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4412 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4316]),
			.N(gen[4317]),
			.NE(gen[4318]),

			.O(gen[4411]),
			.E(gen[4413]),

			.SO(gen[4506]),
			.S(gen[4507]),
			.SE(gen[4508]),

			.SELF(gen[4412]),
			.cell_state(gen[4412])
		); 

/******************* CELL 4413 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4413 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4317]),
			.N(gen[4318]),
			.NE(gen[4319]),

			.O(gen[4412]),
			.E(gen[4414]),

			.SO(gen[4507]),
			.S(gen[4508]),
			.SE(gen[4509]),

			.SELF(gen[4413]),
			.cell_state(gen[4413])
		); 

/******************* CELL 4414 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4414 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4318]),
			.N(gen[4319]),
			.NE(gen[4320]),

			.O(gen[4413]),
			.E(gen[4415]),

			.SO(gen[4508]),
			.S(gen[4509]),
			.SE(gen[4510]),

			.SELF(gen[4414]),
			.cell_state(gen[4414])
		); 

/******************* CELL 4415 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4415 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4319]),
			.N(gen[4320]),
			.NE(gen[4321]),

			.O(gen[4414]),
			.E(gen[4416]),

			.SO(gen[4509]),
			.S(gen[4510]),
			.SE(gen[4511]),

			.SELF(gen[4415]),
			.cell_state(gen[4415])
		); 

/******************* CELL 4416 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4416 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4320]),
			.N(gen[4321]),
			.NE(gen[4322]),

			.O(gen[4415]),
			.E(gen[4417]),

			.SO(gen[4510]),
			.S(gen[4511]),
			.SE(gen[4512]),

			.SELF(gen[4416]),
			.cell_state(gen[4416])
		); 

/******************* CELL 4417 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4417 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4321]),
			.N(gen[4322]),
			.NE(gen[4323]),

			.O(gen[4416]),
			.E(gen[4418]),

			.SO(gen[4511]),
			.S(gen[4512]),
			.SE(gen[4513]),

			.SELF(gen[4417]),
			.cell_state(gen[4417])
		); 

/******************* CELL 4418 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4418 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4322]),
			.N(gen[4323]),
			.NE(gen[4324]),

			.O(gen[4417]),
			.E(gen[4419]),

			.SO(gen[4512]),
			.S(gen[4513]),
			.SE(gen[4514]),

			.SELF(gen[4418]),
			.cell_state(gen[4418])
		); 

/******************* CELL 4419 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4419 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4323]),
			.N(gen[4324]),
			.NE(gen[4325]),

			.O(gen[4418]),
			.E(gen[4420]),

			.SO(gen[4513]),
			.S(gen[4514]),
			.SE(gen[4515]),

			.SELF(gen[4419]),
			.cell_state(gen[4419])
		); 

/******************* CELL 4420 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4420 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4324]),
			.N(gen[4325]),
			.NE(gen[4326]),

			.O(gen[4419]),
			.E(gen[4421]),

			.SO(gen[4514]),
			.S(gen[4515]),
			.SE(gen[4516]),

			.SELF(gen[4420]),
			.cell_state(gen[4420])
		); 

/******************* CELL 4421 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4421 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4325]),
			.N(gen[4326]),
			.NE(gen[4327]),

			.O(gen[4420]),
			.E(gen[4422]),

			.SO(gen[4515]),
			.S(gen[4516]),
			.SE(gen[4517]),

			.SELF(gen[4421]),
			.cell_state(gen[4421])
		); 

/******************* CELL 4422 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4422 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4326]),
			.N(gen[4327]),
			.NE(gen[4328]),

			.O(gen[4421]),
			.E(gen[4423]),

			.SO(gen[4516]),
			.S(gen[4517]),
			.SE(gen[4518]),

			.SELF(gen[4422]),
			.cell_state(gen[4422])
		); 

/******************* CELL 4423 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4423 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4327]),
			.N(gen[4328]),
			.NE(gen[4329]),

			.O(gen[4422]),
			.E(gen[4424]),

			.SO(gen[4517]),
			.S(gen[4518]),
			.SE(gen[4519]),

			.SELF(gen[4423]),
			.cell_state(gen[4423])
		); 

/******************* CELL 4424 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4424 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4328]),
			.N(gen[4329]),
			.NE(gen[4330]),

			.O(gen[4423]),
			.E(gen[4425]),

			.SO(gen[4518]),
			.S(gen[4519]),
			.SE(gen[4520]),

			.SELF(gen[4424]),
			.cell_state(gen[4424])
		); 

/******************* CELL 4425 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4425 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4329]),
			.N(gen[4330]),
			.NE(gen[4331]),

			.O(gen[4424]),
			.E(gen[4426]),

			.SO(gen[4519]),
			.S(gen[4520]),
			.SE(gen[4521]),

			.SELF(gen[4425]),
			.cell_state(gen[4425])
		); 

/******************* CELL 4426 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4426 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4330]),
			.N(gen[4331]),
			.NE(gen[4332]),

			.O(gen[4425]),
			.E(gen[4427]),

			.SO(gen[4520]),
			.S(gen[4521]),
			.SE(gen[4522]),

			.SELF(gen[4426]),
			.cell_state(gen[4426])
		); 

/******************* CELL 4427 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4427 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4331]),
			.N(gen[4332]),
			.NE(gen[4333]),

			.O(gen[4426]),
			.E(gen[4428]),

			.SO(gen[4521]),
			.S(gen[4522]),
			.SE(gen[4523]),

			.SELF(gen[4427]),
			.cell_state(gen[4427])
		); 

/******************* CELL 4428 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4428 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4332]),
			.N(gen[4333]),
			.NE(gen[4334]),

			.O(gen[4427]),
			.E(gen[4429]),

			.SO(gen[4522]),
			.S(gen[4523]),
			.SE(gen[4524]),

			.SELF(gen[4428]),
			.cell_state(gen[4428])
		); 

/******************* CELL 4429 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4429 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4333]),
			.N(gen[4334]),
			.NE(gen[4335]),

			.O(gen[4428]),
			.E(gen[4430]),

			.SO(gen[4523]),
			.S(gen[4524]),
			.SE(gen[4525]),

			.SELF(gen[4429]),
			.cell_state(gen[4429])
		); 

/******************* CELL 4430 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4430 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4334]),
			.N(gen[4335]),
			.NE(gen[4336]),

			.O(gen[4429]),
			.E(gen[4431]),

			.SO(gen[4524]),
			.S(gen[4525]),
			.SE(gen[4526]),

			.SELF(gen[4430]),
			.cell_state(gen[4430])
		); 

/******************* CELL 4431 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4431 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4335]),
			.N(gen[4336]),
			.NE(gen[4337]),

			.O(gen[4430]),
			.E(gen[4432]),

			.SO(gen[4525]),
			.S(gen[4526]),
			.SE(gen[4527]),

			.SELF(gen[4431]),
			.cell_state(gen[4431])
		); 

/******************* CELL 4432 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4432 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4336]),
			.N(gen[4337]),
			.NE(gen[4338]),

			.O(gen[4431]),
			.E(gen[4433]),

			.SO(gen[4526]),
			.S(gen[4527]),
			.SE(gen[4528]),

			.SELF(gen[4432]),
			.cell_state(gen[4432])
		); 

/******************* CELL 4433 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4433 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4337]),
			.N(gen[4338]),
			.NE(gen[4339]),

			.O(gen[4432]),
			.E(gen[4434]),

			.SO(gen[4527]),
			.S(gen[4528]),
			.SE(gen[4529]),

			.SELF(gen[4433]),
			.cell_state(gen[4433])
		); 

/******************* CELL 4434 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4434 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4338]),
			.N(gen[4339]),
			.NE(gen[4340]),

			.O(gen[4433]),
			.E(gen[4435]),

			.SO(gen[4528]),
			.S(gen[4529]),
			.SE(gen[4530]),

			.SELF(gen[4434]),
			.cell_state(gen[4434])
		); 

/******************* CELL 4435 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4435 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4339]),
			.N(gen[4340]),
			.NE(gen[4341]),

			.O(gen[4434]),
			.E(gen[4436]),

			.SO(gen[4529]),
			.S(gen[4530]),
			.SE(gen[4531]),

			.SELF(gen[4435]),
			.cell_state(gen[4435])
		); 

/******************* CELL 4436 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4436 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4340]),
			.N(gen[4341]),
			.NE(gen[4342]),

			.O(gen[4435]),
			.E(gen[4437]),

			.SO(gen[4530]),
			.S(gen[4531]),
			.SE(gen[4532]),

			.SELF(gen[4436]),
			.cell_state(gen[4436])
		); 

/******************* CELL 4437 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4437 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4341]),
			.N(gen[4342]),
			.NE(gen[4343]),

			.O(gen[4436]),
			.E(gen[4438]),

			.SO(gen[4531]),
			.S(gen[4532]),
			.SE(gen[4533]),

			.SELF(gen[4437]),
			.cell_state(gen[4437])
		); 

/******************* CELL 4438 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4438 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4342]),
			.N(gen[4343]),
			.NE(gen[4344]),

			.O(gen[4437]),
			.E(gen[4439]),

			.SO(gen[4532]),
			.S(gen[4533]),
			.SE(gen[4534]),

			.SELF(gen[4438]),
			.cell_state(gen[4438])
		); 

/******************* CELL 4439 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4439 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4343]),
			.N(gen[4344]),
			.NE(gen[4345]),

			.O(gen[4438]),
			.E(gen[4440]),

			.SO(gen[4533]),
			.S(gen[4534]),
			.SE(gen[4535]),

			.SELF(gen[4439]),
			.cell_state(gen[4439])
		); 

/******************* CELL 4440 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4440 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4344]),
			.N(gen[4345]),
			.NE(gen[4346]),

			.O(gen[4439]),
			.E(gen[4441]),

			.SO(gen[4534]),
			.S(gen[4535]),
			.SE(gen[4536]),

			.SELF(gen[4440]),
			.cell_state(gen[4440])
		); 

/******************* CELL 4441 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4441 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4345]),
			.N(gen[4346]),
			.NE(gen[4347]),

			.O(gen[4440]),
			.E(gen[4442]),

			.SO(gen[4535]),
			.S(gen[4536]),
			.SE(gen[4537]),

			.SELF(gen[4441]),
			.cell_state(gen[4441])
		); 

/******************* CELL 4442 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4442 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4346]),
			.N(gen[4347]),
			.NE(gen[4348]),

			.O(gen[4441]),
			.E(gen[4443]),

			.SO(gen[4536]),
			.S(gen[4537]),
			.SE(gen[4538]),

			.SELF(gen[4442]),
			.cell_state(gen[4442])
		); 

/******************* CELL 4443 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4443 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4347]),
			.N(gen[4348]),
			.NE(gen[4349]),

			.O(gen[4442]),
			.E(gen[4444]),

			.SO(gen[4537]),
			.S(gen[4538]),
			.SE(gen[4539]),

			.SELF(gen[4443]),
			.cell_state(gen[4443])
		); 

/******************* CELL 4444 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4444 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4348]),
			.N(gen[4349]),
			.NE(gen[4350]),

			.O(gen[4443]),
			.E(gen[4445]),

			.SO(gen[4538]),
			.S(gen[4539]),
			.SE(gen[4540]),

			.SELF(gen[4444]),
			.cell_state(gen[4444])
		); 

/******************* CELL 4445 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4445 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4349]),
			.N(gen[4350]),
			.NE(gen[4351]),

			.O(gen[4444]),
			.E(gen[4446]),

			.SO(gen[4539]),
			.S(gen[4540]),
			.SE(gen[4541]),

			.SELF(gen[4445]),
			.cell_state(gen[4445])
		); 

/******************* CELL 4446 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4446 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4350]),
			.N(gen[4351]),
			.NE(gen[4352]),

			.O(gen[4445]),
			.E(gen[4447]),

			.SO(gen[4540]),
			.S(gen[4541]),
			.SE(gen[4542]),

			.SELF(gen[4446]),
			.cell_state(gen[4446])
		); 

/******************* CELL 4447 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4447 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4351]),
			.N(gen[4352]),
			.NE(gen[4353]),

			.O(gen[4446]),
			.E(gen[4448]),

			.SO(gen[4541]),
			.S(gen[4542]),
			.SE(gen[4543]),

			.SELF(gen[4447]),
			.cell_state(gen[4447])
		); 

/******************* CELL 4448 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4448 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4352]),
			.N(gen[4353]),
			.NE(gen[4354]),

			.O(gen[4447]),
			.E(gen[4449]),

			.SO(gen[4542]),
			.S(gen[4543]),
			.SE(gen[4544]),

			.SELF(gen[4448]),
			.cell_state(gen[4448])
		); 

/******************* CELL 4449 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4449 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4353]),
			.N(gen[4354]),
			.NE(gen[4355]),

			.O(gen[4448]),
			.E(gen[4450]),

			.SO(gen[4543]),
			.S(gen[4544]),
			.SE(gen[4545]),

			.SELF(gen[4449]),
			.cell_state(gen[4449])
		); 

/******************* CELL 4450 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4450 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4354]),
			.N(gen[4355]),
			.NE(gen[4356]),

			.O(gen[4449]),
			.E(gen[4451]),

			.SO(gen[4544]),
			.S(gen[4545]),
			.SE(gen[4546]),

			.SELF(gen[4450]),
			.cell_state(gen[4450])
		); 

/******************* CELL 4451 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4451 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4355]),
			.N(gen[4356]),
			.NE(gen[4357]),

			.O(gen[4450]),
			.E(gen[4452]),

			.SO(gen[4545]),
			.S(gen[4546]),
			.SE(gen[4547]),

			.SELF(gen[4451]),
			.cell_state(gen[4451])
		); 

/******************* CELL 4452 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4452 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4356]),
			.N(gen[4357]),
			.NE(gen[4358]),

			.O(gen[4451]),
			.E(gen[4453]),

			.SO(gen[4546]),
			.S(gen[4547]),
			.SE(gen[4548]),

			.SELF(gen[4452]),
			.cell_state(gen[4452])
		); 

/******************* CELL 4453 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4453 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4357]),
			.N(gen[4358]),
			.NE(gen[4359]),

			.O(gen[4452]),
			.E(gen[4454]),

			.SO(gen[4547]),
			.S(gen[4548]),
			.SE(gen[4549]),

			.SELF(gen[4453]),
			.cell_state(gen[4453])
		); 

/******************* CELL 4454 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4454 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4358]),
			.N(gen[4359]),
			.NE(gen[4360]),

			.O(gen[4453]),
			.E(gen[4455]),

			.SO(gen[4548]),
			.S(gen[4549]),
			.SE(gen[4550]),

			.SELF(gen[4454]),
			.cell_state(gen[4454])
		); 

/******************* CELL 4455 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4455 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4359]),
			.N(gen[4360]),
			.NE(gen[4361]),

			.O(gen[4454]),
			.E(gen[4456]),

			.SO(gen[4549]),
			.S(gen[4550]),
			.SE(gen[4551]),

			.SELF(gen[4455]),
			.cell_state(gen[4455])
		); 

/******************* CELL 4456 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4456 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4360]),
			.N(gen[4361]),
			.NE(gen[4362]),

			.O(gen[4455]),
			.E(gen[4457]),

			.SO(gen[4550]),
			.S(gen[4551]),
			.SE(gen[4552]),

			.SELF(gen[4456]),
			.cell_state(gen[4456])
		); 

/******************* CELL 4457 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4457 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4361]),
			.N(gen[4362]),
			.NE(gen[4363]),

			.O(gen[4456]),
			.E(gen[4458]),

			.SO(gen[4551]),
			.S(gen[4552]),
			.SE(gen[4553]),

			.SELF(gen[4457]),
			.cell_state(gen[4457])
		); 

/******************* CELL 4458 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4458 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4362]),
			.N(gen[4363]),
			.NE(gen[4364]),

			.O(gen[4457]),
			.E(gen[4459]),

			.SO(gen[4552]),
			.S(gen[4553]),
			.SE(gen[4554]),

			.SELF(gen[4458]),
			.cell_state(gen[4458])
		); 

/******************* CELL 4459 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4459 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4363]),
			.N(gen[4364]),
			.NE(gen[4365]),

			.O(gen[4458]),
			.E(gen[4460]),

			.SO(gen[4553]),
			.S(gen[4554]),
			.SE(gen[4555]),

			.SELF(gen[4459]),
			.cell_state(gen[4459])
		); 

/******************* CELL 4460 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4460 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4364]),
			.N(gen[4365]),
			.NE(gen[4366]),

			.O(gen[4459]),
			.E(gen[4461]),

			.SO(gen[4554]),
			.S(gen[4555]),
			.SE(gen[4556]),

			.SELF(gen[4460]),
			.cell_state(gen[4460])
		); 

/******************* CELL 4461 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4461 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4365]),
			.N(gen[4366]),
			.NE(gen[4367]),

			.O(gen[4460]),
			.E(gen[4462]),

			.SO(gen[4555]),
			.S(gen[4556]),
			.SE(gen[4557]),

			.SELF(gen[4461]),
			.cell_state(gen[4461])
		); 

/******************* CELL 4462 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4462 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4366]),
			.N(gen[4367]),
			.NE(gen[4368]),

			.O(gen[4461]),
			.E(gen[4463]),

			.SO(gen[4556]),
			.S(gen[4557]),
			.SE(gen[4558]),

			.SELF(gen[4462]),
			.cell_state(gen[4462])
		); 

/******************* CELL 4463 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4463 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4367]),
			.N(gen[4368]),
			.NE(gen[4369]),

			.O(gen[4462]),
			.E(gen[4464]),

			.SO(gen[4557]),
			.S(gen[4558]),
			.SE(gen[4559]),

			.SELF(gen[4463]),
			.cell_state(gen[4463])
		); 

/******************* CELL 4464 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4464 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4368]),
			.N(gen[4369]),
			.NE(gen[4368]),

			.O(gen[4463]),
			.E(gen[4463]),

			.SO(gen[4558]),
			.S(gen[4559]),
			.SE(gen[4558]),

			.SELF(gen[4464]),
			.cell_state(gen[4464])
		); 

/******************* CELL 4465 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4465 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4371]),
			.N(gen[4370]),
			.NE(gen[4371]),

			.O(gen[4466]),
			.E(gen[4466]),

			.SO(gen[4561]),
			.S(gen[4560]),
			.SE(gen[4561]),

			.SELF(gen[4465]),
			.cell_state(gen[4465])
		); 

/******************* CELL 4466 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4466 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4370]),
			.N(gen[4371]),
			.NE(gen[4372]),

			.O(gen[4465]),
			.E(gen[4467]),

			.SO(gen[4560]),
			.S(gen[4561]),
			.SE(gen[4562]),

			.SELF(gen[4466]),
			.cell_state(gen[4466])
		); 

/******************* CELL 4467 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4467 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4371]),
			.N(gen[4372]),
			.NE(gen[4373]),

			.O(gen[4466]),
			.E(gen[4468]),

			.SO(gen[4561]),
			.S(gen[4562]),
			.SE(gen[4563]),

			.SELF(gen[4467]),
			.cell_state(gen[4467])
		); 

/******************* CELL 4468 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4468 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4372]),
			.N(gen[4373]),
			.NE(gen[4374]),

			.O(gen[4467]),
			.E(gen[4469]),

			.SO(gen[4562]),
			.S(gen[4563]),
			.SE(gen[4564]),

			.SELF(gen[4468]),
			.cell_state(gen[4468])
		); 

/******************* CELL 4469 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4469 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4373]),
			.N(gen[4374]),
			.NE(gen[4375]),

			.O(gen[4468]),
			.E(gen[4470]),

			.SO(gen[4563]),
			.S(gen[4564]),
			.SE(gen[4565]),

			.SELF(gen[4469]),
			.cell_state(gen[4469])
		); 

/******************* CELL 4470 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4470 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4374]),
			.N(gen[4375]),
			.NE(gen[4376]),

			.O(gen[4469]),
			.E(gen[4471]),

			.SO(gen[4564]),
			.S(gen[4565]),
			.SE(gen[4566]),

			.SELF(gen[4470]),
			.cell_state(gen[4470])
		); 

/******************* CELL 4471 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4471 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4375]),
			.N(gen[4376]),
			.NE(gen[4377]),

			.O(gen[4470]),
			.E(gen[4472]),

			.SO(gen[4565]),
			.S(gen[4566]),
			.SE(gen[4567]),

			.SELF(gen[4471]),
			.cell_state(gen[4471])
		); 

/******************* CELL 4472 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4472 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4376]),
			.N(gen[4377]),
			.NE(gen[4378]),

			.O(gen[4471]),
			.E(gen[4473]),

			.SO(gen[4566]),
			.S(gen[4567]),
			.SE(gen[4568]),

			.SELF(gen[4472]),
			.cell_state(gen[4472])
		); 

/******************* CELL 4473 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4473 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4377]),
			.N(gen[4378]),
			.NE(gen[4379]),

			.O(gen[4472]),
			.E(gen[4474]),

			.SO(gen[4567]),
			.S(gen[4568]),
			.SE(gen[4569]),

			.SELF(gen[4473]),
			.cell_state(gen[4473])
		); 

/******************* CELL 4474 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4474 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4378]),
			.N(gen[4379]),
			.NE(gen[4380]),

			.O(gen[4473]),
			.E(gen[4475]),

			.SO(gen[4568]),
			.S(gen[4569]),
			.SE(gen[4570]),

			.SELF(gen[4474]),
			.cell_state(gen[4474])
		); 

/******************* CELL 4475 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4475 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4379]),
			.N(gen[4380]),
			.NE(gen[4381]),

			.O(gen[4474]),
			.E(gen[4476]),

			.SO(gen[4569]),
			.S(gen[4570]),
			.SE(gen[4571]),

			.SELF(gen[4475]),
			.cell_state(gen[4475])
		); 

/******************* CELL 4476 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4476 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4380]),
			.N(gen[4381]),
			.NE(gen[4382]),

			.O(gen[4475]),
			.E(gen[4477]),

			.SO(gen[4570]),
			.S(gen[4571]),
			.SE(gen[4572]),

			.SELF(gen[4476]),
			.cell_state(gen[4476])
		); 

/******************* CELL 4477 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4477 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4381]),
			.N(gen[4382]),
			.NE(gen[4383]),

			.O(gen[4476]),
			.E(gen[4478]),

			.SO(gen[4571]),
			.S(gen[4572]),
			.SE(gen[4573]),

			.SELF(gen[4477]),
			.cell_state(gen[4477])
		); 

/******************* CELL 4478 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4478 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4382]),
			.N(gen[4383]),
			.NE(gen[4384]),

			.O(gen[4477]),
			.E(gen[4479]),

			.SO(gen[4572]),
			.S(gen[4573]),
			.SE(gen[4574]),

			.SELF(gen[4478]),
			.cell_state(gen[4478])
		); 

/******************* CELL 4479 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4479 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4383]),
			.N(gen[4384]),
			.NE(gen[4385]),

			.O(gen[4478]),
			.E(gen[4480]),

			.SO(gen[4573]),
			.S(gen[4574]),
			.SE(gen[4575]),

			.SELF(gen[4479]),
			.cell_state(gen[4479])
		); 

/******************* CELL 4480 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4480 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4384]),
			.N(gen[4385]),
			.NE(gen[4386]),

			.O(gen[4479]),
			.E(gen[4481]),

			.SO(gen[4574]),
			.S(gen[4575]),
			.SE(gen[4576]),

			.SELF(gen[4480]),
			.cell_state(gen[4480])
		); 

/******************* CELL 4481 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4481 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4385]),
			.N(gen[4386]),
			.NE(gen[4387]),

			.O(gen[4480]),
			.E(gen[4482]),

			.SO(gen[4575]),
			.S(gen[4576]),
			.SE(gen[4577]),

			.SELF(gen[4481]),
			.cell_state(gen[4481])
		); 

/******************* CELL 4482 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4482 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4386]),
			.N(gen[4387]),
			.NE(gen[4388]),

			.O(gen[4481]),
			.E(gen[4483]),

			.SO(gen[4576]),
			.S(gen[4577]),
			.SE(gen[4578]),

			.SELF(gen[4482]),
			.cell_state(gen[4482])
		); 

/******************* CELL 4483 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4483 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4387]),
			.N(gen[4388]),
			.NE(gen[4389]),

			.O(gen[4482]),
			.E(gen[4484]),

			.SO(gen[4577]),
			.S(gen[4578]),
			.SE(gen[4579]),

			.SELF(gen[4483]),
			.cell_state(gen[4483])
		); 

/******************* CELL 4484 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4484 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4388]),
			.N(gen[4389]),
			.NE(gen[4390]),

			.O(gen[4483]),
			.E(gen[4485]),

			.SO(gen[4578]),
			.S(gen[4579]),
			.SE(gen[4580]),

			.SELF(gen[4484]),
			.cell_state(gen[4484])
		); 

/******************* CELL 4485 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4485 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4389]),
			.N(gen[4390]),
			.NE(gen[4391]),

			.O(gen[4484]),
			.E(gen[4486]),

			.SO(gen[4579]),
			.S(gen[4580]),
			.SE(gen[4581]),

			.SELF(gen[4485]),
			.cell_state(gen[4485])
		); 

/******************* CELL 4486 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4486 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4390]),
			.N(gen[4391]),
			.NE(gen[4392]),

			.O(gen[4485]),
			.E(gen[4487]),

			.SO(gen[4580]),
			.S(gen[4581]),
			.SE(gen[4582]),

			.SELF(gen[4486]),
			.cell_state(gen[4486])
		); 

/******************* CELL 4487 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4487 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4391]),
			.N(gen[4392]),
			.NE(gen[4393]),

			.O(gen[4486]),
			.E(gen[4488]),

			.SO(gen[4581]),
			.S(gen[4582]),
			.SE(gen[4583]),

			.SELF(gen[4487]),
			.cell_state(gen[4487])
		); 

/******************* CELL 4488 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4488 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4392]),
			.N(gen[4393]),
			.NE(gen[4394]),

			.O(gen[4487]),
			.E(gen[4489]),

			.SO(gen[4582]),
			.S(gen[4583]),
			.SE(gen[4584]),

			.SELF(gen[4488]),
			.cell_state(gen[4488])
		); 

/******************* CELL 4489 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4489 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4393]),
			.N(gen[4394]),
			.NE(gen[4395]),

			.O(gen[4488]),
			.E(gen[4490]),

			.SO(gen[4583]),
			.S(gen[4584]),
			.SE(gen[4585]),

			.SELF(gen[4489]),
			.cell_state(gen[4489])
		); 

/******************* CELL 4490 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4490 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4394]),
			.N(gen[4395]),
			.NE(gen[4396]),

			.O(gen[4489]),
			.E(gen[4491]),

			.SO(gen[4584]),
			.S(gen[4585]),
			.SE(gen[4586]),

			.SELF(gen[4490]),
			.cell_state(gen[4490])
		); 

/******************* CELL 4491 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4491 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4395]),
			.N(gen[4396]),
			.NE(gen[4397]),

			.O(gen[4490]),
			.E(gen[4492]),

			.SO(gen[4585]),
			.S(gen[4586]),
			.SE(gen[4587]),

			.SELF(gen[4491]),
			.cell_state(gen[4491])
		); 

/******************* CELL 4492 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4492 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4396]),
			.N(gen[4397]),
			.NE(gen[4398]),

			.O(gen[4491]),
			.E(gen[4493]),

			.SO(gen[4586]),
			.S(gen[4587]),
			.SE(gen[4588]),

			.SELF(gen[4492]),
			.cell_state(gen[4492])
		); 

/******************* CELL 4493 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4493 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4397]),
			.N(gen[4398]),
			.NE(gen[4399]),

			.O(gen[4492]),
			.E(gen[4494]),

			.SO(gen[4587]),
			.S(gen[4588]),
			.SE(gen[4589]),

			.SELF(gen[4493]),
			.cell_state(gen[4493])
		); 

/******************* CELL 4494 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4494 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4398]),
			.N(gen[4399]),
			.NE(gen[4400]),

			.O(gen[4493]),
			.E(gen[4495]),

			.SO(gen[4588]),
			.S(gen[4589]),
			.SE(gen[4590]),

			.SELF(gen[4494]),
			.cell_state(gen[4494])
		); 

/******************* CELL 4495 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4495 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4399]),
			.N(gen[4400]),
			.NE(gen[4401]),

			.O(gen[4494]),
			.E(gen[4496]),

			.SO(gen[4589]),
			.S(gen[4590]),
			.SE(gen[4591]),

			.SELF(gen[4495]),
			.cell_state(gen[4495])
		); 

/******************* CELL 4496 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4496 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4400]),
			.N(gen[4401]),
			.NE(gen[4402]),

			.O(gen[4495]),
			.E(gen[4497]),

			.SO(gen[4590]),
			.S(gen[4591]),
			.SE(gen[4592]),

			.SELF(gen[4496]),
			.cell_state(gen[4496])
		); 

/******************* CELL 4497 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4497 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4401]),
			.N(gen[4402]),
			.NE(gen[4403]),

			.O(gen[4496]),
			.E(gen[4498]),

			.SO(gen[4591]),
			.S(gen[4592]),
			.SE(gen[4593]),

			.SELF(gen[4497]),
			.cell_state(gen[4497])
		); 

/******************* CELL 4498 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4498 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4402]),
			.N(gen[4403]),
			.NE(gen[4404]),

			.O(gen[4497]),
			.E(gen[4499]),

			.SO(gen[4592]),
			.S(gen[4593]),
			.SE(gen[4594]),

			.SELF(gen[4498]),
			.cell_state(gen[4498])
		); 

/******************* CELL 4499 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4499 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4403]),
			.N(gen[4404]),
			.NE(gen[4405]),

			.O(gen[4498]),
			.E(gen[4500]),

			.SO(gen[4593]),
			.S(gen[4594]),
			.SE(gen[4595]),

			.SELF(gen[4499]),
			.cell_state(gen[4499])
		); 

/******************* CELL 4500 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4500 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4404]),
			.N(gen[4405]),
			.NE(gen[4406]),

			.O(gen[4499]),
			.E(gen[4501]),

			.SO(gen[4594]),
			.S(gen[4595]),
			.SE(gen[4596]),

			.SELF(gen[4500]),
			.cell_state(gen[4500])
		); 

/******************* CELL 4501 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4501 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4405]),
			.N(gen[4406]),
			.NE(gen[4407]),

			.O(gen[4500]),
			.E(gen[4502]),

			.SO(gen[4595]),
			.S(gen[4596]),
			.SE(gen[4597]),

			.SELF(gen[4501]),
			.cell_state(gen[4501])
		); 

/******************* CELL 4502 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4502 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4406]),
			.N(gen[4407]),
			.NE(gen[4408]),

			.O(gen[4501]),
			.E(gen[4503]),

			.SO(gen[4596]),
			.S(gen[4597]),
			.SE(gen[4598]),

			.SELF(gen[4502]),
			.cell_state(gen[4502])
		); 

/******************* CELL 4503 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4503 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4407]),
			.N(gen[4408]),
			.NE(gen[4409]),

			.O(gen[4502]),
			.E(gen[4504]),

			.SO(gen[4597]),
			.S(gen[4598]),
			.SE(gen[4599]),

			.SELF(gen[4503]),
			.cell_state(gen[4503])
		); 

/******************* CELL 4504 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4504 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4408]),
			.N(gen[4409]),
			.NE(gen[4410]),

			.O(gen[4503]),
			.E(gen[4505]),

			.SO(gen[4598]),
			.S(gen[4599]),
			.SE(gen[4600]),

			.SELF(gen[4504]),
			.cell_state(gen[4504])
		); 

/******************* CELL 4505 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4505 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4409]),
			.N(gen[4410]),
			.NE(gen[4411]),

			.O(gen[4504]),
			.E(gen[4506]),

			.SO(gen[4599]),
			.S(gen[4600]),
			.SE(gen[4601]),

			.SELF(gen[4505]),
			.cell_state(gen[4505])
		); 

/******************* CELL 4506 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4506 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4410]),
			.N(gen[4411]),
			.NE(gen[4412]),

			.O(gen[4505]),
			.E(gen[4507]),

			.SO(gen[4600]),
			.S(gen[4601]),
			.SE(gen[4602]),

			.SELF(gen[4506]),
			.cell_state(gen[4506])
		); 

/******************* CELL 4507 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4507 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4411]),
			.N(gen[4412]),
			.NE(gen[4413]),

			.O(gen[4506]),
			.E(gen[4508]),

			.SO(gen[4601]),
			.S(gen[4602]),
			.SE(gen[4603]),

			.SELF(gen[4507]),
			.cell_state(gen[4507])
		); 

/******************* CELL 4508 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4508 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4412]),
			.N(gen[4413]),
			.NE(gen[4414]),

			.O(gen[4507]),
			.E(gen[4509]),

			.SO(gen[4602]),
			.S(gen[4603]),
			.SE(gen[4604]),

			.SELF(gen[4508]),
			.cell_state(gen[4508])
		); 

/******************* CELL 4509 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4509 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4413]),
			.N(gen[4414]),
			.NE(gen[4415]),

			.O(gen[4508]),
			.E(gen[4510]),

			.SO(gen[4603]),
			.S(gen[4604]),
			.SE(gen[4605]),

			.SELF(gen[4509]),
			.cell_state(gen[4509])
		); 

/******************* CELL 4510 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4510 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4414]),
			.N(gen[4415]),
			.NE(gen[4416]),

			.O(gen[4509]),
			.E(gen[4511]),

			.SO(gen[4604]),
			.S(gen[4605]),
			.SE(gen[4606]),

			.SELF(gen[4510]),
			.cell_state(gen[4510])
		); 

/******************* CELL 4511 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4511 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4415]),
			.N(gen[4416]),
			.NE(gen[4417]),

			.O(gen[4510]),
			.E(gen[4512]),

			.SO(gen[4605]),
			.S(gen[4606]),
			.SE(gen[4607]),

			.SELF(gen[4511]),
			.cell_state(gen[4511])
		); 

/******************* CELL 4512 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4512 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4416]),
			.N(gen[4417]),
			.NE(gen[4418]),

			.O(gen[4511]),
			.E(gen[4513]),

			.SO(gen[4606]),
			.S(gen[4607]),
			.SE(gen[4608]),

			.SELF(gen[4512]),
			.cell_state(gen[4512])
		); 

/******************* CELL 4513 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4513 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4417]),
			.N(gen[4418]),
			.NE(gen[4419]),

			.O(gen[4512]),
			.E(gen[4514]),

			.SO(gen[4607]),
			.S(gen[4608]),
			.SE(gen[4609]),

			.SELF(gen[4513]),
			.cell_state(gen[4513])
		); 

/******************* CELL 4514 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4514 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4418]),
			.N(gen[4419]),
			.NE(gen[4420]),

			.O(gen[4513]),
			.E(gen[4515]),

			.SO(gen[4608]),
			.S(gen[4609]),
			.SE(gen[4610]),

			.SELF(gen[4514]),
			.cell_state(gen[4514])
		); 

/******************* CELL 4515 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4515 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4419]),
			.N(gen[4420]),
			.NE(gen[4421]),

			.O(gen[4514]),
			.E(gen[4516]),

			.SO(gen[4609]),
			.S(gen[4610]),
			.SE(gen[4611]),

			.SELF(gen[4515]),
			.cell_state(gen[4515])
		); 

/******************* CELL 4516 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4516 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4420]),
			.N(gen[4421]),
			.NE(gen[4422]),

			.O(gen[4515]),
			.E(gen[4517]),

			.SO(gen[4610]),
			.S(gen[4611]),
			.SE(gen[4612]),

			.SELF(gen[4516]),
			.cell_state(gen[4516])
		); 

/******************* CELL 4517 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4517 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4421]),
			.N(gen[4422]),
			.NE(gen[4423]),

			.O(gen[4516]),
			.E(gen[4518]),

			.SO(gen[4611]),
			.S(gen[4612]),
			.SE(gen[4613]),

			.SELF(gen[4517]),
			.cell_state(gen[4517])
		); 

/******************* CELL 4518 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4518 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4422]),
			.N(gen[4423]),
			.NE(gen[4424]),

			.O(gen[4517]),
			.E(gen[4519]),

			.SO(gen[4612]),
			.S(gen[4613]),
			.SE(gen[4614]),

			.SELF(gen[4518]),
			.cell_state(gen[4518])
		); 

/******************* CELL 4519 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4519 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4423]),
			.N(gen[4424]),
			.NE(gen[4425]),

			.O(gen[4518]),
			.E(gen[4520]),

			.SO(gen[4613]),
			.S(gen[4614]),
			.SE(gen[4615]),

			.SELF(gen[4519]),
			.cell_state(gen[4519])
		); 

/******************* CELL 4520 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4520 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4424]),
			.N(gen[4425]),
			.NE(gen[4426]),

			.O(gen[4519]),
			.E(gen[4521]),

			.SO(gen[4614]),
			.S(gen[4615]),
			.SE(gen[4616]),

			.SELF(gen[4520]),
			.cell_state(gen[4520])
		); 

/******************* CELL 4521 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4521 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4425]),
			.N(gen[4426]),
			.NE(gen[4427]),

			.O(gen[4520]),
			.E(gen[4522]),

			.SO(gen[4615]),
			.S(gen[4616]),
			.SE(gen[4617]),

			.SELF(gen[4521]),
			.cell_state(gen[4521])
		); 

/******************* CELL 4522 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4522 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4426]),
			.N(gen[4427]),
			.NE(gen[4428]),

			.O(gen[4521]),
			.E(gen[4523]),

			.SO(gen[4616]),
			.S(gen[4617]),
			.SE(gen[4618]),

			.SELF(gen[4522]),
			.cell_state(gen[4522])
		); 

/******************* CELL 4523 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4523 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4427]),
			.N(gen[4428]),
			.NE(gen[4429]),

			.O(gen[4522]),
			.E(gen[4524]),

			.SO(gen[4617]),
			.S(gen[4618]),
			.SE(gen[4619]),

			.SELF(gen[4523]),
			.cell_state(gen[4523])
		); 

/******************* CELL 4524 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4524 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4428]),
			.N(gen[4429]),
			.NE(gen[4430]),

			.O(gen[4523]),
			.E(gen[4525]),

			.SO(gen[4618]),
			.S(gen[4619]),
			.SE(gen[4620]),

			.SELF(gen[4524]),
			.cell_state(gen[4524])
		); 

/******************* CELL 4525 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4525 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4429]),
			.N(gen[4430]),
			.NE(gen[4431]),

			.O(gen[4524]),
			.E(gen[4526]),

			.SO(gen[4619]),
			.S(gen[4620]),
			.SE(gen[4621]),

			.SELF(gen[4525]),
			.cell_state(gen[4525])
		); 

/******************* CELL 4526 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4526 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4430]),
			.N(gen[4431]),
			.NE(gen[4432]),

			.O(gen[4525]),
			.E(gen[4527]),

			.SO(gen[4620]),
			.S(gen[4621]),
			.SE(gen[4622]),

			.SELF(gen[4526]),
			.cell_state(gen[4526])
		); 

/******************* CELL 4527 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4527 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4431]),
			.N(gen[4432]),
			.NE(gen[4433]),

			.O(gen[4526]),
			.E(gen[4528]),

			.SO(gen[4621]),
			.S(gen[4622]),
			.SE(gen[4623]),

			.SELF(gen[4527]),
			.cell_state(gen[4527])
		); 

/******************* CELL 4528 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4528 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4432]),
			.N(gen[4433]),
			.NE(gen[4434]),

			.O(gen[4527]),
			.E(gen[4529]),

			.SO(gen[4622]),
			.S(gen[4623]),
			.SE(gen[4624]),

			.SELF(gen[4528]),
			.cell_state(gen[4528])
		); 

/******************* CELL 4529 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4529 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4433]),
			.N(gen[4434]),
			.NE(gen[4435]),

			.O(gen[4528]),
			.E(gen[4530]),

			.SO(gen[4623]),
			.S(gen[4624]),
			.SE(gen[4625]),

			.SELF(gen[4529]),
			.cell_state(gen[4529])
		); 

/******************* CELL 4530 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4530 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4434]),
			.N(gen[4435]),
			.NE(gen[4436]),

			.O(gen[4529]),
			.E(gen[4531]),

			.SO(gen[4624]),
			.S(gen[4625]),
			.SE(gen[4626]),

			.SELF(gen[4530]),
			.cell_state(gen[4530])
		); 

/******************* CELL 4531 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4531 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4435]),
			.N(gen[4436]),
			.NE(gen[4437]),

			.O(gen[4530]),
			.E(gen[4532]),

			.SO(gen[4625]),
			.S(gen[4626]),
			.SE(gen[4627]),

			.SELF(gen[4531]),
			.cell_state(gen[4531])
		); 

/******************* CELL 4532 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4532 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4436]),
			.N(gen[4437]),
			.NE(gen[4438]),

			.O(gen[4531]),
			.E(gen[4533]),

			.SO(gen[4626]),
			.S(gen[4627]),
			.SE(gen[4628]),

			.SELF(gen[4532]),
			.cell_state(gen[4532])
		); 

/******************* CELL 4533 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4533 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4437]),
			.N(gen[4438]),
			.NE(gen[4439]),

			.O(gen[4532]),
			.E(gen[4534]),

			.SO(gen[4627]),
			.S(gen[4628]),
			.SE(gen[4629]),

			.SELF(gen[4533]),
			.cell_state(gen[4533])
		); 

/******************* CELL 4534 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4534 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4438]),
			.N(gen[4439]),
			.NE(gen[4440]),

			.O(gen[4533]),
			.E(gen[4535]),

			.SO(gen[4628]),
			.S(gen[4629]),
			.SE(gen[4630]),

			.SELF(gen[4534]),
			.cell_state(gen[4534])
		); 

/******************* CELL 4535 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4535 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4439]),
			.N(gen[4440]),
			.NE(gen[4441]),

			.O(gen[4534]),
			.E(gen[4536]),

			.SO(gen[4629]),
			.S(gen[4630]),
			.SE(gen[4631]),

			.SELF(gen[4535]),
			.cell_state(gen[4535])
		); 

/******************* CELL 4536 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4536 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4440]),
			.N(gen[4441]),
			.NE(gen[4442]),

			.O(gen[4535]),
			.E(gen[4537]),

			.SO(gen[4630]),
			.S(gen[4631]),
			.SE(gen[4632]),

			.SELF(gen[4536]),
			.cell_state(gen[4536])
		); 

/******************* CELL 4537 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4537 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4441]),
			.N(gen[4442]),
			.NE(gen[4443]),

			.O(gen[4536]),
			.E(gen[4538]),

			.SO(gen[4631]),
			.S(gen[4632]),
			.SE(gen[4633]),

			.SELF(gen[4537]),
			.cell_state(gen[4537])
		); 

/******************* CELL 4538 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4538 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4442]),
			.N(gen[4443]),
			.NE(gen[4444]),

			.O(gen[4537]),
			.E(gen[4539]),

			.SO(gen[4632]),
			.S(gen[4633]),
			.SE(gen[4634]),

			.SELF(gen[4538]),
			.cell_state(gen[4538])
		); 

/******************* CELL 4539 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4539 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4443]),
			.N(gen[4444]),
			.NE(gen[4445]),

			.O(gen[4538]),
			.E(gen[4540]),

			.SO(gen[4633]),
			.S(gen[4634]),
			.SE(gen[4635]),

			.SELF(gen[4539]),
			.cell_state(gen[4539])
		); 

/******************* CELL 4540 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4540 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4444]),
			.N(gen[4445]),
			.NE(gen[4446]),

			.O(gen[4539]),
			.E(gen[4541]),

			.SO(gen[4634]),
			.S(gen[4635]),
			.SE(gen[4636]),

			.SELF(gen[4540]),
			.cell_state(gen[4540])
		); 

/******************* CELL 4541 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4541 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4445]),
			.N(gen[4446]),
			.NE(gen[4447]),

			.O(gen[4540]),
			.E(gen[4542]),

			.SO(gen[4635]),
			.S(gen[4636]),
			.SE(gen[4637]),

			.SELF(gen[4541]),
			.cell_state(gen[4541])
		); 

/******************* CELL 4542 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4542 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4446]),
			.N(gen[4447]),
			.NE(gen[4448]),

			.O(gen[4541]),
			.E(gen[4543]),

			.SO(gen[4636]),
			.S(gen[4637]),
			.SE(gen[4638]),

			.SELF(gen[4542]),
			.cell_state(gen[4542])
		); 

/******************* CELL 4543 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4543 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4447]),
			.N(gen[4448]),
			.NE(gen[4449]),

			.O(gen[4542]),
			.E(gen[4544]),

			.SO(gen[4637]),
			.S(gen[4638]),
			.SE(gen[4639]),

			.SELF(gen[4543]),
			.cell_state(gen[4543])
		); 

/******************* CELL 4544 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4544 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4448]),
			.N(gen[4449]),
			.NE(gen[4450]),

			.O(gen[4543]),
			.E(gen[4545]),

			.SO(gen[4638]),
			.S(gen[4639]),
			.SE(gen[4640]),

			.SELF(gen[4544]),
			.cell_state(gen[4544])
		); 

/******************* CELL 4545 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4545 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4449]),
			.N(gen[4450]),
			.NE(gen[4451]),

			.O(gen[4544]),
			.E(gen[4546]),

			.SO(gen[4639]),
			.S(gen[4640]),
			.SE(gen[4641]),

			.SELF(gen[4545]),
			.cell_state(gen[4545])
		); 

/******************* CELL 4546 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4546 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4450]),
			.N(gen[4451]),
			.NE(gen[4452]),

			.O(gen[4545]),
			.E(gen[4547]),

			.SO(gen[4640]),
			.S(gen[4641]),
			.SE(gen[4642]),

			.SELF(gen[4546]),
			.cell_state(gen[4546])
		); 

/******************* CELL 4547 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4547 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4451]),
			.N(gen[4452]),
			.NE(gen[4453]),

			.O(gen[4546]),
			.E(gen[4548]),

			.SO(gen[4641]),
			.S(gen[4642]),
			.SE(gen[4643]),

			.SELF(gen[4547]),
			.cell_state(gen[4547])
		); 

/******************* CELL 4548 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4548 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4452]),
			.N(gen[4453]),
			.NE(gen[4454]),

			.O(gen[4547]),
			.E(gen[4549]),

			.SO(gen[4642]),
			.S(gen[4643]),
			.SE(gen[4644]),

			.SELF(gen[4548]),
			.cell_state(gen[4548])
		); 

/******************* CELL 4549 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4549 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4453]),
			.N(gen[4454]),
			.NE(gen[4455]),

			.O(gen[4548]),
			.E(gen[4550]),

			.SO(gen[4643]),
			.S(gen[4644]),
			.SE(gen[4645]),

			.SELF(gen[4549]),
			.cell_state(gen[4549])
		); 

/******************* CELL 4550 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4550 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4454]),
			.N(gen[4455]),
			.NE(gen[4456]),

			.O(gen[4549]),
			.E(gen[4551]),

			.SO(gen[4644]),
			.S(gen[4645]),
			.SE(gen[4646]),

			.SELF(gen[4550]),
			.cell_state(gen[4550])
		); 

/******************* CELL 4551 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4551 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4455]),
			.N(gen[4456]),
			.NE(gen[4457]),

			.O(gen[4550]),
			.E(gen[4552]),

			.SO(gen[4645]),
			.S(gen[4646]),
			.SE(gen[4647]),

			.SELF(gen[4551]),
			.cell_state(gen[4551])
		); 

/******************* CELL 4552 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4552 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4456]),
			.N(gen[4457]),
			.NE(gen[4458]),

			.O(gen[4551]),
			.E(gen[4553]),

			.SO(gen[4646]),
			.S(gen[4647]),
			.SE(gen[4648]),

			.SELF(gen[4552]),
			.cell_state(gen[4552])
		); 

/******************* CELL 4553 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4553 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4457]),
			.N(gen[4458]),
			.NE(gen[4459]),

			.O(gen[4552]),
			.E(gen[4554]),

			.SO(gen[4647]),
			.S(gen[4648]),
			.SE(gen[4649]),

			.SELF(gen[4553]),
			.cell_state(gen[4553])
		); 

/******************* CELL 4554 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4554 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4458]),
			.N(gen[4459]),
			.NE(gen[4460]),

			.O(gen[4553]),
			.E(gen[4555]),

			.SO(gen[4648]),
			.S(gen[4649]),
			.SE(gen[4650]),

			.SELF(gen[4554]),
			.cell_state(gen[4554])
		); 

/******************* CELL 4555 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4555 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4459]),
			.N(gen[4460]),
			.NE(gen[4461]),

			.O(gen[4554]),
			.E(gen[4556]),

			.SO(gen[4649]),
			.S(gen[4650]),
			.SE(gen[4651]),

			.SELF(gen[4555]),
			.cell_state(gen[4555])
		); 

/******************* CELL 4556 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4556 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4460]),
			.N(gen[4461]),
			.NE(gen[4462]),

			.O(gen[4555]),
			.E(gen[4557]),

			.SO(gen[4650]),
			.S(gen[4651]),
			.SE(gen[4652]),

			.SELF(gen[4556]),
			.cell_state(gen[4556])
		); 

/******************* CELL 4557 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4557 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4461]),
			.N(gen[4462]),
			.NE(gen[4463]),

			.O(gen[4556]),
			.E(gen[4558]),

			.SO(gen[4651]),
			.S(gen[4652]),
			.SE(gen[4653]),

			.SELF(gen[4557]),
			.cell_state(gen[4557])
		); 

/******************* CELL 4558 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4558 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4462]),
			.N(gen[4463]),
			.NE(gen[4464]),

			.O(gen[4557]),
			.E(gen[4559]),

			.SO(gen[4652]),
			.S(gen[4653]),
			.SE(gen[4654]),

			.SELF(gen[4558]),
			.cell_state(gen[4558])
		); 

/******************* CELL 4559 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4559 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4463]),
			.N(gen[4464]),
			.NE(gen[4463]),

			.O(gen[4558]),
			.E(gen[4558]),

			.SO(gen[4653]),
			.S(gen[4654]),
			.SE(gen[4653]),

			.SELF(gen[4559]),
			.cell_state(gen[4559])
		); 

/******************* CELL 4560 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4560 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4466]),
			.N(gen[4465]),
			.NE(gen[4466]),

			.O(gen[4561]),
			.E(gen[4561]),

			.SO(gen[4656]),
			.S(gen[4655]),
			.SE(gen[4656]),

			.SELF(gen[4560]),
			.cell_state(gen[4560])
		); 

/******************* CELL 4561 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4561 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4465]),
			.N(gen[4466]),
			.NE(gen[4467]),

			.O(gen[4560]),
			.E(gen[4562]),

			.SO(gen[4655]),
			.S(gen[4656]),
			.SE(gen[4657]),

			.SELF(gen[4561]),
			.cell_state(gen[4561])
		); 

/******************* CELL 4562 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4562 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4466]),
			.N(gen[4467]),
			.NE(gen[4468]),

			.O(gen[4561]),
			.E(gen[4563]),

			.SO(gen[4656]),
			.S(gen[4657]),
			.SE(gen[4658]),

			.SELF(gen[4562]),
			.cell_state(gen[4562])
		); 

/******************* CELL 4563 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4563 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4467]),
			.N(gen[4468]),
			.NE(gen[4469]),

			.O(gen[4562]),
			.E(gen[4564]),

			.SO(gen[4657]),
			.S(gen[4658]),
			.SE(gen[4659]),

			.SELF(gen[4563]),
			.cell_state(gen[4563])
		); 

/******************* CELL 4564 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4564 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4468]),
			.N(gen[4469]),
			.NE(gen[4470]),

			.O(gen[4563]),
			.E(gen[4565]),

			.SO(gen[4658]),
			.S(gen[4659]),
			.SE(gen[4660]),

			.SELF(gen[4564]),
			.cell_state(gen[4564])
		); 

/******************* CELL 4565 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4565 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4469]),
			.N(gen[4470]),
			.NE(gen[4471]),

			.O(gen[4564]),
			.E(gen[4566]),

			.SO(gen[4659]),
			.S(gen[4660]),
			.SE(gen[4661]),

			.SELF(gen[4565]),
			.cell_state(gen[4565])
		); 

/******************* CELL 4566 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4566 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4470]),
			.N(gen[4471]),
			.NE(gen[4472]),

			.O(gen[4565]),
			.E(gen[4567]),

			.SO(gen[4660]),
			.S(gen[4661]),
			.SE(gen[4662]),

			.SELF(gen[4566]),
			.cell_state(gen[4566])
		); 

/******************* CELL 4567 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4567 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4471]),
			.N(gen[4472]),
			.NE(gen[4473]),

			.O(gen[4566]),
			.E(gen[4568]),

			.SO(gen[4661]),
			.S(gen[4662]),
			.SE(gen[4663]),

			.SELF(gen[4567]),
			.cell_state(gen[4567])
		); 

/******************* CELL 4568 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4568 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4472]),
			.N(gen[4473]),
			.NE(gen[4474]),

			.O(gen[4567]),
			.E(gen[4569]),

			.SO(gen[4662]),
			.S(gen[4663]),
			.SE(gen[4664]),

			.SELF(gen[4568]),
			.cell_state(gen[4568])
		); 

/******************* CELL 4569 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4569 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4473]),
			.N(gen[4474]),
			.NE(gen[4475]),

			.O(gen[4568]),
			.E(gen[4570]),

			.SO(gen[4663]),
			.S(gen[4664]),
			.SE(gen[4665]),

			.SELF(gen[4569]),
			.cell_state(gen[4569])
		); 

/******************* CELL 4570 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4570 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4474]),
			.N(gen[4475]),
			.NE(gen[4476]),

			.O(gen[4569]),
			.E(gen[4571]),

			.SO(gen[4664]),
			.S(gen[4665]),
			.SE(gen[4666]),

			.SELF(gen[4570]),
			.cell_state(gen[4570])
		); 

/******************* CELL 4571 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4571 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4475]),
			.N(gen[4476]),
			.NE(gen[4477]),

			.O(gen[4570]),
			.E(gen[4572]),

			.SO(gen[4665]),
			.S(gen[4666]),
			.SE(gen[4667]),

			.SELF(gen[4571]),
			.cell_state(gen[4571])
		); 

/******************* CELL 4572 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4572 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4476]),
			.N(gen[4477]),
			.NE(gen[4478]),

			.O(gen[4571]),
			.E(gen[4573]),

			.SO(gen[4666]),
			.S(gen[4667]),
			.SE(gen[4668]),

			.SELF(gen[4572]),
			.cell_state(gen[4572])
		); 

/******************* CELL 4573 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4573 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4477]),
			.N(gen[4478]),
			.NE(gen[4479]),

			.O(gen[4572]),
			.E(gen[4574]),

			.SO(gen[4667]),
			.S(gen[4668]),
			.SE(gen[4669]),

			.SELF(gen[4573]),
			.cell_state(gen[4573])
		); 

/******************* CELL 4574 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4574 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4478]),
			.N(gen[4479]),
			.NE(gen[4480]),

			.O(gen[4573]),
			.E(gen[4575]),

			.SO(gen[4668]),
			.S(gen[4669]),
			.SE(gen[4670]),

			.SELF(gen[4574]),
			.cell_state(gen[4574])
		); 

/******************* CELL 4575 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4575 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4479]),
			.N(gen[4480]),
			.NE(gen[4481]),

			.O(gen[4574]),
			.E(gen[4576]),

			.SO(gen[4669]),
			.S(gen[4670]),
			.SE(gen[4671]),

			.SELF(gen[4575]),
			.cell_state(gen[4575])
		); 

/******************* CELL 4576 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4576 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4480]),
			.N(gen[4481]),
			.NE(gen[4482]),

			.O(gen[4575]),
			.E(gen[4577]),

			.SO(gen[4670]),
			.S(gen[4671]),
			.SE(gen[4672]),

			.SELF(gen[4576]),
			.cell_state(gen[4576])
		); 

/******************* CELL 4577 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4577 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4481]),
			.N(gen[4482]),
			.NE(gen[4483]),

			.O(gen[4576]),
			.E(gen[4578]),

			.SO(gen[4671]),
			.S(gen[4672]),
			.SE(gen[4673]),

			.SELF(gen[4577]),
			.cell_state(gen[4577])
		); 

/******************* CELL 4578 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4578 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4482]),
			.N(gen[4483]),
			.NE(gen[4484]),

			.O(gen[4577]),
			.E(gen[4579]),

			.SO(gen[4672]),
			.S(gen[4673]),
			.SE(gen[4674]),

			.SELF(gen[4578]),
			.cell_state(gen[4578])
		); 

/******************* CELL 4579 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4579 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4483]),
			.N(gen[4484]),
			.NE(gen[4485]),

			.O(gen[4578]),
			.E(gen[4580]),

			.SO(gen[4673]),
			.S(gen[4674]),
			.SE(gen[4675]),

			.SELF(gen[4579]),
			.cell_state(gen[4579])
		); 

/******************* CELL 4580 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4580 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4484]),
			.N(gen[4485]),
			.NE(gen[4486]),

			.O(gen[4579]),
			.E(gen[4581]),

			.SO(gen[4674]),
			.S(gen[4675]),
			.SE(gen[4676]),

			.SELF(gen[4580]),
			.cell_state(gen[4580])
		); 

/******************* CELL 4581 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4581 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4485]),
			.N(gen[4486]),
			.NE(gen[4487]),

			.O(gen[4580]),
			.E(gen[4582]),

			.SO(gen[4675]),
			.S(gen[4676]),
			.SE(gen[4677]),

			.SELF(gen[4581]),
			.cell_state(gen[4581])
		); 

/******************* CELL 4582 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4582 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4486]),
			.N(gen[4487]),
			.NE(gen[4488]),

			.O(gen[4581]),
			.E(gen[4583]),

			.SO(gen[4676]),
			.S(gen[4677]),
			.SE(gen[4678]),

			.SELF(gen[4582]),
			.cell_state(gen[4582])
		); 

/******************* CELL 4583 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4583 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4487]),
			.N(gen[4488]),
			.NE(gen[4489]),

			.O(gen[4582]),
			.E(gen[4584]),

			.SO(gen[4677]),
			.S(gen[4678]),
			.SE(gen[4679]),

			.SELF(gen[4583]),
			.cell_state(gen[4583])
		); 

/******************* CELL 4584 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4584 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4488]),
			.N(gen[4489]),
			.NE(gen[4490]),

			.O(gen[4583]),
			.E(gen[4585]),

			.SO(gen[4678]),
			.S(gen[4679]),
			.SE(gen[4680]),

			.SELF(gen[4584]),
			.cell_state(gen[4584])
		); 

/******************* CELL 4585 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4585 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4489]),
			.N(gen[4490]),
			.NE(gen[4491]),

			.O(gen[4584]),
			.E(gen[4586]),

			.SO(gen[4679]),
			.S(gen[4680]),
			.SE(gen[4681]),

			.SELF(gen[4585]),
			.cell_state(gen[4585])
		); 

/******************* CELL 4586 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4586 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4490]),
			.N(gen[4491]),
			.NE(gen[4492]),

			.O(gen[4585]),
			.E(gen[4587]),

			.SO(gen[4680]),
			.S(gen[4681]),
			.SE(gen[4682]),

			.SELF(gen[4586]),
			.cell_state(gen[4586])
		); 

/******************* CELL 4587 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4587 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4491]),
			.N(gen[4492]),
			.NE(gen[4493]),

			.O(gen[4586]),
			.E(gen[4588]),

			.SO(gen[4681]),
			.S(gen[4682]),
			.SE(gen[4683]),

			.SELF(gen[4587]),
			.cell_state(gen[4587])
		); 

/******************* CELL 4588 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4588 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4492]),
			.N(gen[4493]),
			.NE(gen[4494]),

			.O(gen[4587]),
			.E(gen[4589]),

			.SO(gen[4682]),
			.S(gen[4683]),
			.SE(gen[4684]),

			.SELF(gen[4588]),
			.cell_state(gen[4588])
		); 

/******************* CELL 4589 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4589 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4493]),
			.N(gen[4494]),
			.NE(gen[4495]),

			.O(gen[4588]),
			.E(gen[4590]),

			.SO(gen[4683]),
			.S(gen[4684]),
			.SE(gen[4685]),

			.SELF(gen[4589]),
			.cell_state(gen[4589])
		); 

/******************* CELL 4590 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4590 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4494]),
			.N(gen[4495]),
			.NE(gen[4496]),

			.O(gen[4589]),
			.E(gen[4591]),

			.SO(gen[4684]),
			.S(gen[4685]),
			.SE(gen[4686]),

			.SELF(gen[4590]),
			.cell_state(gen[4590])
		); 

/******************* CELL 4591 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4591 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4495]),
			.N(gen[4496]),
			.NE(gen[4497]),

			.O(gen[4590]),
			.E(gen[4592]),

			.SO(gen[4685]),
			.S(gen[4686]),
			.SE(gen[4687]),

			.SELF(gen[4591]),
			.cell_state(gen[4591])
		); 

/******************* CELL 4592 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4592 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4496]),
			.N(gen[4497]),
			.NE(gen[4498]),

			.O(gen[4591]),
			.E(gen[4593]),

			.SO(gen[4686]),
			.S(gen[4687]),
			.SE(gen[4688]),

			.SELF(gen[4592]),
			.cell_state(gen[4592])
		); 

/******************* CELL 4593 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4593 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4497]),
			.N(gen[4498]),
			.NE(gen[4499]),

			.O(gen[4592]),
			.E(gen[4594]),

			.SO(gen[4687]),
			.S(gen[4688]),
			.SE(gen[4689]),

			.SELF(gen[4593]),
			.cell_state(gen[4593])
		); 

/******************* CELL 4594 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4594 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4498]),
			.N(gen[4499]),
			.NE(gen[4500]),

			.O(gen[4593]),
			.E(gen[4595]),

			.SO(gen[4688]),
			.S(gen[4689]),
			.SE(gen[4690]),

			.SELF(gen[4594]),
			.cell_state(gen[4594])
		); 

/******************* CELL 4595 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4595 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4499]),
			.N(gen[4500]),
			.NE(gen[4501]),

			.O(gen[4594]),
			.E(gen[4596]),

			.SO(gen[4689]),
			.S(gen[4690]),
			.SE(gen[4691]),

			.SELF(gen[4595]),
			.cell_state(gen[4595])
		); 

/******************* CELL 4596 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4596 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4500]),
			.N(gen[4501]),
			.NE(gen[4502]),

			.O(gen[4595]),
			.E(gen[4597]),

			.SO(gen[4690]),
			.S(gen[4691]),
			.SE(gen[4692]),

			.SELF(gen[4596]),
			.cell_state(gen[4596])
		); 

/******************* CELL 4597 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4597 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4501]),
			.N(gen[4502]),
			.NE(gen[4503]),

			.O(gen[4596]),
			.E(gen[4598]),

			.SO(gen[4691]),
			.S(gen[4692]),
			.SE(gen[4693]),

			.SELF(gen[4597]),
			.cell_state(gen[4597])
		); 

/******************* CELL 4598 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4598 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4502]),
			.N(gen[4503]),
			.NE(gen[4504]),

			.O(gen[4597]),
			.E(gen[4599]),

			.SO(gen[4692]),
			.S(gen[4693]),
			.SE(gen[4694]),

			.SELF(gen[4598]),
			.cell_state(gen[4598])
		); 

/******************* CELL 4599 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4599 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4503]),
			.N(gen[4504]),
			.NE(gen[4505]),

			.O(gen[4598]),
			.E(gen[4600]),

			.SO(gen[4693]),
			.S(gen[4694]),
			.SE(gen[4695]),

			.SELF(gen[4599]),
			.cell_state(gen[4599])
		); 

/******************* CELL 4600 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4600 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4504]),
			.N(gen[4505]),
			.NE(gen[4506]),

			.O(gen[4599]),
			.E(gen[4601]),

			.SO(gen[4694]),
			.S(gen[4695]),
			.SE(gen[4696]),

			.SELF(gen[4600]),
			.cell_state(gen[4600])
		); 

/******************* CELL 4601 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4601 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4505]),
			.N(gen[4506]),
			.NE(gen[4507]),

			.O(gen[4600]),
			.E(gen[4602]),

			.SO(gen[4695]),
			.S(gen[4696]),
			.SE(gen[4697]),

			.SELF(gen[4601]),
			.cell_state(gen[4601])
		); 

/******************* CELL 4602 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4602 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4506]),
			.N(gen[4507]),
			.NE(gen[4508]),

			.O(gen[4601]),
			.E(gen[4603]),

			.SO(gen[4696]),
			.S(gen[4697]),
			.SE(gen[4698]),

			.SELF(gen[4602]),
			.cell_state(gen[4602])
		); 

/******************* CELL 4603 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4603 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4507]),
			.N(gen[4508]),
			.NE(gen[4509]),

			.O(gen[4602]),
			.E(gen[4604]),

			.SO(gen[4697]),
			.S(gen[4698]),
			.SE(gen[4699]),

			.SELF(gen[4603]),
			.cell_state(gen[4603])
		); 

/******************* CELL 4604 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4604 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4508]),
			.N(gen[4509]),
			.NE(gen[4510]),

			.O(gen[4603]),
			.E(gen[4605]),

			.SO(gen[4698]),
			.S(gen[4699]),
			.SE(gen[4700]),

			.SELF(gen[4604]),
			.cell_state(gen[4604])
		); 

/******************* CELL 4605 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4605 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4509]),
			.N(gen[4510]),
			.NE(gen[4511]),

			.O(gen[4604]),
			.E(gen[4606]),

			.SO(gen[4699]),
			.S(gen[4700]),
			.SE(gen[4701]),

			.SELF(gen[4605]),
			.cell_state(gen[4605])
		); 

/******************* CELL 4606 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4606 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4510]),
			.N(gen[4511]),
			.NE(gen[4512]),

			.O(gen[4605]),
			.E(gen[4607]),

			.SO(gen[4700]),
			.S(gen[4701]),
			.SE(gen[4702]),

			.SELF(gen[4606]),
			.cell_state(gen[4606])
		); 

/******************* CELL 4607 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4607 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4511]),
			.N(gen[4512]),
			.NE(gen[4513]),

			.O(gen[4606]),
			.E(gen[4608]),

			.SO(gen[4701]),
			.S(gen[4702]),
			.SE(gen[4703]),

			.SELF(gen[4607]),
			.cell_state(gen[4607])
		); 

/******************* CELL 4608 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4608 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4512]),
			.N(gen[4513]),
			.NE(gen[4514]),

			.O(gen[4607]),
			.E(gen[4609]),

			.SO(gen[4702]),
			.S(gen[4703]),
			.SE(gen[4704]),

			.SELF(gen[4608]),
			.cell_state(gen[4608])
		); 

/******************* CELL 4609 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4609 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4513]),
			.N(gen[4514]),
			.NE(gen[4515]),

			.O(gen[4608]),
			.E(gen[4610]),

			.SO(gen[4703]),
			.S(gen[4704]),
			.SE(gen[4705]),

			.SELF(gen[4609]),
			.cell_state(gen[4609])
		); 

/******************* CELL 4610 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4610 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4514]),
			.N(gen[4515]),
			.NE(gen[4516]),

			.O(gen[4609]),
			.E(gen[4611]),

			.SO(gen[4704]),
			.S(gen[4705]),
			.SE(gen[4706]),

			.SELF(gen[4610]),
			.cell_state(gen[4610])
		); 

/******************* CELL 4611 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4611 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4515]),
			.N(gen[4516]),
			.NE(gen[4517]),

			.O(gen[4610]),
			.E(gen[4612]),

			.SO(gen[4705]),
			.S(gen[4706]),
			.SE(gen[4707]),

			.SELF(gen[4611]),
			.cell_state(gen[4611])
		); 

/******************* CELL 4612 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4612 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4516]),
			.N(gen[4517]),
			.NE(gen[4518]),

			.O(gen[4611]),
			.E(gen[4613]),

			.SO(gen[4706]),
			.S(gen[4707]),
			.SE(gen[4708]),

			.SELF(gen[4612]),
			.cell_state(gen[4612])
		); 

/******************* CELL 4613 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4613 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4517]),
			.N(gen[4518]),
			.NE(gen[4519]),

			.O(gen[4612]),
			.E(gen[4614]),

			.SO(gen[4707]),
			.S(gen[4708]),
			.SE(gen[4709]),

			.SELF(gen[4613]),
			.cell_state(gen[4613])
		); 

/******************* CELL 4614 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4614 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4518]),
			.N(gen[4519]),
			.NE(gen[4520]),

			.O(gen[4613]),
			.E(gen[4615]),

			.SO(gen[4708]),
			.S(gen[4709]),
			.SE(gen[4710]),

			.SELF(gen[4614]),
			.cell_state(gen[4614])
		); 

/******************* CELL 4615 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4615 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4519]),
			.N(gen[4520]),
			.NE(gen[4521]),

			.O(gen[4614]),
			.E(gen[4616]),

			.SO(gen[4709]),
			.S(gen[4710]),
			.SE(gen[4711]),

			.SELF(gen[4615]),
			.cell_state(gen[4615])
		); 

/******************* CELL 4616 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4616 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4520]),
			.N(gen[4521]),
			.NE(gen[4522]),

			.O(gen[4615]),
			.E(gen[4617]),

			.SO(gen[4710]),
			.S(gen[4711]),
			.SE(gen[4712]),

			.SELF(gen[4616]),
			.cell_state(gen[4616])
		); 

/******************* CELL 4617 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4617 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4521]),
			.N(gen[4522]),
			.NE(gen[4523]),

			.O(gen[4616]),
			.E(gen[4618]),

			.SO(gen[4711]),
			.S(gen[4712]),
			.SE(gen[4713]),

			.SELF(gen[4617]),
			.cell_state(gen[4617])
		); 

/******************* CELL 4618 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4618 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4522]),
			.N(gen[4523]),
			.NE(gen[4524]),

			.O(gen[4617]),
			.E(gen[4619]),

			.SO(gen[4712]),
			.S(gen[4713]),
			.SE(gen[4714]),

			.SELF(gen[4618]),
			.cell_state(gen[4618])
		); 

/******************* CELL 4619 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4619 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4523]),
			.N(gen[4524]),
			.NE(gen[4525]),

			.O(gen[4618]),
			.E(gen[4620]),

			.SO(gen[4713]),
			.S(gen[4714]),
			.SE(gen[4715]),

			.SELF(gen[4619]),
			.cell_state(gen[4619])
		); 

/******************* CELL 4620 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4620 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4524]),
			.N(gen[4525]),
			.NE(gen[4526]),

			.O(gen[4619]),
			.E(gen[4621]),

			.SO(gen[4714]),
			.S(gen[4715]),
			.SE(gen[4716]),

			.SELF(gen[4620]),
			.cell_state(gen[4620])
		); 

/******************* CELL 4621 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4621 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4525]),
			.N(gen[4526]),
			.NE(gen[4527]),

			.O(gen[4620]),
			.E(gen[4622]),

			.SO(gen[4715]),
			.S(gen[4716]),
			.SE(gen[4717]),

			.SELF(gen[4621]),
			.cell_state(gen[4621])
		); 

/******************* CELL 4622 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4622 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4526]),
			.N(gen[4527]),
			.NE(gen[4528]),

			.O(gen[4621]),
			.E(gen[4623]),

			.SO(gen[4716]),
			.S(gen[4717]),
			.SE(gen[4718]),

			.SELF(gen[4622]),
			.cell_state(gen[4622])
		); 

/******************* CELL 4623 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4623 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4527]),
			.N(gen[4528]),
			.NE(gen[4529]),

			.O(gen[4622]),
			.E(gen[4624]),

			.SO(gen[4717]),
			.S(gen[4718]),
			.SE(gen[4719]),

			.SELF(gen[4623]),
			.cell_state(gen[4623])
		); 

/******************* CELL 4624 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4624 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4528]),
			.N(gen[4529]),
			.NE(gen[4530]),

			.O(gen[4623]),
			.E(gen[4625]),

			.SO(gen[4718]),
			.S(gen[4719]),
			.SE(gen[4720]),

			.SELF(gen[4624]),
			.cell_state(gen[4624])
		); 

/******************* CELL 4625 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4625 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4529]),
			.N(gen[4530]),
			.NE(gen[4531]),

			.O(gen[4624]),
			.E(gen[4626]),

			.SO(gen[4719]),
			.S(gen[4720]),
			.SE(gen[4721]),

			.SELF(gen[4625]),
			.cell_state(gen[4625])
		); 

/******************* CELL 4626 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4626 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4530]),
			.N(gen[4531]),
			.NE(gen[4532]),

			.O(gen[4625]),
			.E(gen[4627]),

			.SO(gen[4720]),
			.S(gen[4721]),
			.SE(gen[4722]),

			.SELF(gen[4626]),
			.cell_state(gen[4626])
		); 

/******************* CELL 4627 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4627 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4531]),
			.N(gen[4532]),
			.NE(gen[4533]),

			.O(gen[4626]),
			.E(gen[4628]),

			.SO(gen[4721]),
			.S(gen[4722]),
			.SE(gen[4723]),

			.SELF(gen[4627]),
			.cell_state(gen[4627])
		); 

/******************* CELL 4628 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4628 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4532]),
			.N(gen[4533]),
			.NE(gen[4534]),

			.O(gen[4627]),
			.E(gen[4629]),

			.SO(gen[4722]),
			.S(gen[4723]),
			.SE(gen[4724]),

			.SELF(gen[4628]),
			.cell_state(gen[4628])
		); 

/******************* CELL 4629 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4629 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4533]),
			.N(gen[4534]),
			.NE(gen[4535]),

			.O(gen[4628]),
			.E(gen[4630]),

			.SO(gen[4723]),
			.S(gen[4724]),
			.SE(gen[4725]),

			.SELF(gen[4629]),
			.cell_state(gen[4629])
		); 

/******************* CELL 4630 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4630 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4534]),
			.N(gen[4535]),
			.NE(gen[4536]),

			.O(gen[4629]),
			.E(gen[4631]),

			.SO(gen[4724]),
			.S(gen[4725]),
			.SE(gen[4726]),

			.SELF(gen[4630]),
			.cell_state(gen[4630])
		); 

/******************* CELL 4631 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4631 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4535]),
			.N(gen[4536]),
			.NE(gen[4537]),

			.O(gen[4630]),
			.E(gen[4632]),

			.SO(gen[4725]),
			.S(gen[4726]),
			.SE(gen[4727]),

			.SELF(gen[4631]),
			.cell_state(gen[4631])
		); 

/******************* CELL 4632 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4632 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4536]),
			.N(gen[4537]),
			.NE(gen[4538]),

			.O(gen[4631]),
			.E(gen[4633]),

			.SO(gen[4726]),
			.S(gen[4727]),
			.SE(gen[4728]),

			.SELF(gen[4632]),
			.cell_state(gen[4632])
		); 

/******************* CELL 4633 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4633 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4537]),
			.N(gen[4538]),
			.NE(gen[4539]),

			.O(gen[4632]),
			.E(gen[4634]),

			.SO(gen[4727]),
			.S(gen[4728]),
			.SE(gen[4729]),

			.SELF(gen[4633]),
			.cell_state(gen[4633])
		); 

/******************* CELL 4634 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4634 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4538]),
			.N(gen[4539]),
			.NE(gen[4540]),

			.O(gen[4633]),
			.E(gen[4635]),

			.SO(gen[4728]),
			.S(gen[4729]),
			.SE(gen[4730]),

			.SELF(gen[4634]),
			.cell_state(gen[4634])
		); 

/******************* CELL 4635 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4635 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4539]),
			.N(gen[4540]),
			.NE(gen[4541]),

			.O(gen[4634]),
			.E(gen[4636]),

			.SO(gen[4729]),
			.S(gen[4730]),
			.SE(gen[4731]),

			.SELF(gen[4635]),
			.cell_state(gen[4635])
		); 

/******************* CELL 4636 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4636 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4540]),
			.N(gen[4541]),
			.NE(gen[4542]),

			.O(gen[4635]),
			.E(gen[4637]),

			.SO(gen[4730]),
			.S(gen[4731]),
			.SE(gen[4732]),

			.SELF(gen[4636]),
			.cell_state(gen[4636])
		); 

/******************* CELL 4637 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4637 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4541]),
			.N(gen[4542]),
			.NE(gen[4543]),

			.O(gen[4636]),
			.E(gen[4638]),

			.SO(gen[4731]),
			.S(gen[4732]),
			.SE(gen[4733]),

			.SELF(gen[4637]),
			.cell_state(gen[4637])
		); 

/******************* CELL 4638 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4638 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4542]),
			.N(gen[4543]),
			.NE(gen[4544]),

			.O(gen[4637]),
			.E(gen[4639]),

			.SO(gen[4732]),
			.S(gen[4733]),
			.SE(gen[4734]),

			.SELF(gen[4638]),
			.cell_state(gen[4638])
		); 

/******************* CELL 4639 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4639 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4543]),
			.N(gen[4544]),
			.NE(gen[4545]),

			.O(gen[4638]),
			.E(gen[4640]),

			.SO(gen[4733]),
			.S(gen[4734]),
			.SE(gen[4735]),

			.SELF(gen[4639]),
			.cell_state(gen[4639])
		); 

/******************* CELL 4640 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4640 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4544]),
			.N(gen[4545]),
			.NE(gen[4546]),

			.O(gen[4639]),
			.E(gen[4641]),

			.SO(gen[4734]),
			.S(gen[4735]),
			.SE(gen[4736]),

			.SELF(gen[4640]),
			.cell_state(gen[4640])
		); 

/******************* CELL 4641 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4641 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4545]),
			.N(gen[4546]),
			.NE(gen[4547]),

			.O(gen[4640]),
			.E(gen[4642]),

			.SO(gen[4735]),
			.S(gen[4736]),
			.SE(gen[4737]),

			.SELF(gen[4641]),
			.cell_state(gen[4641])
		); 

/******************* CELL 4642 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4642 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4546]),
			.N(gen[4547]),
			.NE(gen[4548]),

			.O(gen[4641]),
			.E(gen[4643]),

			.SO(gen[4736]),
			.S(gen[4737]),
			.SE(gen[4738]),

			.SELF(gen[4642]),
			.cell_state(gen[4642])
		); 

/******************* CELL 4643 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4643 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4547]),
			.N(gen[4548]),
			.NE(gen[4549]),

			.O(gen[4642]),
			.E(gen[4644]),

			.SO(gen[4737]),
			.S(gen[4738]),
			.SE(gen[4739]),

			.SELF(gen[4643]),
			.cell_state(gen[4643])
		); 

/******************* CELL 4644 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4644 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4548]),
			.N(gen[4549]),
			.NE(gen[4550]),

			.O(gen[4643]),
			.E(gen[4645]),

			.SO(gen[4738]),
			.S(gen[4739]),
			.SE(gen[4740]),

			.SELF(gen[4644]),
			.cell_state(gen[4644])
		); 

/******************* CELL 4645 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4645 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4549]),
			.N(gen[4550]),
			.NE(gen[4551]),

			.O(gen[4644]),
			.E(gen[4646]),

			.SO(gen[4739]),
			.S(gen[4740]),
			.SE(gen[4741]),

			.SELF(gen[4645]),
			.cell_state(gen[4645])
		); 

/******************* CELL 4646 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4646 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4550]),
			.N(gen[4551]),
			.NE(gen[4552]),

			.O(gen[4645]),
			.E(gen[4647]),

			.SO(gen[4740]),
			.S(gen[4741]),
			.SE(gen[4742]),

			.SELF(gen[4646]),
			.cell_state(gen[4646])
		); 

/******************* CELL 4647 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4647 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4551]),
			.N(gen[4552]),
			.NE(gen[4553]),

			.O(gen[4646]),
			.E(gen[4648]),

			.SO(gen[4741]),
			.S(gen[4742]),
			.SE(gen[4743]),

			.SELF(gen[4647]),
			.cell_state(gen[4647])
		); 

/******************* CELL 4648 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4648 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4552]),
			.N(gen[4553]),
			.NE(gen[4554]),

			.O(gen[4647]),
			.E(gen[4649]),

			.SO(gen[4742]),
			.S(gen[4743]),
			.SE(gen[4744]),

			.SELF(gen[4648]),
			.cell_state(gen[4648])
		); 

/******************* CELL 4649 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4649 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4553]),
			.N(gen[4554]),
			.NE(gen[4555]),

			.O(gen[4648]),
			.E(gen[4650]),

			.SO(gen[4743]),
			.S(gen[4744]),
			.SE(gen[4745]),

			.SELF(gen[4649]),
			.cell_state(gen[4649])
		); 

/******************* CELL 4650 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4650 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4554]),
			.N(gen[4555]),
			.NE(gen[4556]),

			.O(gen[4649]),
			.E(gen[4651]),

			.SO(gen[4744]),
			.S(gen[4745]),
			.SE(gen[4746]),

			.SELF(gen[4650]),
			.cell_state(gen[4650])
		); 

/******************* CELL 4651 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4651 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4555]),
			.N(gen[4556]),
			.NE(gen[4557]),

			.O(gen[4650]),
			.E(gen[4652]),

			.SO(gen[4745]),
			.S(gen[4746]),
			.SE(gen[4747]),

			.SELF(gen[4651]),
			.cell_state(gen[4651])
		); 

/******************* CELL 4652 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4652 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4556]),
			.N(gen[4557]),
			.NE(gen[4558]),

			.O(gen[4651]),
			.E(gen[4653]),

			.SO(gen[4746]),
			.S(gen[4747]),
			.SE(gen[4748]),

			.SELF(gen[4652]),
			.cell_state(gen[4652])
		); 

/******************* CELL 4653 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4653 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4557]),
			.N(gen[4558]),
			.NE(gen[4559]),

			.O(gen[4652]),
			.E(gen[4654]),

			.SO(gen[4747]),
			.S(gen[4748]),
			.SE(gen[4749]),

			.SELF(gen[4653]),
			.cell_state(gen[4653])
		); 

/******************* CELL 4654 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4654 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4558]),
			.N(gen[4559]),
			.NE(gen[4558]),

			.O(gen[4653]),
			.E(gen[4653]),

			.SO(gen[4748]),
			.S(gen[4749]),
			.SE(gen[4748]),

			.SELF(gen[4654]),
			.cell_state(gen[4654])
		); 

/******************* CELL 4655 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4655 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4561]),
			.N(gen[4560]),
			.NE(gen[4561]),

			.O(gen[4656]),
			.E(gen[4656]),

			.SO(gen[4751]),
			.S(gen[4750]),
			.SE(gen[4751]),

			.SELF(gen[4655]),
			.cell_state(gen[4655])
		); 

/******************* CELL 4656 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4656 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4560]),
			.N(gen[4561]),
			.NE(gen[4562]),

			.O(gen[4655]),
			.E(gen[4657]),

			.SO(gen[4750]),
			.S(gen[4751]),
			.SE(gen[4752]),

			.SELF(gen[4656]),
			.cell_state(gen[4656])
		); 

/******************* CELL 4657 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4657 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4561]),
			.N(gen[4562]),
			.NE(gen[4563]),

			.O(gen[4656]),
			.E(gen[4658]),

			.SO(gen[4751]),
			.S(gen[4752]),
			.SE(gen[4753]),

			.SELF(gen[4657]),
			.cell_state(gen[4657])
		); 

/******************* CELL 4658 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4658 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4562]),
			.N(gen[4563]),
			.NE(gen[4564]),

			.O(gen[4657]),
			.E(gen[4659]),

			.SO(gen[4752]),
			.S(gen[4753]),
			.SE(gen[4754]),

			.SELF(gen[4658]),
			.cell_state(gen[4658])
		); 

/******************* CELL 4659 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4659 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4563]),
			.N(gen[4564]),
			.NE(gen[4565]),

			.O(gen[4658]),
			.E(gen[4660]),

			.SO(gen[4753]),
			.S(gen[4754]),
			.SE(gen[4755]),

			.SELF(gen[4659]),
			.cell_state(gen[4659])
		); 

/******************* CELL 4660 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4660 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4564]),
			.N(gen[4565]),
			.NE(gen[4566]),

			.O(gen[4659]),
			.E(gen[4661]),

			.SO(gen[4754]),
			.S(gen[4755]),
			.SE(gen[4756]),

			.SELF(gen[4660]),
			.cell_state(gen[4660])
		); 

/******************* CELL 4661 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4661 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4565]),
			.N(gen[4566]),
			.NE(gen[4567]),

			.O(gen[4660]),
			.E(gen[4662]),

			.SO(gen[4755]),
			.S(gen[4756]),
			.SE(gen[4757]),

			.SELF(gen[4661]),
			.cell_state(gen[4661])
		); 

/******************* CELL 4662 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4662 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4566]),
			.N(gen[4567]),
			.NE(gen[4568]),

			.O(gen[4661]),
			.E(gen[4663]),

			.SO(gen[4756]),
			.S(gen[4757]),
			.SE(gen[4758]),

			.SELF(gen[4662]),
			.cell_state(gen[4662])
		); 

/******************* CELL 4663 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4663 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4567]),
			.N(gen[4568]),
			.NE(gen[4569]),

			.O(gen[4662]),
			.E(gen[4664]),

			.SO(gen[4757]),
			.S(gen[4758]),
			.SE(gen[4759]),

			.SELF(gen[4663]),
			.cell_state(gen[4663])
		); 

/******************* CELL 4664 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4664 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4568]),
			.N(gen[4569]),
			.NE(gen[4570]),

			.O(gen[4663]),
			.E(gen[4665]),

			.SO(gen[4758]),
			.S(gen[4759]),
			.SE(gen[4760]),

			.SELF(gen[4664]),
			.cell_state(gen[4664])
		); 

/******************* CELL 4665 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4665 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4569]),
			.N(gen[4570]),
			.NE(gen[4571]),

			.O(gen[4664]),
			.E(gen[4666]),

			.SO(gen[4759]),
			.S(gen[4760]),
			.SE(gen[4761]),

			.SELF(gen[4665]),
			.cell_state(gen[4665])
		); 

/******************* CELL 4666 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4666 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4570]),
			.N(gen[4571]),
			.NE(gen[4572]),

			.O(gen[4665]),
			.E(gen[4667]),

			.SO(gen[4760]),
			.S(gen[4761]),
			.SE(gen[4762]),

			.SELF(gen[4666]),
			.cell_state(gen[4666])
		); 

/******************* CELL 4667 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4667 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4571]),
			.N(gen[4572]),
			.NE(gen[4573]),

			.O(gen[4666]),
			.E(gen[4668]),

			.SO(gen[4761]),
			.S(gen[4762]),
			.SE(gen[4763]),

			.SELF(gen[4667]),
			.cell_state(gen[4667])
		); 

/******************* CELL 4668 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4668 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4572]),
			.N(gen[4573]),
			.NE(gen[4574]),

			.O(gen[4667]),
			.E(gen[4669]),

			.SO(gen[4762]),
			.S(gen[4763]),
			.SE(gen[4764]),

			.SELF(gen[4668]),
			.cell_state(gen[4668])
		); 

/******************* CELL 4669 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4669 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4573]),
			.N(gen[4574]),
			.NE(gen[4575]),

			.O(gen[4668]),
			.E(gen[4670]),

			.SO(gen[4763]),
			.S(gen[4764]),
			.SE(gen[4765]),

			.SELF(gen[4669]),
			.cell_state(gen[4669])
		); 

/******************* CELL 4670 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4670 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4574]),
			.N(gen[4575]),
			.NE(gen[4576]),

			.O(gen[4669]),
			.E(gen[4671]),

			.SO(gen[4764]),
			.S(gen[4765]),
			.SE(gen[4766]),

			.SELF(gen[4670]),
			.cell_state(gen[4670])
		); 

/******************* CELL 4671 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4671 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4575]),
			.N(gen[4576]),
			.NE(gen[4577]),

			.O(gen[4670]),
			.E(gen[4672]),

			.SO(gen[4765]),
			.S(gen[4766]),
			.SE(gen[4767]),

			.SELF(gen[4671]),
			.cell_state(gen[4671])
		); 

/******************* CELL 4672 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4672 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4576]),
			.N(gen[4577]),
			.NE(gen[4578]),

			.O(gen[4671]),
			.E(gen[4673]),

			.SO(gen[4766]),
			.S(gen[4767]),
			.SE(gen[4768]),

			.SELF(gen[4672]),
			.cell_state(gen[4672])
		); 

/******************* CELL 4673 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4673 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4577]),
			.N(gen[4578]),
			.NE(gen[4579]),

			.O(gen[4672]),
			.E(gen[4674]),

			.SO(gen[4767]),
			.S(gen[4768]),
			.SE(gen[4769]),

			.SELF(gen[4673]),
			.cell_state(gen[4673])
		); 

/******************* CELL 4674 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4674 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4578]),
			.N(gen[4579]),
			.NE(gen[4580]),

			.O(gen[4673]),
			.E(gen[4675]),

			.SO(gen[4768]),
			.S(gen[4769]),
			.SE(gen[4770]),

			.SELF(gen[4674]),
			.cell_state(gen[4674])
		); 

/******************* CELL 4675 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4675 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4579]),
			.N(gen[4580]),
			.NE(gen[4581]),

			.O(gen[4674]),
			.E(gen[4676]),

			.SO(gen[4769]),
			.S(gen[4770]),
			.SE(gen[4771]),

			.SELF(gen[4675]),
			.cell_state(gen[4675])
		); 

/******************* CELL 4676 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4676 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4580]),
			.N(gen[4581]),
			.NE(gen[4582]),

			.O(gen[4675]),
			.E(gen[4677]),

			.SO(gen[4770]),
			.S(gen[4771]),
			.SE(gen[4772]),

			.SELF(gen[4676]),
			.cell_state(gen[4676])
		); 

/******************* CELL 4677 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4677 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4581]),
			.N(gen[4582]),
			.NE(gen[4583]),

			.O(gen[4676]),
			.E(gen[4678]),

			.SO(gen[4771]),
			.S(gen[4772]),
			.SE(gen[4773]),

			.SELF(gen[4677]),
			.cell_state(gen[4677])
		); 

/******************* CELL 4678 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4678 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4582]),
			.N(gen[4583]),
			.NE(gen[4584]),

			.O(gen[4677]),
			.E(gen[4679]),

			.SO(gen[4772]),
			.S(gen[4773]),
			.SE(gen[4774]),

			.SELF(gen[4678]),
			.cell_state(gen[4678])
		); 

/******************* CELL 4679 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4679 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4583]),
			.N(gen[4584]),
			.NE(gen[4585]),

			.O(gen[4678]),
			.E(gen[4680]),

			.SO(gen[4773]),
			.S(gen[4774]),
			.SE(gen[4775]),

			.SELF(gen[4679]),
			.cell_state(gen[4679])
		); 

/******************* CELL 4680 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4680 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4584]),
			.N(gen[4585]),
			.NE(gen[4586]),

			.O(gen[4679]),
			.E(gen[4681]),

			.SO(gen[4774]),
			.S(gen[4775]),
			.SE(gen[4776]),

			.SELF(gen[4680]),
			.cell_state(gen[4680])
		); 

/******************* CELL 4681 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4681 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4585]),
			.N(gen[4586]),
			.NE(gen[4587]),

			.O(gen[4680]),
			.E(gen[4682]),

			.SO(gen[4775]),
			.S(gen[4776]),
			.SE(gen[4777]),

			.SELF(gen[4681]),
			.cell_state(gen[4681])
		); 

/******************* CELL 4682 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4682 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4586]),
			.N(gen[4587]),
			.NE(gen[4588]),

			.O(gen[4681]),
			.E(gen[4683]),

			.SO(gen[4776]),
			.S(gen[4777]),
			.SE(gen[4778]),

			.SELF(gen[4682]),
			.cell_state(gen[4682])
		); 

/******************* CELL 4683 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4683 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4587]),
			.N(gen[4588]),
			.NE(gen[4589]),

			.O(gen[4682]),
			.E(gen[4684]),

			.SO(gen[4777]),
			.S(gen[4778]),
			.SE(gen[4779]),

			.SELF(gen[4683]),
			.cell_state(gen[4683])
		); 

/******************* CELL 4684 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4684 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4588]),
			.N(gen[4589]),
			.NE(gen[4590]),

			.O(gen[4683]),
			.E(gen[4685]),

			.SO(gen[4778]),
			.S(gen[4779]),
			.SE(gen[4780]),

			.SELF(gen[4684]),
			.cell_state(gen[4684])
		); 

/******************* CELL 4685 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4685 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4589]),
			.N(gen[4590]),
			.NE(gen[4591]),

			.O(gen[4684]),
			.E(gen[4686]),

			.SO(gen[4779]),
			.S(gen[4780]),
			.SE(gen[4781]),

			.SELF(gen[4685]),
			.cell_state(gen[4685])
		); 

/******************* CELL 4686 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4686 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4590]),
			.N(gen[4591]),
			.NE(gen[4592]),

			.O(gen[4685]),
			.E(gen[4687]),

			.SO(gen[4780]),
			.S(gen[4781]),
			.SE(gen[4782]),

			.SELF(gen[4686]),
			.cell_state(gen[4686])
		); 

/******************* CELL 4687 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4687 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4591]),
			.N(gen[4592]),
			.NE(gen[4593]),

			.O(gen[4686]),
			.E(gen[4688]),

			.SO(gen[4781]),
			.S(gen[4782]),
			.SE(gen[4783]),

			.SELF(gen[4687]),
			.cell_state(gen[4687])
		); 

/******************* CELL 4688 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4688 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4592]),
			.N(gen[4593]),
			.NE(gen[4594]),

			.O(gen[4687]),
			.E(gen[4689]),

			.SO(gen[4782]),
			.S(gen[4783]),
			.SE(gen[4784]),

			.SELF(gen[4688]),
			.cell_state(gen[4688])
		); 

/******************* CELL 4689 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4689 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4593]),
			.N(gen[4594]),
			.NE(gen[4595]),

			.O(gen[4688]),
			.E(gen[4690]),

			.SO(gen[4783]),
			.S(gen[4784]),
			.SE(gen[4785]),

			.SELF(gen[4689]),
			.cell_state(gen[4689])
		); 

/******************* CELL 4690 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4690 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4594]),
			.N(gen[4595]),
			.NE(gen[4596]),

			.O(gen[4689]),
			.E(gen[4691]),

			.SO(gen[4784]),
			.S(gen[4785]),
			.SE(gen[4786]),

			.SELF(gen[4690]),
			.cell_state(gen[4690])
		); 

/******************* CELL 4691 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4691 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4595]),
			.N(gen[4596]),
			.NE(gen[4597]),

			.O(gen[4690]),
			.E(gen[4692]),

			.SO(gen[4785]),
			.S(gen[4786]),
			.SE(gen[4787]),

			.SELF(gen[4691]),
			.cell_state(gen[4691])
		); 

/******************* CELL 4692 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4692 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4596]),
			.N(gen[4597]),
			.NE(gen[4598]),

			.O(gen[4691]),
			.E(gen[4693]),

			.SO(gen[4786]),
			.S(gen[4787]),
			.SE(gen[4788]),

			.SELF(gen[4692]),
			.cell_state(gen[4692])
		); 

/******************* CELL 4693 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4693 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4597]),
			.N(gen[4598]),
			.NE(gen[4599]),

			.O(gen[4692]),
			.E(gen[4694]),

			.SO(gen[4787]),
			.S(gen[4788]),
			.SE(gen[4789]),

			.SELF(gen[4693]),
			.cell_state(gen[4693])
		); 

/******************* CELL 4694 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4694 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4598]),
			.N(gen[4599]),
			.NE(gen[4600]),

			.O(gen[4693]),
			.E(gen[4695]),

			.SO(gen[4788]),
			.S(gen[4789]),
			.SE(gen[4790]),

			.SELF(gen[4694]),
			.cell_state(gen[4694])
		); 

/******************* CELL 4695 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4695 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4599]),
			.N(gen[4600]),
			.NE(gen[4601]),

			.O(gen[4694]),
			.E(gen[4696]),

			.SO(gen[4789]),
			.S(gen[4790]),
			.SE(gen[4791]),

			.SELF(gen[4695]),
			.cell_state(gen[4695])
		); 

/******************* CELL 4696 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4696 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4600]),
			.N(gen[4601]),
			.NE(gen[4602]),

			.O(gen[4695]),
			.E(gen[4697]),

			.SO(gen[4790]),
			.S(gen[4791]),
			.SE(gen[4792]),

			.SELF(gen[4696]),
			.cell_state(gen[4696])
		); 

/******************* CELL 4697 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4697 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4601]),
			.N(gen[4602]),
			.NE(gen[4603]),

			.O(gen[4696]),
			.E(gen[4698]),

			.SO(gen[4791]),
			.S(gen[4792]),
			.SE(gen[4793]),

			.SELF(gen[4697]),
			.cell_state(gen[4697])
		); 

/******************* CELL 4698 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4698 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4602]),
			.N(gen[4603]),
			.NE(gen[4604]),

			.O(gen[4697]),
			.E(gen[4699]),

			.SO(gen[4792]),
			.S(gen[4793]),
			.SE(gen[4794]),

			.SELF(gen[4698]),
			.cell_state(gen[4698])
		); 

/******************* CELL 4699 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4699 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4603]),
			.N(gen[4604]),
			.NE(gen[4605]),

			.O(gen[4698]),
			.E(gen[4700]),

			.SO(gen[4793]),
			.S(gen[4794]),
			.SE(gen[4795]),

			.SELF(gen[4699]),
			.cell_state(gen[4699])
		); 

/******************* CELL 4700 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4700 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4604]),
			.N(gen[4605]),
			.NE(gen[4606]),

			.O(gen[4699]),
			.E(gen[4701]),

			.SO(gen[4794]),
			.S(gen[4795]),
			.SE(gen[4796]),

			.SELF(gen[4700]),
			.cell_state(gen[4700])
		); 

/******************* CELL 4701 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4701 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4605]),
			.N(gen[4606]),
			.NE(gen[4607]),

			.O(gen[4700]),
			.E(gen[4702]),

			.SO(gen[4795]),
			.S(gen[4796]),
			.SE(gen[4797]),

			.SELF(gen[4701]),
			.cell_state(gen[4701])
		); 

/******************* CELL 4702 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4702 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4606]),
			.N(gen[4607]),
			.NE(gen[4608]),

			.O(gen[4701]),
			.E(gen[4703]),

			.SO(gen[4796]),
			.S(gen[4797]),
			.SE(gen[4798]),

			.SELF(gen[4702]),
			.cell_state(gen[4702])
		); 

/******************* CELL 4703 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4703 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4607]),
			.N(gen[4608]),
			.NE(gen[4609]),

			.O(gen[4702]),
			.E(gen[4704]),

			.SO(gen[4797]),
			.S(gen[4798]),
			.SE(gen[4799]),

			.SELF(gen[4703]),
			.cell_state(gen[4703])
		); 

/******************* CELL 4704 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4704 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4608]),
			.N(gen[4609]),
			.NE(gen[4610]),

			.O(gen[4703]),
			.E(gen[4705]),

			.SO(gen[4798]),
			.S(gen[4799]),
			.SE(gen[4800]),

			.SELF(gen[4704]),
			.cell_state(gen[4704])
		); 

/******************* CELL 4705 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4705 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4609]),
			.N(gen[4610]),
			.NE(gen[4611]),

			.O(gen[4704]),
			.E(gen[4706]),

			.SO(gen[4799]),
			.S(gen[4800]),
			.SE(gen[4801]),

			.SELF(gen[4705]),
			.cell_state(gen[4705])
		); 

/******************* CELL 4706 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4706 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4610]),
			.N(gen[4611]),
			.NE(gen[4612]),

			.O(gen[4705]),
			.E(gen[4707]),

			.SO(gen[4800]),
			.S(gen[4801]),
			.SE(gen[4802]),

			.SELF(gen[4706]),
			.cell_state(gen[4706])
		); 

/******************* CELL 4707 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4707 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4611]),
			.N(gen[4612]),
			.NE(gen[4613]),

			.O(gen[4706]),
			.E(gen[4708]),

			.SO(gen[4801]),
			.S(gen[4802]),
			.SE(gen[4803]),

			.SELF(gen[4707]),
			.cell_state(gen[4707])
		); 

/******************* CELL 4708 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4708 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4612]),
			.N(gen[4613]),
			.NE(gen[4614]),

			.O(gen[4707]),
			.E(gen[4709]),

			.SO(gen[4802]),
			.S(gen[4803]),
			.SE(gen[4804]),

			.SELF(gen[4708]),
			.cell_state(gen[4708])
		); 

/******************* CELL 4709 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4709 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4613]),
			.N(gen[4614]),
			.NE(gen[4615]),

			.O(gen[4708]),
			.E(gen[4710]),

			.SO(gen[4803]),
			.S(gen[4804]),
			.SE(gen[4805]),

			.SELF(gen[4709]),
			.cell_state(gen[4709])
		); 

/******************* CELL 4710 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4710 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4614]),
			.N(gen[4615]),
			.NE(gen[4616]),

			.O(gen[4709]),
			.E(gen[4711]),

			.SO(gen[4804]),
			.S(gen[4805]),
			.SE(gen[4806]),

			.SELF(gen[4710]),
			.cell_state(gen[4710])
		); 

/******************* CELL 4711 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4711 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4615]),
			.N(gen[4616]),
			.NE(gen[4617]),

			.O(gen[4710]),
			.E(gen[4712]),

			.SO(gen[4805]),
			.S(gen[4806]),
			.SE(gen[4807]),

			.SELF(gen[4711]),
			.cell_state(gen[4711])
		); 

/******************* CELL 4712 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4712 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4616]),
			.N(gen[4617]),
			.NE(gen[4618]),

			.O(gen[4711]),
			.E(gen[4713]),

			.SO(gen[4806]),
			.S(gen[4807]),
			.SE(gen[4808]),

			.SELF(gen[4712]),
			.cell_state(gen[4712])
		); 

/******************* CELL 4713 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4713 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4617]),
			.N(gen[4618]),
			.NE(gen[4619]),

			.O(gen[4712]),
			.E(gen[4714]),

			.SO(gen[4807]),
			.S(gen[4808]),
			.SE(gen[4809]),

			.SELF(gen[4713]),
			.cell_state(gen[4713])
		); 

/******************* CELL 4714 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4714 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4618]),
			.N(gen[4619]),
			.NE(gen[4620]),

			.O(gen[4713]),
			.E(gen[4715]),

			.SO(gen[4808]),
			.S(gen[4809]),
			.SE(gen[4810]),

			.SELF(gen[4714]),
			.cell_state(gen[4714])
		); 

/******************* CELL 4715 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4715 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4619]),
			.N(gen[4620]),
			.NE(gen[4621]),

			.O(gen[4714]),
			.E(gen[4716]),

			.SO(gen[4809]),
			.S(gen[4810]),
			.SE(gen[4811]),

			.SELF(gen[4715]),
			.cell_state(gen[4715])
		); 

/******************* CELL 4716 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4716 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4620]),
			.N(gen[4621]),
			.NE(gen[4622]),

			.O(gen[4715]),
			.E(gen[4717]),

			.SO(gen[4810]),
			.S(gen[4811]),
			.SE(gen[4812]),

			.SELF(gen[4716]),
			.cell_state(gen[4716])
		); 

/******************* CELL 4717 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4717 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4621]),
			.N(gen[4622]),
			.NE(gen[4623]),

			.O(gen[4716]),
			.E(gen[4718]),

			.SO(gen[4811]),
			.S(gen[4812]),
			.SE(gen[4813]),

			.SELF(gen[4717]),
			.cell_state(gen[4717])
		); 

/******************* CELL 4718 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4718 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4622]),
			.N(gen[4623]),
			.NE(gen[4624]),

			.O(gen[4717]),
			.E(gen[4719]),

			.SO(gen[4812]),
			.S(gen[4813]),
			.SE(gen[4814]),

			.SELF(gen[4718]),
			.cell_state(gen[4718])
		); 

/******************* CELL 4719 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4719 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4623]),
			.N(gen[4624]),
			.NE(gen[4625]),

			.O(gen[4718]),
			.E(gen[4720]),

			.SO(gen[4813]),
			.S(gen[4814]),
			.SE(gen[4815]),

			.SELF(gen[4719]),
			.cell_state(gen[4719])
		); 

/******************* CELL 4720 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4720 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4624]),
			.N(gen[4625]),
			.NE(gen[4626]),

			.O(gen[4719]),
			.E(gen[4721]),

			.SO(gen[4814]),
			.S(gen[4815]),
			.SE(gen[4816]),

			.SELF(gen[4720]),
			.cell_state(gen[4720])
		); 

/******************* CELL 4721 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4721 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4625]),
			.N(gen[4626]),
			.NE(gen[4627]),

			.O(gen[4720]),
			.E(gen[4722]),

			.SO(gen[4815]),
			.S(gen[4816]),
			.SE(gen[4817]),

			.SELF(gen[4721]),
			.cell_state(gen[4721])
		); 

/******************* CELL 4722 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4722 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4626]),
			.N(gen[4627]),
			.NE(gen[4628]),

			.O(gen[4721]),
			.E(gen[4723]),

			.SO(gen[4816]),
			.S(gen[4817]),
			.SE(gen[4818]),

			.SELF(gen[4722]),
			.cell_state(gen[4722])
		); 

/******************* CELL 4723 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4723 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4627]),
			.N(gen[4628]),
			.NE(gen[4629]),

			.O(gen[4722]),
			.E(gen[4724]),

			.SO(gen[4817]),
			.S(gen[4818]),
			.SE(gen[4819]),

			.SELF(gen[4723]),
			.cell_state(gen[4723])
		); 

/******************* CELL 4724 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4724 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4628]),
			.N(gen[4629]),
			.NE(gen[4630]),

			.O(gen[4723]),
			.E(gen[4725]),

			.SO(gen[4818]),
			.S(gen[4819]),
			.SE(gen[4820]),

			.SELF(gen[4724]),
			.cell_state(gen[4724])
		); 

/******************* CELL 4725 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4725 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4629]),
			.N(gen[4630]),
			.NE(gen[4631]),

			.O(gen[4724]),
			.E(gen[4726]),

			.SO(gen[4819]),
			.S(gen[4820]),
			.SE(gen[4821]),

			.SELF(gen[4725]),
			.cell_state(gen[4725])
		); 

/******************* CELL 4726 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4726 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4630]),
			.N(gen[4631]),
			.NE(gen[4632]),

			.O(gen[4725]),
			.E(gen[4727]),

			.SO(gen[4820]),
			.S(gen[4821]),
			.SE(gen[4822]),

			.SELF(gen[4726]),
			.cell_state(gen[4726])
		); 

/******************* CELL 4727 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4727 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4631]),
			.N(gen[4632]),
			.NE(gen[4633]),

			.O(gen[4726]),
			.E(gen[4728]),

			.SO(gen[4821]),
			.S(gen[4822]),
			.SE(gen[4823]),

			.SELF(gen[4727]),
			.cell_state(gen[4727])
		); 

/******************* CELL 4728 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4728 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4632]),
			.N(gen[4633]),
			.NE(gen[4634]),

			.O(gen[4727]),
			.E(gen[4729]),

			.SO(gen[4822]),
			.S(gen[4823]),
			.SE(gen[4824]),

			.SELF(gen[4728]),
			.cell_state(gen[4728])
		); 

/******************* CELL 4729 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4729 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4633]),
			.N(gen[4634]),
			.NE(gen[4635]),

			.O(gen[4728]),
			.E(gen[4730]),

			.SO(gen[4823]),
			.S(gen[4824]),
			.SE(gen[4825]),

			.SELF(gen[4729]),
			.cell_state(gen[4729])
		); 

/******************* CELL 4730 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4730 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4634]),
			.N(gen[4635]),
			.NE(gen[4636]),

			.O(gen[4729]),
			.E(gen[4731]),

			.SO(gen[4824]),
			.S(gen[4825]),
			.SE(gen[4826]),

			.SELF(gen[4730]),
			.cell_state(gen[4730])
		); 

/******************* CELL 4731 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4731 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4635]),
			.N(gen[4636]),
			.NE(gen[4637]),

			.O(gen[4730]),
			.E(gen[4732]),

			.SO(gen[4825]),
			.S(gen[4826]),
			.SE(gen[4827]),

			.SELF(gen[4731]),
			.cell_state(gen[4731])
		); 

/******************* CELL 4732 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4732 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4636]),
			.N(gen[4637]),
			.NE(gen[4638]),

			.O(gen[4731]),
			.E(gen[4733]),

			.SO(gen[4826]),
			.S(gen[4827]),
			.SE(gen[4828]),

			.SELF(gen[4732]),
			.cell_state(gen[4732])
		); 

/******************* CELL 4733 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4733 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4637]),
			.N(gen[4638]),
			.NE(gen[4639]),

			.O(gen[4732]),
			.E(gen[4734]),

			.SO(gen[4827]),
			.S(gen[4828]),
			.SE(gen[4829]),

			.SELF(gen[4733]),
			.cell_state(gen[4733])
		); 

/******************* CELL 4734 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4734 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4638]),
			.N(gen[4639]),
			.NE(gen[4640]),

			.O(gen[4733]),
			.E(gen[4735]),

			.SO(gen[4828]),
			.S(gen[4829]),
			.SE(gen[4830]),

			.SELF(gen[4734]),
			.cell_state(gen[4734])
		); 

/******************* CELL 4735 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4735 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4639]),
			.N(gen[4640]),
			.NE(gen[4641]),

			.O(gen[4734]),
			.E(gen[4736]),

			.SO(gen[4829]),
			.S(gen[4830]),
			.SE(gen[4831]),

			.SELF(gen[4735]),
			.cell_state(gen[4735])
		); 

/******************* CELL 4736 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4736 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4640]),
			.N(gen[4641]),
			.NE(gen[4642]),

			.O(gen[4735]),
			.E(gen[4737]),

			.SO(gen[4830]),
			.S(gen[4831]),
			.SE(gen[4832]),

			.SELF(gen[4736]),
			.cell_state(gen[4736])
		); 

/******************* CELL 4737 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4737 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4641]),
			.N(gen[4642]),
			.NE(gen[4643]),

			.O(gen[4736]),
			.E(gen[4738]),

			.SO(gen[4831]),
			.S(gen[4832]),
			.SE(gen[4833]),

			.SELF(gen[4737]),
			.cell_state(gen[4737])
		); 

/******************* CELL 4738 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4738 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4642]),
			.N(gen[4643]),
			.NE(gen[4644]),

			.O(gen[4737]),
			.E(gen[4739]),

			.SO(gen[4832]),
			.S(gen[4833]),
			.SE(gen[4834]),

			.SELF(gen[4738]),
			.cell_state(gen[4738])
		); 

/******************* CELL 4739 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4739 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4643]),
			.N(gen[4644]),
			.NE(gen[4645]),

			.O(gen[4738]),
			.E(gen[4740]),

			.SO(gen[4833]),
			.S(gen[4834]),
			.SE(gen[4835]),

			.SELF(gen[4739]),
			.cell_state(gen[4739])
		); 

/******************* CELL 4740 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4740 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4644]),
			.N(gen[4645]),
			.NE(gen[4646]),

			.O(gen[4739]),
			.E(gen[4741]),

			.SO(gen[4834]),
			.S(gen[4835]),
			.SE(gen[4836]),

			.SELF(gen[4740]),
			.cell_state(gen[4740])
		); 

/******************* CELL 4741 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4741 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4645]),
			.N(gen[4646]),
			.NE(gen[4647]),

			.O(gen[4740]),
			.E(gen[4742]),

			.SO(gen[4835]),
			.S(gen[4836]),
			.SE(gen[4837]),

			.SELF(gen[4741]),
			.cell_state(gen[4741])
		); 

/******************* CELL 4742 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4742 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4646]),
			.N(gen[4647]),
			.NE(gen[4648]),

			.O(gen[4741]),
			.E(gen[4743]),

			.SO(gen[4836]),
			.S(gen[4837]),
			.SE(gen[4838]),

			.SELF(gen[4742]),
			.cell_state(gen[4742])
		); 

/******************* CELL 4743 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4743 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4647]),
			.N(gen[4648]),
			.NE(gen[4649]),

			.O(gen[4742]),
			.E(gen[4744]),

			.SO(gen[4837]),
			.S(gen[4838]),
			.SE(gen[4839]),

			.SELF(gen[4743]),
			.cell_state(gen[4743])
		); 

/******************* CELL 4744 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4744 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4648]),
			.N(gen[4649]),
			.NE(gen[4650]),

			.O(gen[4743]),
			.E(gen[4745]),

			.SO(gen[4838]),
			.S(gen[4839]),
			.SE(gen[4840]),

			.SELF(gen[4744]),
			.cell_state(gen[4744])
		); 

/******************* CELL 4745 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4745 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4649]),
			.N(gen[4650]),
			.NE(gen[4651]),

			.O(gen[4744]),
			.E(gen[4746]),

			.SO(gen[4839]),
			.S(gen[4840]),
			.SE(gen[4841]),

			.SELF(gen[4745]),
			.cell_state(gen[4745])
		); 

/******************* CELL 4746 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4746 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4650]),
			.N(gen[4651]),
			.NE(gen[4652]),

			.O(gen[4745]),
			.E(gen[4747]),

			.SO(gen[4840]),
			.S(gen[4841]),
			.SE(gen[4842]),

			.SELF(gen[4746]),
			.cell_state(gen[4746])
		); 

/******************* CELL 4747 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4747 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4651]),
			.N(gen[4652]),
			.NE(gen[4653]),

			.O(gen[4746]),
			.E(gen[4748]),

			.SO(gen[4841]),
			.S(gen[4842]),
			.SE(gen[4843]),

			.SELF(gen[4747]),
			.cell_state(gen[4747])
		); 

/******************* CELL 4748 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4748 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4652]),
			.N(gen[4653]),
			.NE(gen[4654]),

			.O(gen[4747]),
			.E(gen[4749]),

			.SO(gen[4842]),
			.S(gen[4843]),
			.SE(gen[4844]),

			.SELF(gen[4748]),
			.cell_state(gen[4748])
		); 

/******************* CELL 4749 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4749 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4653]),
			.N(gen[4654]),
			.NE(gen[4653]),

			.O(gen[4748]),
			.E(gen[4748]),

			.SO(gen[4843]),
			.S(gen[4844]),
			.SE(gen[4843]),

			.SELF(gen[4749]),
			.cell_state(gen[4749])
		); 

/******************* CELL 4750 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4750 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4656]),
			.N(gen[4655]),
			.NE(gen[4656]),

			.O(gen[4751]),
			.E(gen[4751]),

			.SO(gen[4846]),
			.S(gen[4845]),
			.SE(gen[4846]),

			.SELF(gen[4750]),
			.cell_state(gen[4750])
		); 

/******************* CELL 4751 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4751 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4655]),
			.N(gen[4656]),
			.NE(gen[4657]),

			.O(gen[4750]),
			.E(gen[4752]),

			.SO(gen[4845]),
			.S(gen[4846]),
			.SE(gen[4847]),

			.SELF(gen[4751]),
			.cell_state(gen[4751])
		); 

/******************* CELL 4752 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4752 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4656]),
			.N(gen[4657]),
			.NE(gen[4658]),

			.O(gen[4751]),
			.E(gen[4753]),

			.SO(gen[4846]),
			.S(gen[4847]),
			.SE(gen[4848]),

			.SELF(gen[4752]),
			.cell_state(gen[4752])
		); 

/******************* CELL 4753 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4753 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4657]),
			.N(gen[4658]),
			.NE(gen[4659]),

			.O(gen[4752]),
			.E(gen[4754]),

			.SO(gen[4847]),
			.S(gen[4848]),
			.SE(gen[4849]),

			.SELF(gen[4753]),
			.cell_state(gen[4753])
		); 

/******************* CELL 4754 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4754 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4658]),
			.N(gen[4659]),
			.NE(gen[4660]),

			.O(gen[4753]),
			.E(gen[4755]),

			.SO(gen[4848]),
			.S(gen[4849]),
			.SE(gen[4850]),

			.SELF(gen[4754]),
			.cell_state(gen[4754])
		); 

/******************* CELL 4755 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4755 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4659]),
			.N(gen[4660]),
			.NE(gen[4661]),

			.O(gen[4754]),
			.E(gen[4756]),

			.SO(gen[4849]),
			.S(gen[4850]),
			.SE(gen[4851]),

			.SELF(gen[4755]),
			.cell_state(gen[4755])
		); 

/******************* CELL 4756 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4756 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4660]),
			.N(gen[4661]),
			.NE(gen[4662]),

			.O(gen[4755]),
			.E(gen[4757]),

			.SO(gen[4850]),
			.S(gen[4851]),
			.SE(gen[4852]),

			.SELF(gen[4756]),
			.cell_state(gen[4756])
		); 

/******************* CELL 4757 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4757 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4661]),
			.N(gen[4662]),
			.NE(gen[4663]),

			.O(gen[4756]),
			.E(gen[4758]),

			.SO(gen[4851]),
			.S(gen[4852]),
			.SE(gen[4853]),

			.SELF(gen[4757]),
			.cell_state(gen[4757])
		); 

/******************* CELL 4758 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4758 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4662]),
			.N(gen[4663]),
			.NE(gen[4664]),

			.O(gen[4757]),
			.E(gen[4759]),

			.SO(gen[4852]),
			.S(gen[4853]),
			.SE(gen[4854]),

			.SELF(gen[4758]),
			.cell_state(gen[4758])
		); 

/******************* CELL 4759 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4759 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4663]),
			.N(gen[4664]),
			.NE(gen[4665]),

			.O(gen[4758]),
			.E(gen[4760]),

			.SO(gen[4853]),
			.S(gen[4854]),
			.SE(gen[4855]),

			.SELF(gen[4759]),
			.cell_state(gen[4759])
		); 

/******************* CELL 4760 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4760 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4664]),
			.N(gen[4665]),
			.NE(gen[4666]),

			.O(gen[4759]),
			.E(gen[4761]),

			.SO(gen[4854]),
			.S(gen[4855]),
			.SE(gen[4856]),

			.SELF(gen[4760]),
			.cell_state(gen[4760])
		); 

/******************* CELL 4761 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4761 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4665]),
			.N(gen[4666]),
			.NE(gen[4667]),

			.O(gen[4760]),
			.E(gen[4762]),

			.SO(gen[4855]),
			.S(gen[4856]),
			.SE(gen[4857]),

			.SELF(gen[4761]),
			.cell_state(gen[4761])
		); 

/******************* CELL 4762 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4762 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4666]),
			.N(gen[4667]),
			.NE(gen[4668]),

			.O(gen[4761]),
			.E(gen[4763]),

			.SO(gen[4856]),
			.S(gen[4857]),
			.SE(gen[4858]),

			.SELF(gen[4762]),
			.cell_state(gen[4762])
		); 

/******************* CELL 4763 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4763 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4667]),
			.N(gen[4668]),
			.NE(gen[4669]),

			.O(gen[4762]),
			.E(gen[4764]),

			.SO(gen[4857]),
			.S(gen[4858]),
			.SE(gen[4859]),

			.SELF(gen[4763]),
			.cell_state(gen[4763])
		); 

/******************* CELL 4764 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4764 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4668]),
			.N(gen[4669]),
			.NE(gen[4670]),

			.O(gen[4763]),
			.E(gen[4765]),

			.SO(gen[4858]),
			.S(gen[4859]),
			.SE(gen[4860]),

			.SELF(gen[4764]),
			.cell_state(gen[4764])
		); 

/******************* CELL 4765 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4765 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4669]),
			.N(gen[4670]),
			.NE(gen[4671]),

			.O(gen[4764]),
			.E(gen[4766]),

			.SO(gen[4859]),
			.S(gen[4860]),
			.SE(gen[4861]),

			.SELF(gen[4765]),
			.cell_state(gen[4765])
		); 

/******************* CELL 4766 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4766 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4670]),
			.N(gen[4671]),
			.NE(gen[4672]),

			.O(gen[4765]),
			.E(gen[4767]),

			.SO(gen[4860]),
			.S(gen[4861]),
			.SE(gen[4862]),

			.SELF(gen[4766]),
			.cell_state(gen[4766])
		); 

/******************* CELL 4767 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4767 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4671]),
			.N(gen[4672]),
			.NE(gen[4673]),

			.O(gen[4766]),
			.E(gen[4768]),

			.SO(gen[4861]),
			.S(gen[4862]),
			.SE(gen[4863]),

			.SELF(gen[4767]),
			.cell_state(gen[4767])
		); 

/******************* CELL 4768 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4768 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4672]),
			.N(gen[4673]),
			.NE(gen[4674]),

			.O(gen[4767]),
			.E(gen[4769]),

			.SO(gen[4862]),
			.S(gen[4863]),
			.SE(gen[4864]),

			.SELF(gen[4768]),
			.cell_state(gen[4768])
		); 

/******************* CELL 4769 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4769 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4673]),
			.N(gen[4674]),
			.NE(gen[4675]),

			.O(gen[4768]),
			.E(gen[4770]),

			.SO(gen[4863]),
			.S(gen[4864]),
			.SE(gen[4865]),

			.SELF(gen[4769]),
			.cell_state(gen[4769])
		); 

/******************* CELL 4770 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4770 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4674]),
			.N(gen[4675]),
			.NE(gen[4676]),

			.O(gen[4769]),
			.E(gen[4771]),

			.SO(gen[4864]),
			.S(gen[4865]),
			.SE(gen[4866]),

			.SELF(gen[4770]),
			.cell_state(gen[4770])
		); 

/******************* CELL 4771 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4771 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4675]),
			.N(gen[4676]),
			.NE(gen[4677]),

			.O(gen[4770]),
			.E(gen[4772]),

			.SO(gen[4865]),
			.S(gen[4866]),
			.SE(gen[4867]),

			.SELF(gen[4771]),
			.cell_state(gen[4771])
		); 

/******************* CELL 4772 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4772 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4676]),
			.N(gen[4677]),
			.NE(gen[4678]),

			.O(gen[4771]),
			.E(gen[4773]),

			.SO(gen[4866]),
			.S(gen[4867]),
			.SE(gen[4868]),

			.SELF(gen[4772]),
			.cell_state(gen[4772])
		); 

/******************* CELL 4773 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4773 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4677]),
			.N(gen[4678]),
			.NE(gen[4679]),

			.O(gen[4772]),
			.E(gen[4774]),

			.SO(gen[4867]),
			.S(gen[4868]),
			.SE(gen[4869]),

			.SELF(gen[4773]),
			.cell_state(gen[4773])
		); 

/******************* CELL 4774 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4774 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4678]),
			.N(gen[4679]),
			.NE(gen[4680]),

			.O(gen[4773]),
			.E(gen[4775]),

			.SO(gen[4868]),
			.S(gen[4869]),
			.SE(gen[4870]),

			.SELF(gen[4774]),
			.cell_state(gen[4774])
		); 

/******************* CELL 4775 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4775 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4679]),
			.N(gen[4680]),
			.NE(gen[4681]),

			.O(gen[4774]),
			.E(gen[4776]),

			.SO(gen[4869]),
			.S(gen[4870]),
			.SE(gen[4871]),

			.SELF(gen[4775]),
			.cell_state(gen[4775])
		); 

/******************* CELL 4776 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4776 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4680]),
			.N(gen[4681]),
			.NE(gen[4682]),

			.O(gen[4775]),
			.E(gen[4777]),

			.SO(gen[4870]),
			.S(gen[4871]),
			.SE(gen[4872]),

			.SELF(gen[4776]),
			.cell_state(gen[4776])
		); 

/******************* CELL 4777 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4777 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4681]),
			.N(gen[4682]),
			.NE(gen[4683]),

			.O(gen[4776]),
			.E(gen[4778]),

			.SO(gen[4871]),
			.S(gen[4872]),
			.SE(gen[4873]),

			.SELF(gen[4777]),
			.cell_state(gen[4777])
		); 

/******************* CELL 4778 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4778 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4682]),
			.N(gen[4683]),
			.NE(gen[4684]),

			.O(gen[4777]),
			.E(gen[4779]),

			.SO(gen[4872]),
			.S(gen[4873]),
			.SE(gen[4874]),

			.SELF(gen[4778]),
			.cell_state(gen[4778])
		); 

/******************* CELL 4779 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4779 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4683]),
			.N(gen[4684]),
			.NE(gen[4685]),

			.O(gen[4778]),
			.E(gen[4780]),

			.SO(gen[4873]),
			.S(gen[4874]),
			.SE(gen[4875]),

			.SELF(gen[4779]),
			.cell_state(gen[4779])
		); 

/******************* CELL 4780 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4780 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4684]),
			.N(gen[4685]),
			.NE(gen[4686]),

			.O(gen[4779]),
			.E(gen[4781]),

			.SO(gen[4874]),
			.S(gen[4875]),
			.SE(gen[4876]),

			.SELF(gen[4780]),
			.cell_state(gen[4780])
		); 

/******************* CELL 4781 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4781 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4685]),
			.N(gen[4686]),
			.NE(gen[4687]),

			.O(gen[4780]),
			.E(gen[4782]),

			.SO(gen[4875]),
			.S(gen[4876]),
			.SE(gen[4877]),

			.SELF(gen[4781]),
			.cell_state(gen[4781])
		); 

/******************* CELL 4782 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4782 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4686]),
			.N(gen[4687]),
			.NE(gen[4688]),

			.O(gen[4781]),
			.E(gen[4783]),

			.SO(gen[4876]),
			.S(gen[4877]),
			.SE(gen[4878]),

			.SELF(gen[4782]),
			.cell_state(gen[4782])
		); 

/******************* CELL 4783 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4783 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4687]),
			.N(gen[4688]),
			.NE(gen[4689]),

			.O(gen[4782]),
			.E(gen[4784]),

			.SO(gen[4877]),
			.S(gen[4878]),
			.SE(gen[4879]),

			.SELF(gen[4783]),
			.cell_state(gen[4783])
		); 

/******************* CELL 4784 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4784 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4688]),
			.N(gen[4689]),
			.NE(gen[4690]),

			.O(gen[4783]),
			.E(gen[4785]),

			.SO(gen[4878]),
			.S(gen[4879]),
			.SE(gen[4880]),

			.SELF(gen[4784]),
			.cell_state(gen[4784])
		); 

/******************* CELL 4785 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4785 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4689]),
			.N(gen[4690]),
			.NE(gen[4691]),

			.O(gen[4784]),
			.E(gen[4786]),

			.SO(gen[4879]),
			.S(gen[4880]),
			.SE(gen[4881]),

			.SELF(gen[4785]),
			.cell_state(gen[4785])
		); 

/******************* CELL 4786 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4786 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4690]),
			.N(gen[4691]),
			.NE(gen[4692]),

			.O(gen[4785]),
			.E(gen[4787]),

			.SO(gen[4880]),
			.S(gen[4881]),
			.SE(gen[4882]),

			.SELF(gen[4786]),
			.cell_state(gen[4786])
		); 

/******************* CELL 4787 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4787 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4691]),
			.N(gen[4692]),
			.NE(gen[4693]),

			.O(gen[4786]),
			.E(gen[4788]),

			.SO(gen[4881]),
			.S(gen[4882]),
			.SE(gen[4883]),

			.SELF(gen[4787]),
			.cell_state(gen[4787])
		); 

/******************* CELL 4788 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4788 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4692]),
			.N(gen[4693]),
			.NE(gen[4694]),

			.O(gen[4787]),
			.E(gen[4789]),

			.SO(gen[4882]),
			.S(gen[4883]),
			.SE(gen[4884]),

			.SELF(gen[4788]),
			.cell_state(gen[4788])
		); 

/******************* CELL 4789 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4789 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4693]),
			.N(gen[4694]),
			.NE(gen[4695]),

			.O(gen[4788]),
			.E(gen[4790]),

			.SO(gen[4883]),
			.S(gen[4884]),
			.SE(gen[4885]),

			.SELF(gen[4789]),
			.cell_state(gen[4789])
		); 

/******************* CELL 4790 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4790 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4694]),
			.N(gen[4695]),
			.NE(gen[4696]),

			.O(gen[4789]),
			.E(gen[4791]),

			.SO(gen[4884]),
			.S(gen[4885]),
			.SE(gen[4886]),

			.SELF(gen[4790]),
			.cell_state(gen[4790])
		); 

/******************* CELL 4791 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4791 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4695]),
			.N(gen[4696]),
			.NE(gen[4697]),

			.O(gen[4790]),
			.E(gen[4792]),

			.SO(gen[4885]),
			.S(gen[4886]),
			.SE(gen[4887]),

			.SELF(gen[4791]),
			.cell_state(gen[4791])
		); 

/******************* CELL 4792 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4792 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4696]),
			.N(gen[4697]),
			.NE(gen[4698]),

			.O(gen[4791]),
			.E(gen[4793]),

			.SO(gen[4886]),
			.S(gen[4887]),
			.SE(gen[4888]),

			.SELF(gen[4792]),
			.cell_state(gen[4792])
		); 

/******************* CELL 4793 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4793 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4697]),
			.N(gen[4698]),
			.NE(gen[4699]),

			.O(gen[4792]),
			.E(gen[4794]),

			.SO(gen[4887]),
			.S(gen[4888]),
			.SE(gen[4889]),

			.SELF(gen[4793]),
			.cell_state(gen[4793])
		); 

/******************* CELL 4794 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4794 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4698]),
			.N(gen[4699]),
			.NE(gen[4700]),

			.O(gen[4793]),
			.E(gen[4795]),

			.SO(gen[4888]),
			.S(gen[4889]),
			.SE(gen[4890]),

			.SELF(gen[4794]),
			.cell_state(gen[4794])
		); 

/******************* CELL 4795 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4795 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4699]),
			.N(gen[4700]),
			.NE(gen[4701]),

			.O(gen[4794]),
			.E(gen[4796]),

			.SO(gen[4889]),
			.S(gen[4890]),
			.SE(gen[4891]),

			.SELF(gen[4795]),
			.cell_state(gen[4795])
		); 

/******************* CELL 4796 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4796 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4700]),
			.N(gen[4701]),
			.NE(gen[4702]),

			.O(gen[4795]),
			.E(gen[4797]),

			.SO(gen[4890]),
			.S(gen[4891]),
			.SE(gen[4892]),

			.SELF(gen[4796]),
			.cell_state(gen[4796])
		); 

/******************* CELL 4797 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4797 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4701]),
			.N(gen[4702]),
			.NE(gen[4703]),

			.O(gen[4796]),
			.E(gen[4798]),

			.SO(gen[4891]),
			.S(gen[4892]),
			.SE(gen[4893]),

			.SELF(gen[4797]),
			.cell_state(gen[4797])
		); 

/******************* CELL 4798 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4798 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4702]),
			.N(gen[4703]),
			.NE(gen[4704]),

			.O(gen[4797]),
			.E(gen[4799]),

			.SO(gen[4892]),
			.S(gen[4893]),
			.SE(gen[4894]),

			.SELF(gen[4798]),
			.cell_state(gen[4798])
		); 

/******************* CELL 4799 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4799 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4703]),
			.N(gen[4704]),
			.NE(gen[4705]),

			.O(gen[4798]),
			.E(gen[4800]),

			.SO(gen[4893]),
			.S(gen[4894]),
			.SE(gen[4895]),

			.SELF(gen[4799]),
			.cell_state(gen[4799])
		); 

/******************* CELL 4800 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4800 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4704]),
			.N(gen[4705]),
			.NE(gen[4706]),

			.O(gen[4799]),
			.E(gen[4801]),

			.SO(gen[4894]),
			.S(gen[4895]),
			.SE(gen[4896]),

			.SELF(gen[4800]),
			.cell_state(gen[4800])
		); 

/******************* CELL 4801 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4801 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4705]),
			.N(gen[4706]),
			.NE(gen[4707]),

			.O(gen[4800]),
			.E(gen[4802]),

			.SO(gen[4895]),
			.S(gen[4896]),
			.SE(gen[4897]),

			.SELF(gen[4801]),
			.cell_state(gen[4801])
		); 

/******************* CELL 4802 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4802 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4706]),
			.N(gen[4707]),
			.NE(gen[4708]),

			.O(gen[4801]),
			.E(gen[4803]),

			.SO(gen[4896]),
			.S(gen[4897]),
			.SE(gen[4898]),

			.SELF(gen[4802]),
			.cell_state(gen[4802])
		); 

/******************* CELL 4803 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4803 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4707]),
			.N(gen[4708]),
			.NE(gen[4709]),

			.O(gen[4802]),
			.E(gen[4804]),

			.SO(gen[4897]),
			.S(gen[4898]),
			.SE(gen[4899]),

			.SELF(gen[4803]),
			.cell_state(gen[4803])
		); 

/******************* CELL 4804 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4804 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4708]),
			.N(gen[4709]),
			.NE(gen[4710]),

			.O(gen[4803]),
			.E(gen[4805]),

			.SO(gen[4898]),
			.S(gen[4899]),
			.SE(gen[4900]),

			.SELF(gen[4804]),
			.cell_state(gen[4804])
		); 

/******************* CELL 4805 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4805 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4709]),
			.N(gen[4710]),
			.NE(gen[4711]),

			.O(gen[4804]),
			.E(gen[4806]),

			.SO(gen[4899]),
			.S(gen[4900]),
			.SE(gen[4901]),

			.SELF(gen[4805]),
			.cell_state(gen[4805])
		); 

/******************* CELL 4806 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4806 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4710]),
			.N(gen[4711]),
			.NE(gen[4712]),

			.O(gen[4805]),
			.E(gen[4807]),

			.SO(gen[4900]),
			.S(gen[4901]),
			.SE(gen[4902]),

			.SELF(gen[4806]),
			.cell_state(gen[4806])
		); 

/******************* CELL 4807 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4807 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4711]),
			.N(gen[4712]),
			.NE(gen[4713]),

			.O(gen[4806]),
			.E(gen[4808]),

			.SO(gen[4901]),
			.S(gen[4902]),
			.SE(gen[4903]),

			.SELF(gen[4807]),
			.cell_state(gen[4807])
		); 

/******************* CELL 4808 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4808 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4712]),
			.N(gen[4713]),
			.NE(gen[4714]),

			.O(gen[4807]),
			.E(gen[4809]),

			.SO(gen[4902]),
			.S(gen[4903]),
			.SE(gen[4904]),

			.SELF(gen[4808]),
			.cell_state(gen[4808])
		); 

/******************* CELL 4809 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4809 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4713]),
			.N(gen[4714]),
			.NE(gen[4715]),

			.O(gen[4808]),
			.E(gen[4810]),

			.SO(gen[4903]),
			.S(gen[4904]),
			.SE(gen[4905]),

			.SELF(gen[4809]),
			.cell_state(gen[4809])
		); 

/******************* CELL 4810 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4810 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4714]),
			.N(gen[4715]),
			.NE(gen[4716]),

			.O(gen[4809]),
			.E(gen[4811]),

			.SO(gen[4904]),
			.S(gen[4905]),
			.SE(gen[4906]),

			.SELF(gen[4810]),
			.cell_state(gen[4810])
		); 

/******************* CELL 4811 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4811 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4715]),
			.N(gen[4716]),
			.NE(gen[4717]),

			.O(gen[4810]),
			.E(gen[4812]),

			.SO(gen[4905]),
			.S(gen[4906]),
			.SE(gen[4907]),

			.SELF(gen[4811]),
			.cell_state(gen[4811])
		); 

/******************* CELL 4812 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4812 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4716]),
			.N(gen[4717]),
			.NE(gen[4718]),

			.O(gen[4811]),
			.E(gen[4813]),

			.SO(gen[4906]),
			.S(gen[4907]),
			.SE(gen[4908]),

			.SELF(gen[4812]),
			.cell_state(gen[4812])
		); 

/******************* CELL 4813 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4813 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4717]),
			.N(gen[4718]),
			.NE(gen[4719]),

			.O(gen[4812]),
			.E(gen[4814]),

			.SO(gen[4907]),
			.S(gen[4908]),
			.SE(gen[4909]),

			.SELF(gen[4813]),
			.cell_state(gen[4813])
		); 

/******************* CELL 4814 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4814 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4718]),
			.N(gen[4719]),
			.NE(gen[4720]),

			.O(gen[4813]),
			.E(gen[4815]),

			.SO(gen[4908]),
			.S(gen[4909]),
			.SE(gen[4910]),

			.SELF(gen[4814]),
			.cell_state(gen[4814])
		); 

/******************* CELL 4815 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4815 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4719]),
			.N(gen[4720]),
			.NE(gen[4721]),

			.O(gen[4814]),
			.E(gen[4816]),

			.SO(gen[4909]),
			.S(gen[4910]),
			.SE(gen[4911]),

			.SELF(gen[4815]),
			.cell_state(gen[4815])
		); 

/******************* CELL 4816 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4816 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4720]),
			.N(gen[4721]),
			.NE(gen[4722]),

			.O(gen[4815]),
			.E(gen[4817]),

			.SO(gen[4910]),
			.S(gen[4911]),
			.SE(gen[4912]),

			.SELF(gen[4816]),
			.cell_state(gen[4816])
		); 

/******************* CELL 4817 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4817 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4721]),
			.N(gen[4722]),
			.NE(gen[4723]),

			.O(gen[4816]),
			.E(gen[4818]),

			.SO(gen[4911]),
			.S(gen[4912]),
			.SE(gen[4913]),

			.SELF(gen[4817]),
			.cell_state(gen[4817])
		); 

/******************* CELL 4818 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4818 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4722]),
			.N(gen[4723]),
			.NE(gen[4724]),

			.O(gen[4817]),
			.E(gen[4819]),

			.SO(gen[4912]),
			.S(gen[4913]),
			.SE(gen[4914]),

			.SELF(gen[4818]),
			.cell_state(gen[4818])
		); 

/******************* CELL 4819 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4819 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4723]),
			.N(gen[4724]),
			.NE(gen[4725]),

			.O(gen[4818]),
			.E(gen[4820]),

			.SO(gen[4913]),
			.S(gen[4914]),
			.SE(gen[4915]),

			.SELF(gen[4819]),
			.cell_state(gen[4819])
		); 

/******************* CELL 4820 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4820 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4724]),
			.N(gen[4725]),
			.NE(gen[4726]),

			.O(gen[4819]),
			.E(gen[4821]),

			.SO(gen[4914]),
			.S(gen[4915]),
			.SE(gen[4916]),

			.SELF(gen[4820]),
			.cell_state(gen[4820])
		); 

/******************* CELL 4821 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4821 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4725]),
			.N(gen[4726]),
			.NE(gen[4727]),

			.O(gen[4820]),
			.E(gen[4822]),

			.SO(gen[4915]),
			.S(gen[4916]),
			.SE(gen[4917]),

			.SELF(gen[4821]),
			.cell_state(gen[4821])
		); 

/******************* CELL 4822 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4822 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4726]),
			.N(gen[4727]),
			.NE(gen[4728]),

			.O(gen[4821]),
			.E(gen[4823]),

			.SO(gen[4916]),
			.S(gen[4917]),
			.SE(gen[4918]),

			.SELF(gen[4822]),
			.cell_state(gen[4822])
		); 

/******************* CELL 4823 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4823 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4727]),
			.N(gen[4728]),
			.NE(gen[4729]),

			.O(gen[4822]),
			.E(gen[4824]),

			.SO(gen[4917]),
			.S(gen[4918]),
			.SE(gen[4919]),

			.SELF(gen[4823]),
			.cell_state(gen[4823])
		); 

/******************* CELL 4824 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4824 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4728]),
			.N(gen[4729]),
			.NE(gen[4730]),

			.O(gen[4823]),
			.E(gen[4825]),

			.SO(gen[4918]),
			.S(gen[4919]),
			.SE(gen[4920]),

			.SELF(gen[4824]),
			.cell_state(gen[4824])
		); 

/******************* CELL 4825 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4825 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4729]),
			.N(gen[4730]),
			.NE(gen[4731]),

			.O(gen[4824]),
			.E(gen[4826]),

			.SO(gen[4919]),
			.S(gen[4920]),
			.SE(gen[4921]),

			.SELF(gen[4825]),
			.cell_state(gen[4825])
		); 

/******************* CELL 4826 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4826 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4730]),
			.N(gen[4731]),
			.NE(gen[4732]),

			.O(gen[4825]),
			.E(gen[4827]),

			.SO(gen[4920]),
			.S(gen[4921]),
			.SE(gen[4922]),

			.SELF(gen[4826]),
			.cell_state(gen[4826])
		); 

/******************* CELL 4827 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4827 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4731]),
			.N(gen[4732]),
			.NE(gen[4733]),

			.O(gen[4826]),
			.E(gen[4828]),

			.SO(gen[4921]),
			.S(gen[4922]),
			.SE(gen[4923]),

			.SELF(gen[4827]),
			.cell_state(gen[4827])
		); 

/******************* CELL 4828 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4828 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4732]),
			.N(gen[4733]),
			.NE(gen[4734]),

			.O(gen[4827]),
			.E(gen[4829]),

			.SO(gen[4922]),
			.S(gen[4923]),
			.SE(gen[4924]),

			.SELF(gen[4828]),
			.cell_state(gen[4828])
		); 

/******************* CELL 4829 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4829 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4733]),
			.N(gen[4734]),
			.NE(gen[4735]),

			.O(gen[4828]),
			.E(gen[4830]),

			.SO(gen[4923]),
			.S(gen[4924]),
			.SE(gen[4925]),

			.SELF(gen[4829]),
			.cell_state(gen[4829])
		); 

/******************* CELL 4830 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4830 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4734]),
			.N(gen[4735]),
			.NE(gen[4736]),

			.O(gen[4829]),
			.E(gen[4831]),

			.SO(gen[4924]),
			.S(gen[4925]),
			.SE(gen[4926]),

			.SELF(gen[4830]),
			.cell_state(gen[4830])
		); 

/******************* CELL 4831 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4831 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4735]),
			.N(gen[4736]),
			.NE(gen[4737]),

			.O(gen[4830]),
			.E(gen[4832]),

			.SO(gen[4925]),
			.S(gen[4926]),
			.SE(gen[4927]),

			.SELF(gen[4831]),
			.cell_state(gen[4831])
		); 

/******************* CELL 4832 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4832 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4736]),
			.N(gen[4737]),
			.NE(gen[4738]),

			.O(gen[4831]),
			.E(gen[4833]),

			.SO(gen[4926]),
			.S(gen[4927]),
			.SE(gen[4928]),

			.SELF(gen[4832]),
			.cell_state(gen[4832])
		); 

/******************* CELL 4833 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4833 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4737]),
			.N(gen[4738]),
			.NE(gen[4739]),

			.O(gen[4832]),
			.E(gen[4834]),

			.SO(gen[4927]),
			.S(gen[4928]),
			.SE(gen[4929]),

			.SELF(gen[4833]),
			.cell_state(gen[4833])
		); 

/******************* CELL 4834 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4834 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4738]),
			.N(gen[4739]),
			.NE(gen[4740]),

			.O(gen[4833]),
			.E(gen[4835]),

			.SO(gen[4928]),
			.S(gen[4929]),
			.SE(gen[4930]),

			.SELF(gen[4834]),
			.cell_state(gen[4834])
		); 

/******************* CELL 4835 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4835 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4739]),
			.N(gen[4740]),
			.NE(gen[4741]),

			.O(gen[4834]),
			.E(gen[4836]),

			.SO(gen[4929]),
			.S(gen[4930]),
			.SE(gen[4931]),

			.SELF(gen[4835]),
			.cell_state(gen[4835])
		); 

/******************* CELL 4836 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4836 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4740]),
			.N(gen[4741]),
			.NE(gen[4742]),

			.O(gen[4835]),
			.E(gen[4837]),

			.SO(gen[4930]),
			.S(gen[4931]),
			.SE(gen[4932]),

			.SELF(gen[4836]),
			.cell_state(gen[4836])
		); 

/******************* CELL 4837 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4837 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4741]),
			.N(gen[4742]),
			.NE(gen[4743]),

			.O(gen[4836]),
			.E(gen[4838]),

			.SO(gen[4931]),
			.S(gen[4932]),
			.SE(gen[4933]),

			.SELF(gen[4837]),
			.cell_state(gen[4837])
		); 

/******************* CELL 4838 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4838 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4742]),
			.N(gen[4743]),
			.NE(gen[4744]),

			.O(gen[4837]),
			.E(gen[4839]),

			.SO(gen[4932]),
			.S(gen[4933]),
			.SE(gen[4934]),

			.SELF(gen[4838]),
			.cell_state(gen[4838])
		); 

/******************* CELL 4839 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4839 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4743]),
			.N(gen[4744]),
			.NE(gen[4745]),

			.O(gen[4838]),
			.E(gen[4840]),

			.SO(gen[4933]),
			.S(gen[4934]),
			.SE(gen[4935]),

			.SELF(gen[4839]),
			.cell_state(gen[4839])
		); 

/******************* CELL 4840 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4840 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4744]),
			.N(gen[4745]),
			.NE(gen[4746]),

			.O(gen[4839]),
			.E(gen[4841]),

			.SO(gen[4934]),
			.S(gen[4935]),
			.SE(gen[4936]),

			.SELF(gen[4840]),
			.cell_state(gen[4840])
		); 

/******************* CELL 4841 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4841 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4745]),
			.N(gen[4746]),
			.NE(gen[4747]),

			.O(gen[4840]),
			.E(gen[4842]),

			.SO(gen[4935]),
			.S(gen[4936]),
			.SE(gen[4937]),

			.SELF(gen[4841]),
			.cell_state(gen[4841])
		); 

/******************* CELL 4842 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4842 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4746]),
			.N(gen[4747]),
			.NE(gen[4748]),

			.O(gen[4841]),
			.E(gen[4843]),

			.SO(gen[4936]),
			.S(gen[4937]),
			.SE(gen[4938]),

			.SELF(gen[4842]),
			.cell_state(gen[4842])
		); 

/******************* CELL 4843 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4843 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4747]),
			.N(gen[4748]),
			.NE(gen[4749]),

			.O(gen[4842]),
			.E(gen[4844]),

			.SO(gen[4937]),
			.S(gen[4938]),
			.SE(gen[4939]),

			.SELF(gen[4843]),
			.cell_state(gen[4843])
		); 

/******************* CELL 4844 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4844 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4748]),
			.N(gen[4749]),
			.NE(gen[4748]),

			.O(gen[4843]),
			.E(gen[4843]),

			.SO(gen[4938]),
			.S(gen[4939]),
			.SE(gen[4938]),

			.SELF(gen[4844]),
			.cell_state(gen[4844])
		); 

/******************* CELL 4845 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4845 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4751]),
			.N(gen[4750]),
			.NE(gen[4751]),

			.O(gen[4846]),
			.E(gen[4846]),

			.SO(gen[4941]),
			.S(gen[4940]),
			.SE(gen[4941]),

			.SELF(gen[4845]),
			.cell_state(gen[4845])
		); 

/******************* CELL 4846 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4846 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4750]),
			.N(gen[4751]),
			.NE(gen[4752]),

			.O(gen[4845]),
			.E(gen[4847]),

			.SO(gen[4940]),
			.S(gen[4941]),
			.SE(gen[4942]),

			.SELF(gen[4846]),
			.cell_state(gen[4846])
		); 

/******************* CELL 4847 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4847 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4751]),
			.N(gen[4752]),
			.NE(gen[4753]),

			.O(gen[4846]),
			.E(gen[4848]),

			.SO(gen[4941]),
			.S(gen[4942]),
			.SE(gen[4943]),

			.SELF(gen[4847]),
			.cell_state(gen[4847])
		); 

/******************* CELL 4848 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4848 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4752]),
			.N(gen[4753]),
			.NE(gen[4754]),

			.O(gen[4847]),
			.E(gen[4849]),

			.SO(gen[4942]),
			.S(gen[4943]),
			.SE(gen[4944]),

			.SELF(gen[4848]),
			.cell_state(gen[4848])
		); 

/******************* CELL 4849 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4849 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4753]),
			.N(gen[4754]),
			.NE(gen[4755]),

			.O(gen[4848]),
			.E(gen[4850]),

			.SO(gen[4943]),
			.S(gen[4944]),
			.SE(gen[4945]),

			.SELF(gen[4849]),
			.cell_state(gen[4849])
		); 

/******************* CELL 4850 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4850 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4754]),
			.N(gen[4755]),
			.NE(gen[4756]),

			.O(gen[4849]),
			.E(gen[4851]),

			.SO(gen[4944]),
			.S(gen[4945]),
			.SE(gen[4946]),

			.SELF(gen[4850]),
			.cell_state(gen[4850])
		); 

/******************* CELL 4851 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4851 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4755]),
			.N(gen[4756]),
			.NE(gen[4757]),

			.O(gen[4850]),
			.E(gen[4852]),

			.SO(gen[4945]),
			.S(gen[4946]),
			.SE(gen[4947]),

			.SELF(gen[4851]),
			.cell_state(gen[4851])
		); 

/******************* CELL 4852 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4852 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4756]),
			.N(gen[4757]),
			.NE(gen[4758]),

			.O(gen[4851]),
			.E(gen[4853]),

			.SO(gen[4946]),
			.S(gen[4947]),
			.SE(gen[4948]),

			.SELF(gen[4852]),
			.cell_state(gen[4852])
		); 

/******************* CELL 4853 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4853 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4757]),
			.N(gen[4758]),
			.NE(gen[4759]),

			.O(gen[4852]),
			.E(gen[4854]),

			.SO(gen[4947]),
			.S(gen[4948]),
			.SE(gen[4949]),

			.SELF(gen[4853]),
			.cell_state(gen[4853])
		); 

/******************* CELL 4854 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4854 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4758]),
			.N(gen[4759]),
			.NE(gen[4760]),

			.O(gen[4853]),
			.E(gen[4855]),

			.SO(gen[4948]),
			.S(gen[4949]),
			.SE(gen[4950]),

			.SELF(gen[4854]),
			.cell_state(gen[4854])
		); 

/******************* CELL 4855 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4855 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4759]),
			.N(gen[4760]),
			.NE(gen[4761]),

			.O(gen[4854]),
			.E(gen[4856]),

			.SO(gen[4949]),
			.S(gen[4950]),
			.SE(gen[4951]),

			.SELF(gen[4855]),
			.cell_state(gen[4855])
		); 

/******************* CELL 4856 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4856 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4760]),
			.N(gen[4761]),
			.NE(gen[4762]),

			.O(gen[4855]),
			.E(gen[4857]),

			.SO(gen[4950]),
			.S(gen[4951]),
			.SE(gen[4952]),

			.SELF(gen[4856]),
			.cell_state(gen[4856])
		); 

/******************* CELL 4857 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4857 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4761]),
			.N(gen[4762]),
			.NE(gen[4763]),

			.O(gen[4856]),
			.E(gen[4858]),

			.SO(gen[4951]),
			.S(gen[4952]),
			.SE(gen[4953]),

			.SELF(gen[4857]),
			.cell_state(gen[4857])
		); 

/******************* CELL 4858 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4858 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4762]),
			.N(gen[4763]),
			.NE(gen[4764]),

			.O(gen[4857]),
			.E(gen[4859]),

			.SO(gen[4952]),
			.S(gen[4953]),
			.SE(gen[4954]),

			.SELF(gen[4858]),
			.cell_state(gen[4858])
		); 

/******************* CELL 4859 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4859 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4763]),
			.N(gen[4764]),
			.NE(gen[4765]),

			.O(gen[4858]),
			.E(gen[4860]),

			.SO(gen[4953]),
			.S(gen[4954]),
			.SE(gen[4955]),

			.SELF(gen[4859]),
			.cell_state(gen[4859])
		); 

/******************* CELL 4860 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4860 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4764]),
			.N(gen[4765]),
			.NE(gen[4766]),

			.O(gen[4859]),
			.E(gen[4861]),

			.SO(gen[4954]),
			.S(gen[4955]),
			.SE(gen[4956]),

			.SELF(gen[4860]),
			.cell_state(gen[4860])
		); 

/******************* CELL 4861 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4861 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4765]),
			.N(gen[4766]),
			.NE(gen[4767]),

			.O(gen[4860]),
			.E(gen[4862]),

			.SO(gen[4955]),
			.S(gen[4956]),
			.SE(gen[4957]),

			.SELF(gen[4861]),
			.cell_state(gen[4861])
		); 

/******************* CELL 4862 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4862 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4766]),
			.N(gen[4767]),
			.NE(gen[4768]),

			.O(gen[4861]),
			.E(gen[4863]),

			.SO(gen[4956]),
			.S(gen[4957]),
			.SE(gen[4958]),

			.SELF(gen[4862]),
			.cell_state(gen[4862])
		); 

/******************* CELL 4863 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4863 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4767]),
			.N(gen[4768]),
			.NE(gen[4769]),

			.O(gen[4862]),
			.E(gen[4864]),

			.SO(gen[4957]),
			.S(gen[4958]),
			.SE(gen[4959]),

			.SELF(gen[4863]),
			.cell_state(gen[4863])
		); 

/******************* CELL 4864 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4864 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4768]),
			.N(gen[4769]),
			.NE(gen[4770]),

			.O(gen[4863]),
			.E(gen[4865]),

			.SO(gen[4958]),
			.S(gen[4959]),
			.SE(gen[4960]),

			.SELF(gen[4864]),
			.cell_state(gen[4864])
		); 

/******************* CELL 4865 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4865 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4769]),
			.N(gen[4770]),
			.NE(gen[4771]),

			.O(gen[4864]),
			.E(gen[4866]),

			.SO(gen[4959]),
			.S(gen[4960]),
			.SE(gen[4961]),

			.SELF(gen[4865]),
			.cell_state(gen[4865])
		); 

/******************* CELL 4866 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4866 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4770]),
			.N(gen[4771]),
			.NE(gen[4772]),

			.O(gen[4865]),
			.E(gen[4867]),

			.SO(gen[4960]),
			.S(gen[4961]),
			.SE(gen[4962]),

			.SELF(gen[4866]),
			.cell_state(gen[4866])
		); 

/******************* CELL 4867 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4867 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4771]),
			.N(gen[4772]),
			.NE(gen[4773]),

			.O(gen[4866]),
			.E(gen[4868]),

			.SO(gen[4961]),
			.S(gen[4962]),
			.SE(gen[4963]),

			.SELF(gen[4867]),
			.cell_state(gen[4867])
		); 

/******************* CELL 4868 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4868 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4772]),
			.N(gen[4773]),
			.NE(gen[4774]),

			.O(gen[4867]),
			.E(gen[4869]),

			.SO(gen[4962]),
			.S(gen[4963]),
			.SE(gen[4964]),

			.SELF(gen[4868]),
			.cell_state(gen[4868])
		); 

/******************* CELL 4869 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4869 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4773]),
			.N(gen[4774]),
			.NE(gen[4775]),

			.O(gen[4868]),
			.E(gen[4870]),

			.SO(gen[4963]),
			.S(gen[4964]),
			.SE(gen[4965]),

			.SELF(gen[4869]),
			.cell_state(gen[4869])
		); 

/******************* CELL 4870 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4870 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4774]),
			.N(gen[4775]),
			.NE(gen[4776]),

			.O(gen[4869]),
			.E(gen[4871]),

			.SO(gen[4964]),
			.S(gen[4965]),
			.SE(gen[4966]),

			.SELF(gen[4870]),
			.cell_state(gen[4870])
		); 

/******************* CELL 4871 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4871 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4775]),
			.N(gen[4776]),
			.NE(gen[4777]),

			.O(gen[4870]),
			.E(gen[4872]),

			.SO(gen[4965]),
			.S(gen[4966]),
			.SE(gen[4967]),

			.SELF(gen[4871]),
			.cell_state(gen[4871])
		); 

/******************* CELL 4872 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4872 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4776]),
			.N(gen[4777]),
			.NE(gen[4778]),

			.O(gen[4871]),
			.E(gen[4873]),

			.SO(gen[4966]),
			.S(gen[4967]),
			.SE(gen[4968]),

			.SELF(gen[4872]),
			.cell_state(gen[4872])
		); 

/******************* CELL 4873 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4873 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4777]),
			.N(gen[4778]),
			.NE(gen[4779]),

			.O(gen[4872]),
			.E(gen[4874]),

			.SO(gen[4967]),
			.S(gen[4968]),
			.SE(gen[4969]),

			.SELF(gen[4873]),
			.cell_state(gen[4873])
		); 

/******************* CELL 4874 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4874 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4778]),
			.N(gen[4779]),
			.NE(gen[4780]),

			.O(gen[4873]),
			.E(gen[4875]),

			.SO(gen[4968]),
			.S(gen[4969]),
			.SE(gen[4970]),

			.SELF(gen[4874]),
			.cell_state(gen[4874])
		); 

/******************* CELL 4875 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4875 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4779]),
			.N(gen[4780]),
			.NE(gen[4781]),

			.O(gen[4874]),
			.E(gen[4876]),

			.SO(gen[4969]),
			.S(gen[4970]),
			.SE(gen[4971]),

			.SELF(gen[4875]),
			.cell_state(gen[4875])
		); 

/******************* CELL 4876 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4876 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4780]),
			.N(gen[4781]),
			.NE(gen[4782]),

			.O(gen[4875]),
			.E(gen[4877]),

			.SO(gen[4970]),
			.S(gen[4971]),
			.SE(gen[4972]),

			.SELF(gen[4876]),
			.cell_state(gen[4876])
		); 

/******************* CELL 4877 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4877 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4781]),
			.N(gen[4782]),
			.NE(gen[4783]),

			.O(gen[4876]),
			.E(gen[4878]),

			.SO(gen[4971]),
			.S(gen[4972]),
			.SE(gen[4973]),

			.SELF(gen[4877]),
			.cell_state(gen[4877])
		); 

/******************* CELL 4878 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4878 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4782]),
			.N(gen[4783]),
			.NE(gen[4784]),

			.O(gen[4877]),
			.E(gen[4879]),

			.SO(gen[4972]),
			.S(gen[4973]),
			.SE(gen[4974]),

			.SELF(gen[4878]),
			.cell_state(gen[4878])
		); 

/******************* CELL 4879 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4879 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4783]),
			.N(gen[4784]),
			.NE(gen[4785]),

			.O(gen[4878]),
			.E(gen[4880]),

			.SO(gen[4973]),
			.S(gen[4974]),
			.SE(gen[4975]),

			.SELF(gen[4879]),
			.cell_state(gen[4879])
		); 

/******************* CELL 4880 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4880 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4784]),
			.N(gen[4785]),
			.NE(gen[4786]),

			.O(gen[4879]),
			.E(gen[4881]),

			.SO(gen[4974]),
			.S(gen[4975]),
			.SE(gen[4976]),

			.SELF(gen[4880]),
			.cell_state(gen[4880])
		); 

/******************* CELL 4881 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4881 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4785]),
			.N(gen[4786]),
			.NE(gen[4787]),

			.O(gen[4880]),
			.E(gen[4882]),

			.SO(gen[4975]),
			.S(gen[4976]),
			.SE(gen[4977]),

			.SELF(gen[4881]),
			.cell_state(gen[4881])
		); 

/******************* CELL 4882 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4882 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4786]),
			.N(gen[4787]),
			.NE(gen[4788]),

			.O(gen[4881]),
			.E(gen[4883]),

			.SO(gen[4976]),
			.S(gen[4977]),
			.SE(gen[4978]),

			.SELF(gen[4882]),
			.cell_state(gen[4882])
		); 

/******************* CELL 4883 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4883 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4787]),
			.N(gen[4788]),
			.NE(gen[4789]),

			.O(gen[4882]),
			.E(gen[4884]),

			.SO(gen[4977]),
			.S(gen[4978]),
			.SE(gen[4979]),

			.SELF(gen[4883]),
			.cell_state(gen[4883])
		); 

/******************* CELL 4884 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4884 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4788]),
			.N(gen[4789]),
			.NE(gen[4790]),

			.O(gen[4883]),
			.E(gen[4885]),

			.SO(gen[4978]),
			.S(gen[4979]),
			.SE(gen[4980]),

			.SELF(gen[4884]),
			.cell_state(gen[4884])
		); 

/******************* CELL 4885 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4885 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4789]),
			.N(gen[4790]),
			.NE(gen[4791]),

			.O(gen[4884]),
			.E(gen[4886]),

			.SO(gen[4979]),
			.S(gen[4980]),
			.SE(gen[4981]),

			.SELF(gen[4885]),
			.cell_state(gen[4885])
		); 

/******************* CELL 4886 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4886 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4790]),
			.N(gen[4791]),
			.NE(gen[4792]),

			.O(gen[4885]),
			.E(gen[4887]),

			.SO(gen[4980]),
			.S(gen[4981]),
			.SE(gen[4982]),

			.SELF(gen[4886]),
			.cell_state(gen[4886])
		); 

/******************* CELL 4887 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4887 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4791]),
			.N(gen[4792]),
			.NE(gen[4793]),

			.O(gen[4886]),
			.E(gen[4888]),

			.SO(gen[4981]),
			.S(gen[4982]),
			.SE(gen[4983]),

			.SELF(gen[4887]),
			.cell_state(gen[4887])
		); 

/******************* CELL 4888 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4888 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4792]),
			.N(gen[4793]),
			.NE(gen[4794]),

			.O(gen[4887]),
			.E(gen[4889]),

			.SO(gen[4982]),
			.S(gen[4983]),
			.SE(gen[4984]),

			.SELF(gen[4888]),
			.cell_state(gen[4888])
		); 

/******************* CELL 4889 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4889 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4793]),
			.N(gen[4794]),
			.NE(gen[4795]),

			.O(gen[4888]),
			.E(gen[4890]),

			.SO(gen[4983]),
			.S(gen[4984]),
			.SE(gen[4985]),

			.SELF(gen[4889]),
			.cell_state(gen[4889])
		); 

/******************* CELL 4890 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4890 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4794]),
			.N(gen[4795]),
			.NE(gen[4796]),

			.O(gen[4889]),
			.E(gen[4891]),

			.SO(gen[4984]),
			.S(gen[4985]),
			.SE(gen[4986]),

			.SELF(gen[4890]),
			.cell_state(gen[4890])
		); 

/******************* CELL 4891 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4891 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4795]),
			.N(gen[4796]),
			.NE(gen[4797]),

			.O(gen[4890]),
			.E(gen[4892]),

			.SO(gen[4985]),
			.S(gen[4986]),
			.SE(gen[4987]),

			.SELF(gen[4891]),
			.cell_state(gen[4891])
		); 

/******************* CELL 4892 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4892 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4796]),
			.N(gen[4797]),
			.NE(gen[4798]),

			.O(gen[4891]),
			.E(gen[4893]),

			.SO(gen[4986]),
			.S(gen[4987]),
			.SE(gen[4988]),

			.SELF(gen[4892]),
			.cell_state(gen[4892])
		); 

/******************* CELL 4893 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4893 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4797]),
			.N(gen[4798]),
			.NE(gen[4799]),

			.O(gen[4892]),
			.E(gen[4894]),

			.SO(gen[4987]),
			.S(gen[4988]),
			.SE(gen[4989]),

			.SELF(gen[4893]),
			.cell_state(gen[4893])
		); 

/******************* CELL 4894 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4894 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4798]),
			.N(gen[4799]),
			.NE(gen[4800]),

			.O(gen[4893]),
			.E(gen[4895]),

			.SO(gen[4988]),
			.S(gen[4989]),
			.SE(gen[4990]),

			.SELF(gen[4894]),
			.cell_state(gen[4894])
		); 

/******************* CELL 4895 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4895 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4799]),
			.N(gen[4800]),
			.NE(gen[4801]),

			.O(gen[4894]),
			.E(gen[4896]),

			.SO(gen[4989]),
			.S(gen[4990]),
			.SE(gen[4991]),

			.SELF(gen[4895]),
			.cell_state(gen[4895])
		); 

/******************* CELL 4896 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4896 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4800]),
			.N(gen[4801]),
			.NE(gen[4802]),

			.O(gen[4895]),
			.E(gen[4897]),

			.SO(gen[4990]),
			.S(gen[4991]),
			.SE(gen[4992]),

			.SELF(gen[4896]),
			.cell_state(gen[4896])
		); 

/******************* CELL 4897 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4897 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4801]),
			.N(gen[4802]),
			.NE(gen[4803]),

			.O(gen[4896]),
			.E(gen[4898]),

			.SO(gen[4991]),
			.S(gen[4992]),
			.SE(gen[4993]),

			.SELF(gen[4897]),
			.cell_state(gen[4897])
		); 

/******************* CELL 4898 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4898 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4802]),
			.N(gen[4803]),
			.NE(gen[4804]),

			.O(gen[4897]),
			.E(gen[4899]),

			.SO(gen[4992]),
			.S(gen[4993]),
			.SE(gen[4994]),

			.SELF(gen[4898]),
			.cell_state(gen[4898])
		); 

/******************* CELL 4899 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4899 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4803]),
			.N(gen[4804]),
			.NE(gen[4805]),

			.O(gen[4898]),
			.E(gen[4900]),

			.SO(gen[4993]),
			.S(gen[4994]),
			.SE(gen[4995]),

			.SELF(gen[4899]),
			.cell_state(gen[4899])
		); 

/******************* CELL 4900 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4900 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4804]),
			.N(gen[4805]),
			.NE(gen[4806]),

			.O(gen[4899]),
			.E(gen[4901]),

			.SO(gen[4994]),
			.S(gen[4995]),
			.SE(gen[4996]),

			.SELF(gen[4900]),
			.cell_state(gen[4900])
		); 

/******************* CELL 4901 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4901 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4805]),
			.N(gen[4806]),
			.NE(gen[4807]),

			.O(gen[4900]),
			.E(gen[4902]),

			.SO(gen[4995]),
			.S(gen[4996]),
			.SE(gen[4997]),

			.SELF(gen[4901]),
			.cell_state(gen[4901])
		); 

/******************* CELL 4902 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4902 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4806]),
			.N(gen[4807]),
			.NE(gen[4808]),

			.O(gen[4901]),
			.E(gen[4903]),

			.SO(gen[4996]),
			.S(gen[4997]),
			.SE(gen[4998]),

			.SELF(gen[4902]),
			.cell_state(gen[4902])
		); 

/******************* CELL 4903 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4903 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4807]),
			.N(gen[4808]),
			.NE(gen[4809]),

			.O(gen[4902]),
			.E(gen[4904]),

			.SO(gen[4997]),
			.S(gen[4998]),
			.SE(gen[4999]),

			.SELF(gen[4903]),
			.cell_state(gen[4903])
		); 

/******************* CELL 4904 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4904 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4808]),
			.N(gen[4809]),
			.NE(gen[4810]),

			.O(gen[4903]),
			.E(gen[4905]),

			.SO(gen[4998]),
			.S(gen[4999]),
			.SE(gen[5000]),

			.SELF(gen[4904]),
			.cell_state(gen[4904])
		); 

/******************* CELL 4905 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4905 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4809]),
			.N(gen[4810]),
			.NE(gen[4811]),

			.O(gen[4904]),
			.E(gen[4906]),

			.SO(gen[4999]),
			.S(gen[5000]),
			.SE(gen[5001]),

			.SELF(gen[4905]),
			.cell_state(gen[4905])
		); 

/******************* CELL 4906 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4906 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4810]),
			.N(gen[4811]),
			.NE(gen[4812]),

			.O(gen[4905]),
			.E(gen[4907]),

			.SO(gen[5000]),
			.S(gen[5001]),
			.SE(gen[5002]),

			.SELF(gen[4906]),
			.cell_state(gen[4906])
		); 

/******************* CELL 4907 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4907 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4811]),
			.N(gen[4812]),
			.NE(gen[4813]),

			.O(gen[4906]),
			.E(gen[4908]),

			.SO(gen[5001]),
			.S(gen[5002]),
			.SE(gen[5003]),

			.SELF(gen[4907]),
			.cell_state(gen[4907])
		); 

/******************* CELL 4908 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4908 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4812]),
			.N(gen[4813]),
			.NE(gen[4814]),

			.O(gen[4907]),
			.E(gen[4909]),

			.SO(gen[5002]),
			.S(gen[5003]),
			.SE(gen[5004]),

			.SELF(gen[4908]),
			.cell_state(gen[4908])
		); 

/******************* CELL 4909 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4909 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4813]),
			.N(gen[4814]),
			.NE(gen[4815]),

			.O(gen[4908]),
			.E(gen[4910]),

			.SO(gen[5003]),
			.S(gen[5004]),
			.SE(gen[5005]),

			.SELF(gen[4909]),
			.cell_state(gen[4909])
		); 

/******************* CELL 4910 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4910 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4814]),
			.N(gen[4815]),
			.NE(gen[4816]),

			.O(gen[4909]),
			.E(gen[4911]),

			.SO(gen[5004]),
			.S(gen[5005]),
			.SE(gen[5006]),

			.SELF(gen[4910]),
			.cell_state(gen[4910])
		); 

/******************* CELL 4911 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4911 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4815]),
			.N(gen[4816]),
			.NE(gen[4817]),

			.O(gen[4910]),
			.E(gen[4912]),

			.SO(gen[5005]),
			.S(gen[5006]),
			.SE(gen[5007]),

			.SELF(gen[4911]),
			.cell_state(gen[4911])
		); 

/******************* CELL 4912 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4912 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4816]),
			.N(gen[4817]),
			.NE(gen[4818]),

			.O(gen[4911]),
			.E(gen[4913]),

			.SO(gen[5006]),
			.S(gen[5007]),
			.SE(gen[5008]),

			.SELF(gen[4912]),
			.cell_state(gen[4912])
		); 

/******************* CELL 4913 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4913 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4817]),
			.N(gen[4818]),
			.NE(gen[4819]),

			.O(gen[4912]),
			.E(gen[4914]),

			.SO(gen[5007]),
			.S(gen[5008]),
			.SE(gen[5009]),

			.SELF(gen[4913]),
			.cell_state(gen[4913])
		); 

/******************* CELL 4914 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4914 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4818]),
			.N(gen[4819]),
			.NE(gen[4820]),

			.O(gen[4913]),
			.E(gen[4915]),

			.SO(gen[5008]),
			.S(gen[5009]),
			.SE(gen[5010]),

			.SELF(gen[4914]),
			.cell_state(gen[4914])
		); 

/******************* CELL 4915 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4915 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4819]),
			.N(gen[4820]),
			.NE(gen[4821]),

			.O(gen[4914]),
			.E(gen[4916]),

			.SO(gen[5009]),
			.S(gen[5010]),
			.SE(gen[5011]),

			.SELF(gen[4915]),
			.cell_state(gen[4915])
		); 

/******************* CELL 4916 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4916 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4820]),
			.N(gen[4821]),
			.NE(gen[4822]),

			.O(gen[4915]),
			.E(gen[4917]),

			.SO(gen[5010]),
			.S(gen[5011]),
			.SE(gen[5012]),

			.SELF(gen[4916]),
			.cell_state(gen[4916])
		); 

/******************* CELL 4917 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4917 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4821]),
			.N(gen[4822]),
			.NE(gen[4823]),

			.O(gen[4916]),
			.E(gen[4918]),

			.SO(gen[5011]),
			.S(gen[5012]),
			.SE(gen[5013]),

			.SELF(gen[4917]),
			.cell_state(gen[4917])
		); 

/******************* CELL 4918 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4918 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4822]),
			.N(gen[4823]),
			.NE(gen[4824]),

			.O(gen[4917]),
			.E(gen[4919]),

			.SO(gen[5012]),
			.S(gen[5013]),
			.SE(gen[5014]),

			.SELF(gen[4918]),
			.cell_state(gen[4918])
		); 

/******************* CELL 4919 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4919 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4823]),
			.N(gen[4824]),
			.NE(gen[4825]),

			.O(gen[4918]),
			.E(gen[4920]),

			.SO(gen[5013]),
			.S(gen[5014]),
			.SE(gen[5015]),

			.SELF(gen[4919]),
			.cell_state(gen[4919])
		); 

/******************* CELL 4920 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4920 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4824]),
			.N(gen[4825]),
			.NE(gen[4826]),

			.O(gen[4919]),
			.E(gen[4921]),

			.SO(gen[5014]),
			.S(gen[5015]),
			.SE(gen[5016]),

			.SELF(gen[4920]),
			.cell_state(gen[4920])
		); 

/******************* CELL 4921 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4921 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4825]),
			.N(gen[4826]),
			.NE(gen[4827]),

			.O(gen[4920]),
			.E(gen[4922]),

			.SO(gen[5015]),
			.S(gen[5016]),
			.SE(gen[5017]),

			.SELF(gen[4921]),
			.cell_state(gen[4921])
		); 

/******************* CELL 4922 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4922 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4826]),
			.N(gen[4827]),
			.NE(gen[4828]),

			.O(gen[4921]),
			.E(gen[4923]),

			.SO(gen[5016]),
			.S(gen[5017]),
			.SE(gen[5018]),

			.SELF(gen[4922]),
			.cell_state(gen[4922])
		); 

/******************* CELL 4923 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4923 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4827]),
			.N(gen[4828]),
			.NE(gen[4829]),

			.O(gen[4922]),
			.E(gen[4924]),

			.SO(gen[5017]),
			.S(gen[5018]),
			.SE(gen[5019]),

			.SELF(gen[4923]),
			.cell_state(gen[4923])
		); 

/******************* CELL 4924 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4924 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4828]),
			.N(gen[4829]),
			.NE(gen[4830]),

			.O(gen[4923]),
			.E(gen[4925]),

			.SO(gen[5018]),
			.S(gen[5019]),
			.SE(gen[5020]),

			.SELF(gen[4924]),
			.cell_state(gen[4924])
		); 

/******************* CELL 4925 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4925 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4829]),
			.N(gen[4830]),
			.NE(gen[4831]),

			.O(gen[4924]),
			.E(gen[4926]),

			.SO(gen[5019]),
			.S(gen[5020]),
			.SE(gen[5021]),

			.SELF(gen[4925]),
			.cell_state(gen[4925])
		); 

/******************* CELL 4926 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4926 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4830]),
			.N(gen[4831]),
			.NE(gen[4832]),

			.O(gen[4925]),
			.E(gen[4927]),

			.SO(gen[5020]),
			.S(gen[5021]),
			.SE(gen[5022]),

			.SELF(gen[4926]),
			.cell_state(gen[4926])
		); 

/******************* CELL 4927 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4927 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4831]),
			.N(gen[4832]),
			.NE(gen[4833]),

			.O(gen[4926]),
			.E(gen[4928]),

			.SO(gen[5021]),
			.S(gen[5022]),
			.SE(gen[5023]),

			.SELF(gen[4927]),
			.cell_state(gen[4927])
		); 

/******************* CELL 4928 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4928 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4832]),
			.N(gen[4833]),
			.NE(gen[4834]),

			.O(gen[4927]),
			.E(gen[4929]),

			.SO(gen[5022]),
			.S(gen[5023]),
			.SE(gen[5024]),

			.SELF(gen[4928]),
			.cell_state(gen[4928])
		); 

/******************* CELL 4929 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4929 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4833]),
			.N(gen[4834]),
			.NE(gen[4835]),

			.O(gen[4928]),
			.E(gen[4930]),

			.SO(gen[5023]),
			.S(gen[5024]),
			.SE(gen[5025]),

			.SELF(gen[4929]),
			.cell_state(gen[4929])
		); 

/******************* CELL 4930 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4930 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4834]),
			.N(gen[4835]),
			.NE(gen[4836]),

			.O(gen[4929]),
			.E(gen[4931]),

			.SO(gen[5024]),
			.S(gen[5025]),
			.SE(gen[5026]),

			.SELF(gen[4930]),
			.cell_state(gen[4930])
		); 

/******************* CELL 4931 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4931 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4835]),
			.N(gen[4836]),
			.NE(gen[4837]),

			.O(gen[4930]),
			.E(gen[4932]),

			.SO(gen[5025]),
			.S(gen[5026]),
			.SE(gen[5027]),

			.SELF(gen[4931]),
			.cell_state(gen[4931])
		); 

/******************* CELL 4932 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4932 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4836]),
			.N(gen[4837]),
			.NE(gen[4838]),

			.O(gen[4931]),
			.E(gen[4933]),

			.SO(gen[5026]),
			.S(gen[5027]),
			.SE(gen[5028]),

			.SELF(gen[4932]),
			.cell_state(gen[4932])
		); 

/******************* CELL 4933 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4933 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4837]),
			.N(gen[4838]),
			.NE(gen[4839]),

			.O(gen[4932]),
			.E(gen[4934]),

			.SO(gen[5027]),
			.S(gen[5028]),
			.SE(gen[5029]),

			.SELF(gen[4933]),
			.cell_state(gen[4933])
		); 

/******************* CELL 4934 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4934 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4838]),
			.N(gen[4839]),
			.NE(gen[4840]),

			.O(gen[4933]),
			.E(gen[4935]),

			.SO(gen[5028]),
			.S(gen[5029]),
			.SE(gen[5030]),

			.SELF(gen[4934]),
			.cell_state(gen[4934])
		); 

/******************* CELL 4935 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4935 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4839]),
			.N(gen[4840]),
			.NE(gen[4841]),

			.O(gen[4934]),
			.E(gen[4936]),

			.SO(gen[5029]),
			.S(gen[5030]),
			.SE(gen[5031]),

			.SELF(gen[4935]),
			.cell_state(gen[4935])
		); 

/******************* CELL 4936 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4936 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4840]),
			.N(gen[4841]),
			.NE(gen[4842]),

			.O(gen[4935]),
			.E(gen[4937]),

			.SO(gen[5030]),
			.S(gen[5031]),
			.SE(gen[5032]),

			.SELF(gen[4936]),
			.cell_state(gen[4936])
		); 

/******************* CELL 4937 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4937 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4841]),
			.N(gen[4842]),
			.NE(gen[4843]),

			.O(gen[4936]),
			.E(gen[4938]),

			.SO(gen[5031]),
			.S(gen[5032]),
			.SE(gen[5033]),

			.SELF(gen[4937]),
			.cell_state(gen[4937])
		); 

/******************* CELL 4938 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4938 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4842]),
			.N(gen[4843]),
			.NE(gen[4844]),

			.O(gen[4937]),
			.E(gen[4939]),

			.SO(gen[5032]),
			.S(gen[5033]),
			.SE(gen[5034]),

			.SELF(gen[4938]),
			.cell_state(gen[4938])
		); 

/******************* CELL 4939 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4939 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4843]),
			.N(gen[4844]),
			.NE(gen[4843]),

			.O(gen[4938]),
			.E(gen[4938]),

			.SO(gen[5033]),
			.S(gen[5034]),
			.SE(gen[5033]),

			.SELF(gen[4939]),
			.cell_state(gen[4939])
		); 

/******************* CELL 4940 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4940 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4846]),
			.N(gen[4845]),
			.NE(gen[4846]),

			.O(gen[4941]),
			.E(gen[4941]),

			.SO(gen[5036]),
			.S(gen[5035]),
			.SE(gen[5036]),

			.SELF(gen[4940]),
			.cell_state(gen[4940])
		); 

/******************* CELL 4941 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4941 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4845]),
			.N(gen[4846]),
			.NE(gen[4847]),

			.O(gen[4940]),
			.E(gen[4942]),

			.SO(gen[5035]),
			.S(gen[5036]),
			.SE(gen[5037]),

			.SELF(gen[4941]),
			.cell_state(gen[4941])
		); 

/******************* CELL 4942 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4942 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4846]),
			.N(gen[4847]),
			.NE(gen[4848]),

			.O(gen[4941]),
			.E(gen[4943]),

			.SO(gen[5036]),
			.S(gen[5037]),
			.SE(gen[5038]),

			.SELF(gen[4942]),
			.cell_state(gen[4942])
		); 

/******************* CELL 4943 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4943 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4847]),
			.N(gen[4848]),
			.NE(gen[4849]),

			.O(gen[4942]),
			.E(gen[4944]),

			.SO(gen[5037]),
			.S(gen[5038]),
			.SE(gen[5039]),

			.SELF(gen[4943]),
			.cell_state(gen[4943])
		); 

/******************* CELL 4944 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4944 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4848]),
			.N(gen[4849]),
			.NE(gen[4850]),

			.O(gen[4943]),
			.E(gen[4945]),

			.SO(gen[5038]),
			.S(gen[5039]),
			.SE(gen[5040]),

			.SELF(gen[4944]),
			.cell_state(gen[4944])
		); 

/******************* CELL 4945 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4945 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4849]),
			.N(gen[4850]),
			.NE(gen[4851]),

			.O(gen[4944]),
			.E(gen[4946]),

			.SO(gen[5039]),
			.S(gen[5040]),
			.SE(gen[5041]),

			.SELF(gen[4945]),
			.cell_state(gen[4945])
		); 

/******************* CELL 4946 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4946 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4850]),
			.N(gen[4851]),
			.NE(gen[4852]),

			.O(gen[4945]),
			.E(gen[4947]),

			.SO(gen[5040]),
			.S(gen[5041]),
			.SE(gen[5042]),

			.SELF(gen[4946]),
			.cell_state(gen[4946])
		); 

/******************* CELL 4947 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4947 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4851]),
			.N(gen[4852]),
			.NE(gen[4853]),

			.O(gen[4946]),
			.E(gen[4948]),

			.SO(gen[5041]),
			.S(gen[5042]),
			.SE(gen[5043]),

			.SELF(gen[4947]),
			.cell_state(gen[4947])
		); 

/******************* CELL 4948 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4948 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4852]),
			.N(gen[4853]),
			.NE(gen[4854]),

			.O(gen[4947]),
			.E(gen[4949]),

			.SO(gen[5042]),
			.S(gen[5043]),
			.SE(gen[5044]),

			.SELF(gen[4948]),
			.cell_state(gen[4948])
		); 

/******************* CELL 4949 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4949 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4853]),
			.N(gen[4854]),
			.NE(gen[4855]),

			.O(gen[4948]),
			.E(gen[4950]),

			.SO(gen[5043]),
			.S(gen[5044]),
			.SE(gen[5045]),

			.SELF(gen[4949]),
			.cell_state(gen[4949])
		); 

/******************* CELL 4950 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4950 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4854]),
			.N(gen[4855]),
			.NE(gen[4856]),

			.O(gen[4949]),
			.E(gen[4951]),

			.SO(gen[5044]),
			.S(gen[5045]),
			.SE(gen[5046]),

			.SELF(gen[4950]),
			.cell_state(gen[4950])
		); 

/******************* CELL 4951 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4951 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4855]),
			.N(gen[4856]),
			.NE(gen[4857]),

			.O(gen[4950]),
			.E(gen[4952]),

			.SO(gen[5045]),
			.S(gen[5046]),
			.SE(gen[5047]),

			.SELF(gen[4951]),
			.cell_state(gen[4951])
		); 

/******************* CELL 4952 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4952 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4856]),
			.N(gen[4857]),
			.NE(gen[4858]),

			.O(gen[4951]),
			.E(gen[4953]),

			.SO(gen[5046]),
			.S(gen[5047]),
			.SE(gen[5048]),

			.SELF(gen[4952]),
			.cell_state(gen[4952])
		); 

/******************* CELL 4953 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4953 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4857]),
			.N(gen[4858]),
			.NE(gen[4859]),

			.O(gen[4952]),
			.E(gen[4954]),

			.SO(gen[5047]),
			.S(gen[5048]),
			.SE(gen[5049]),

			.SELF(gen[4953]),
			.cell_state(gen[4953])
		); 

/******************* CELL 4954 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4954 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4858]),
			.N(gen[4859]),
			.NE(gen[4860]),

			.O(gen[4953]),
			.E(gen[4955]),

			.SO(gen[5048]),
			.S(gen[5049]),
			.SE(gen[5050]),

			.SELF(gen[4954]),
			.cell_state(gen[4954])
		); 

/******************* CELL 4955 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4955 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4859]),
			.N(gen[4860]),
			.NE(gen[4861]),

			.O(gen[4954]),
			.E(gen[4956]),

			.SO(gen[5049]),
			.S(gen[5050]),
			.SE(gen[5051]),

			.SELF(gen[4955]),
			.cell_state(gen[4955])
		); 

/******************* CELL 4956 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4956 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4860]),
			.N(gen[4861]),
			.NE(gen[4862]),

			.O(gen[4955]),
			.E(gen[4957]),

			.SO(gen[5050]),
			.S(gen[5051]),
			.SE(gen[5052]),

			.SELF(gen[4956]),
			.cell_state(gen[4956])
		); 

/******************* CELL 4957 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4957 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4861]),
			.N(gen[4862]),
			.NE(gen[4863]),

			.O(gen[4956]),
			.E(gen[4958]),

			.SO(gen[5051]),
			.S(gen[5052]),
			.SE(gen[5053]),

			.SELF(gen[4957]),
			.cell_state(gen[4957])
		); 

/******************* CELL 4958 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4958 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4862]),
			.N(gen[4863]),
			.NE(gen[4864]),

			.O(gen[4957]),
			.E(gen[4959]),

			.SO(gen[5052]),
			.S(gen[5053]),
			.SE(gen[5054]),

			.SELF(gen[4958]),
			.cell_state(gen[4958])
		); 

/******************* CELL 4959 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4959 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4863]),
			.N(gen[4864]),
			.NE(gen[4865]),

			.O(gen[4958]),
			.E(gen[4960]),

			.SO(gen[5053]),
			.S(gen[5054]),
			.SE(gen[5055]),

			.SELF(gen[4959]),
			.cell_state(gen[4959])
		); 

/******************* CELL 4960 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4960 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4864]),
			.N(gen[4865]),
			.NE(gen[4866]),

			.O(gen[4959]),
			.E(gen[4961]),

			.SO(gen[5054]),
			.S(gen[5055]),
			.SE(gen[5056]),

			.SELF(gen[4960]),
			.cell_state(gen[4960])
		); 

/******************* CELL 4961 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4961 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4865]),
			.N(gen[4866]),
			.NE(gen[4867]),

			.O(gen[4960]),
			.E(gen[4962]),

			.SO(gen[5055]),
			.S(gen[5056]),
			.SE(gen[5057]),

			.SELF(gen[4961]),
			.cell_state(gen[4961])
		); 

/******************* CELL 4962 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4962 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4866]),
			.N(gen[4867]),
			.NE(gen[4868]),

			.O(gen[4961]),
			.E(gen[4963]),

			.SO(gen[5056]),
			.S(gen[5057]),
			.SE(gen[5058]),

			.SELF(gen[4962]),
			.cell_state(gen[4962])
		); 

/******************* CELL 4963 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4963 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4867]),
			.N(gen[4868]),
			.NE(gen[4869]),

			.O(gen[4962]),
			.E(gen[4964]),

			.SO(gen[5057]),
			.S(gen[5058]),
			.SE(gen[5059]),

			.SELF(gen[4963]),
			.cell_state(gen[4963])
		); 

/******************* CELL 4964 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4964 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4868]),
			.N(gen[4869]),
			.NE(gen[4870]),

			.O(gen[4963]),
			.E(gen[4965]),

			.SO(gen[5058]),
			.S(gen[5059]),
			.SE(gen[5060]),

			.SELF(gen[4964]),
			.cell_state(gen[4964])
		); 

/******************* CELL 4965 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4965 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4869]),
			.N(gen[4870]),
			.NE(gen[4871]),

			.O(gen[4964]),
			.E(gen[4966]),

			.SO(gen[5059]),
			.S(gen[5060]),
			.SE(gen[5061]),

			.SELF(gen[4965]),
			.cell_state(gen[4965])
		); 

/******************* CELL 4966 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4966 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4870]),
			.N(gen[4871]),
			.NE(gen[4872]),

			.O(gen[4965]),
			.E(gen[4967]),

			.SO(gen[5060]),
			.S(gen[5061]),
			.SE(gen[5062]),

			.SELF(gen[4966]),
			.cell_state(gen[4966])
		); 

/******************* CELL 4967 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4967 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4871]),
			.N(gen[4872]),
			.NE(gen[4873]),

			.O(gen[4966]),
			.E(gen[4968]),

			.SO(gen[5061]),
			.S(gen[5062]),
			.SE(gen[5063]),

			.SELF(gen[4967]),
			.cell_state(gen[4967])
		); 

/******************* CELL 4968 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4968 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4872]),
			.N(gen[4873]),
			.NE(gen[4874]),

			.O(gen[4967]),
			.E(gen[4969]),

			.SO(gen[5062]),
			.S(gen[5063]),
			.SE(gen[5064]),

			.SELF(gen[4968]),
			.cell_state(gen[4968])
		); 

/******************* CELL 4969 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4969 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4873]),
			.N(gen[4874]),
			.NE(gen[4875]),

			.O(gen[4968]),
			.E(gen[4970]),

			.SO(gen[5063]),
			.S(gen[5064]),
			.SE(gen[5065]),

			.SELF(gen[4969]),
			.cell_state(gen[4969])
		); 

/******************* CELL 4970 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4970 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4874]),
			.N(gen[4875]),
			.NE(gen[4876]),

			.O(gen[4969]),
			.E(gen[4971]),

			.SO(gen[5064]),
			.S(gen[5065]),
			.SE(gen[5066]),

			.SELF(gen[4970]),
			.cell_state(gen[4970])
		); 

/******************* CELL 4971 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4971 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4875]),
			.N(gen[4876]),
			.NE(gen[4877]),

			.O(gen[4970]),
			.E(gen[4972]),

			.SO(gen[5065]),
			.S(gen[5066]),
			.SE(gen[5067]),

			.SELF(gen[4971]),
			.cell_state(gen[4971])
		); 

/******************* CELL 4972 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4972 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4876]),
			.N(gen[4877]),
			.NE(gen[4878]),

			.O(gen[4971]),
			.E(gen[4973]),

			.SO(gen[5066]),
			.S(gen[5067]),
			.SE(gen[5068]),

			.SELF(gen[4972]),
			.cell_state(gen[4972])
		); 

/******************* CELL 4973 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4973 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4877]),
			.N(gen[4878]),
			.NE(gen[4879]),

			.O(gen[4972]),
			.E(gen[4974]),

			.SO(gen[5067]),
			.S(gen[5068]),
			.SE(gen[5069]),

			.SELF(gen[4973]),
			.cell_state(gen[4973])
		); 

/******************* CELL 4974 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4974 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4878]),
			.N(gen[4879]),
			.NE(gen[4880]),

			.O(gen[4973]),
			.E(gen[4975]),

			.SO(gen[5068]),
			.S(gen[5069]),
			.SE(gen[5070]),

			.SELF(gen[4974]),
			.cell_state(gen[4974])
		); 

/******************* CELL 4975 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4975 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4879]),
			.N(gen[4880]),
			.NE(gen[4881]),

			.O(gen[4974]),
			.E(gen[4976]),

			.SO(gen[5069]),
			.S(gen[5070]),
			.SE(gen[5071]),

			.SELF(gen[4975]),
			.cell_state(gen[4975])
		); 

/******************* CELL 4976 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4976 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4880]),
			.N(gen[4881]),
			.NE(gen[4882]),

			.O(gen[4975]),
			.E(gen[4977]),

			.SO(gen[5070]),
			.S(gen[5071]),
			.SE(gen[5072]),

			.SELF(gen[4976]),
			.cell_state(gen[4976])
		); 

/******************* CELL 4977 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4977 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4881]),
			.N(gen[4882]),
			.NE(gen[4883]),

			.O(gen[4976]),
			.E(gen[4978]),

			.SO(gen[5071]),
			.S(gen[5072]),
			.SE(gen[5073]),

			.SELF(gen[4977]),
			.cell_state(gen[4977])
		); 

/******************* CELL 4978 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4978 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4882]),
			.N(gen[4883]),
			.NE(gen[4884]),

			.O(gen[4977]),
			.E(gen[4979]),

			.SO(gen[5072]),
			.S(gen[5073]),
			.SE(gen[5074]),

			.SELF(gen[4978]),
			.cell_state(gen[4978])
		); 

/******************* CELL 4979 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4979 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4883]),
			.N(gen[4884]),
			.NE(gen[4885]),

			.O(gen[4978]),
			.E(gen[4980]),

			.SO(gen[5073]),
			.S(gen[5074]),
			.SE(gen[5075]),

			.SELF(gen[4979]),
			.cell_state(gen[4979])
		); 

/******************* CELL 4980 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4980 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4884]),
			.N(gen[4885]),
			.NE(gen[4886]),

			.O(gen[4979]),
			.E(gen[4981]),

			.SO(gen[5074]),
			.S(gen[5075]),
			.SE(gen[5076]),

			.SELF(gen[4980]),
			.cell_state(gen[4980])
		); 

/******************* CELL 4981 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4981 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4885]),
			.N(gen[4886]),
			.NE(gen[4887]),

			.O(gen[4980]),
			.E(gen[4982]),

			.SO(gen[5075]),
			.S(gen[5076]),
			.SE(gen[5077]),

			.SELF(gen[4981]),
			.cell_state(gen[4981])
		); 

/******************* CELL 4982 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4982 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4886]),
			.N(gen[4887]),
			.NE(gen[4888]),

			.O(gen[4981]),
			.E(gen[4983]),

			.SO(gen[5076]),
			.S(gen[5077]),
			.SE(gen[5078]),

			.SELF(gen[4982]),
			.cell_state(gen[4982])
		); 

/******************* CELL 4983 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4983 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4887]),
			.N(gen[4888]),
			.NE(gen[4889]),

			.O(gen[4982]),
			.E(gen[4984]),

			.SO(gen[5077]),
			.S(gen[5078]),
			.SE(gen[5079]),

			.SELF(gen[4983]),
			.cell_state(gen[4983])
		); 

/******************* CELL 4984 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4984 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4888]),
			.N(gen[4889]),
			.NE(gen[4890]),

			.O(gen[4983]),
			.E(gen[4985]),

			.SO(gen[5078]),
			.S(gen[5079]),
			.SE(gen[5080]),

			.SELF(gen[4984]),
			.cell_state(gen[4984])
		); 

/******************* CELL 4985 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4985 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4889]),
			.N(gen[4890]),
			.NE(gen[4891]),

			.O(gen[4984]),
			.E(gen[4986]),

			.SO(gen[5079]),
			.S(gen[5080]),
			.SE(gen[5081]),

			.SELF(gen[4985]),
			.cell_state(gen[4985])
		); 

/******************* CELL 4986 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4986 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4890]),
			.N(gen[4891]),
			.NE(gen[4892]),

			.O(gen[4985]),
			.E(gen[4987]),

			.SO(gen[5080]),
			.S(gen[5081]),
			.SE(gen[5082]),

			.SELF(gen[4986]),
			.cell_state(gen[4986])
		); 

/******************* CELL 4987 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4987 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4891]),
			.N(gen[4892]),
			.NE(gen[4893]),

			.O(gen[4986]),
			.E(gen[4988]),

			.SO(gen[5081]),
			.S(gen[5082]),
			.SE(gen[5083]),

			.SELF(gen[4987]),
			.cell_state(gen[4987])
		); 

/******************* CELL 4988 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4988 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4892]),
			.N(gen[4893]),
			.NE(gen[4894]),

			.O(gen[4987]),
			.E(gen[4989]),

			.SO(gen[5082]),
			.S(gen[5083]),
			.SE(gen[5084]),

			.SELF(gen[4988]),
			.cell_state(gen[4988])
		); 

/******************* CELL 4989 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4989 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4893]),
			.N(gen[4894]),
			.NE(gen[4895]),

			.O(gen[4988]),
			.E(gen[4990]),

			.SO(gen[5083]),
			.S(gen[5084]),
			.SE(gen[5085]),

			.SELF(gen[4989]),
			.cell_state(gen[4989])
		); 

/******************* CELL 4990 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4990 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4894]),
			.N(gen[4895]),
			.NE(gen[4896]),

			.O(gen[4989]),
			.E(gen[4991]),

			.SO(gen[5084]),
			.S(gen[5085]),
			.SE(gen[5086]),

			.SELF(gen[4990]),
			.cell_state(gen[4990])
		); 

/******************* CELL 4991 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4991 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4895]),
			.N(gen[4896]),
			.NE(gen[4897]),

			.O(gen[4990]),
			.E(gen[4992]),

			.SO(gen[5085]),
			.S(gen[5086]),
			.SE(gen[5087]),

			.SELF(gen[4991]),
			.cell_state(gen[4991])
		); 

/******************* CELL 4992 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4992 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4896]),
			.N(gen[4897]),
			.NE(gen[4898]),

			.O(gen[4991]),
			.E(gen[4993]),

			.SO(gen[5086]),
			.S(gen[5087]),
			.SE(gen[5088]),

			.SELF(gen[4992]),
			.cell_state(gen[4992])
		); 

/******************* CELL 4993 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4993 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4897]),
			.N(gen[4898]),
			.NE(gen[4899]),

			.O(gen[4992]),
			.E(gen[4994]),

			.SO(gen[5087]),
			.S(gen[5088]),
			.SE(gen[5089]),

			.SELF(gen[4993]),
			.cell_state(gen[4993])
		); 

/******************* CELL 4994 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4994 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4898]),
			.N(gen[4899]),
			.NE(gen[4900]),

			.O(gen[4993]),
			.E(gen[4995]),

			.SO(gen[5088]),
			.S(gen[5089]),
			.SE(gen[5090]),

			.SELF(gen[4994]),
			.cell_state(gen[4994])
		); 

/******************* CELL 4995 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4995 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4899]),
			.N(gen[4900]),
			.NE(gen[4901]),

			.O(gen[4994]),
			.E(gen[4996]),

			.SO(gen[5089]),
			.S(gen[5090]),
			.SE(gen[5091]),

			.SELF(gen[4995]),
			.cell_state(gen[4995])
		); 

/******************* CELL 4996 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4996 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4900]),
			.N(gen[4901]),
			.NE(gen[4902]),

			.O(gen[4995]),
			.E(gen[4997]),

			.SO(gen[5090]),
			.S(gen[5091]),
			.SE(gen[5092]),

			.SELF(gen[4996]),
			.cell_state(gen[4996])
		); 

/******************* CELL 4997 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4997 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4901]),
			.N(gen[4902]),
			.NE(gen[4903]),

			.O(gen[4996]),
			.E(gen[4998]),

			.SO(gen[5091]),
			.S(gen[5092]),
			.SE(gen[5093]),

			.SELF(gen[4997]),
			.cell_state(gen[4997])
		); 

/******************* CELL 4998 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4998 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4902]),
			.N(gen[4903]),
			.NE(gen[4904]),

			.O(gen[4997]),
			.E(gen[4999]),

			.SO(gen[5092]),
			.S(gen[5093]),
			.SE(gen[5094]),

			.SELF(gen[4998]),
			.cell_state(gen[4998])
		); 

/******************* CELL 4999 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell4999 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4903]),
			.N(gen[4904]),
			.NE(gen[4905]),

			.O(gen[4998]),
			.E(gen[5000]),

			.SO(gen[5093]),
			.S(gen[5094]),
			.SE(gen[5095]),

			.SELF(gen[4999]),
			.cell_state(gen[4999])
		); 

/******************* CELL 5000 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5000 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4904]),
			.N(gen[4905]),
			.NE(gen[4906]),

			.O(gen[4999]),
			.E(gen[5001]),

			.SO(gen[5094]),
			.S(gen[5095]),
			.SE(gen[5096]),

			.SELF(gen[5000]),
			.cell_state(gen[5000])
		); 

/******************* CELL 5001 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5001 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4905]),
			.N(gen[4906]),
			.NE(gen[4907]),

			.O(gen[5000]),
			.E(gen[5002]),

			.SO(gen[5095]),
			.S(gen[5096]),
			.SE(gen[5097]),

			.SELF(gen[5001]),
			.cell_state(gen[5001])
		); 

/******************* CELL 5002 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5002 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4906]),
			.N(gen[4907]),
			.NE(gen[4908]),

			.O(gen[5001]),
			.E(gen[5003]),

			.SO(gen[5096]),
			.S(gen[5097]),
			.SE(gen[5098]),

			.SELF(gen[5002]),
			.cell_state(gen[5002])
		); 

/******************* CELL 5003 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5003 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4907]),
			.N(gen[4908]),
			.NE(gen[4909]),

			.O(gen[5002]),
			.E(gen[5004]),

			.SO(gen[5097]),
			.S(gen[5098]),
			.SE(gen[5099]),

			.SELF(gen[5003]),
			.cell_state(gen[5003])
		); 

/******************* CELL 5004 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5004 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4908]),
			.N(gen[4909]),
			.NE(gen[4910]),

			.O(gen[5003]),
			.E(gen[5005]),

			.SO(gen[5098]),
			.S(gen[5099]),
			.SE(gen[5100]),

			.SELF(gen[5004]),
			.cell_state(gen[5004])
		); 

/******************* CELL 5005 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5005 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4909]),
			.N(gen[4910]),
			.NE(gen[4911]),

			.O(gen[5004]),
			.E(gen[5006]),

			.SO(gen[5099]),
			.S(gen[5100]),
			.SE(gen[5101]),

			.SELF(gen[5005]),
			.cell_state(gen[5005])
		); 

/******************* CELL 5006 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5006 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4910]),
			.N(gen[4911]),
			.NE(gen[4912]),

			.O(gen[5005]),
			.E(gen[5007]),

			.SO(gen[5100]),
			.S(gen[5101]),
			.SE(gen[5102]),

			.SELF(gen[5006]),
			.cell_state(gen[5006])
		); 

/******************* CELL 5007 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5007 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4911]),
			.N(gen[4912]),
			.NE(gen[4913]),

			.O(gen[5006]),
			.E(gen[5008]),

			.SO(gen[5101]),
			.S(gen[5102]),
			.SE(gen[5103]),

			.SELF(gen[5007]),
			.cell_state(gen[5007])
		); 

/******************* CELL 5008 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5008 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4912]),
			.N(gen[4913]),
			.NE(gen[4914]),

			.O(gen[5007]),
			.E(gen[5009]),

			.SO(gen[5102]),
			.S(gen[5103]),
			.SE(gen[5104]),

			.SELF(gen[5008]),
			.cell_state(gen[5008])
		); 

/******************* CELL 5009 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5009 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4913]),
			.N(gen[4914]),
			.NE(gen[4915]),

			.O(gen[5008]),
			.E(gen[5010]),

			.SO(gen[5103]),
			.S(gen[5104]),
			.SE(gen[5105]),

			.SELF(gen[5009]),
			.cell_state(gen[5009])
		); 

/******************* CELL 5010 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5010 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4914]),
			.N(gen[4915]),
			.NE(gen[4916]),

			.O(gen[5009]),
			.E(gen[5011]),

			.SO(gen[5104]),
			.S(gen[5105]),
			.SE(gen[5106]),

			.SELF(gen[5010]),
			.cell_state(gen[5010])
		); 

/******************* CELL 5011 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5011 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4915]),
			.N(gen[4916]),
			.NE(gen[4917]),

			.O(gen[5010]),
			.E(gen[5012]),

			.SO(gen[5105]),
			.S(gen[5106]),
			.SE(gen[5107]),

			.SELF(gen[5011]),
			.cell_state(gen[5011])
		); 

/******************* CELL 5012 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5012 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4916]),
			.N(gen[4917]),
			.NE(gen[4918]),

			.O(gen[5011]),
			.E(gen[5013]),

			.SO(gen[5106]),
			.S(gen[5107]),
			.SE(gen[5108]),

			.SELF(gen[5012]),
			.cell_state(gen[5012])
		); 

/******************* CELL 5013 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5013 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4917]),
			.N(gen[4918]),
			.NE(gen[4919]),

			.O(gen[5012]),
			.E(gen[5014]),

			.SO(gen[5107]),
			.S(gen[5108]),
			.SE(gen[5109]),

			.SELF(gen[5013]),
			.cell_state(gen[5013])
		); 

/******************* CELL 5014 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5014 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4918]),
			.N(gen[4919]),
			.NE(gen[4920]),

			.O(gen[5013]),
			.E(gen[5015]),

			.SO(gen[5108]),
			.S(gen[5109]),
			.SE(gen[5110]),

			.SELF(gen[5014]),
			.cell_state(gen[5014])
		); 

/******************* CELL 5015 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5015 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4919]),
			.N(gen[4920]),
			.NE(gen[4921]),

			.O(gen[5014]),
			.E(gen[5016]),

			.SO(gen[5109]),
			.S(gen[5110]),
			.SE(gen[5111]),

			.SELF(gen[5015]),
			.cell_state(gen[5015])
		); 

/******************* CELL 5016 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5016 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4920]),
			.N(gen[4921]),
			.NE(gen[4922]),

			.O(gen[5015]),
			.E(gen[5017]),

			.SO(gen[5110]),
			.S(gen[5111]),
			.SE(gen[5112]),

			.SELF(gen[5016]),
			.cell_state(gen[5016])
		); 

/******************* CELL 5017 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5017 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4921]),
			.N(gen[4922]),
			.NE(gen[4923]),

			.O(gen[5016]),
			.E(gen[5018]),

			.SO(gen[5111]),
			.S(gen[5112]),
			.SE(gen[5113]),

			.SELF(gen[5017]),
			.cell_state(gen[5017])
		); 

/******************* CELL 5018 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5018 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4922]),
			.N(gen[4923]),
			.NE(gen[4924]),

			.O(gen[5017]),
			.E(gen[5019]),

			.SO(gen[5112]),
			.S(gen[5113]),
			.SE(gen[5114]),

			.SELF(gen[5018]),
			.cell_state(gen[5018])
		); 

/******************* CELL 5019 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5019 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4923]),
			.N(gen[4924]),
			.NE(gen[4925]),

			.O(gen[5018]),
			.E(gen[5020]),

			.SO(gen[5113]),
			.S(gen[5114]),
			.SE(gen[5115]),

			.SELF(gen[5019]),
			.cell_state(gen[5019])
		); 

/******************* CELL 5020 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5020 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4924]),
			.N(gen[4925]),
			.NE(gen[4926]),

			.O(gen[5019]),
			.E(gen[5021]),

			.SO(gen[5114]),
			.S(gen[5115]),
			.SE(gen[5116]),

			.SELF(gen[5020]),
			.cell_state(gen[5020])
		); 

/******************* CELL 5021 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5021 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4925]),
			.N(gen[4926]),
			.NE(gen[4927]),

			.O(gen[5020]),
			.E(gen[5022]),

			.SO(gen[5115]),
			.S(gen[5116]),
			.SE(gen[5117]),

			.SELF(gen[5021]),
			.cell_state(gen[5021])
		); 

/******************* CELL 5022 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5022 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4926]),
			.N(gen[4927]),
			.NE(gen[4928]),

			.O(gen[5021]),
			.E(gen[5023]),

			.SO(gen[5116]),
			.S(gen[5117]),
			.SE(gen[5118]),

			.SELF(gen[5022]),
			.cell_state(gen[5022])
		); 

/******************* CELL 5023 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5023 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4927]),
			.N(gen[4928]),
			.NE(gen[4929]),

			.O(gen[5022]),
			.E(gen[5024]),

			.SO(gen[5117]),
			.S(gen[5118]),
			.SE(gen[5119]),

			.SELF(gen[5023]),
			.cell_state(gen[5023])
		); 

/******************* CELL 5024 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5024 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4928]),
			.N(gen[4929]),
			.NE(gen[4930]),

			.O(gen[5023]),
			.E(gen[5025]),

			.SO(gen[5118]),
			.S(gen[5119]),
			.SE(gen[5120]),

			.SELF(gen[5024]),
			.cell_state(gen[5024])
		); 

/******************* CELL 5025 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5025 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4929]),
			.N(gen[4930]),
			.NE(gen[4931]),

			.O(gen[5024]),
			.E(gen[5026]),

			.SO(gen[5119]),
			.S(gen[5120]),
			.SE(gen[5121]),

			.SELF(gen[5025]),
			.cell_state(gen[5025])
		); 

/******************* CELL 5026 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5026 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4930]),
			.N(gen[4931]),
			.NE(gen[4932]),

			.O(gen[5025]),
			.E(gen[5027]),

			.SO(gen[5120]),
			.S(gen[5121]),
			.SE(gen[5122]),

			.SELF(gen[5026]),
			.cell_state(gen[5026])
		); 

/******************* CELL 5027 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5027 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4931]),
			.N(gen[4932]),
			.NE(gen[4933]),

			.O(gen[5026]),
			.E(gen[5028]),

			.SO(gen[5121]),
			.S(gen[5122]),
			.SE(gen[5123]),

			.SELF(gen[5027]),
			.cell_state(gen[5027])
		); 

/******************* CELL 5028 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5028 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4932]),
			.N(gen[4933]),
			.NE(gen[4934]),

			.O(gen[5027]),
			.E(gen[5029]),

			.SO(gen[5122]),
			.S(gen[5123]),
			.SE(gen[5124]),

			.SELF(gen[5028]),
			.cell_state(gen[5028])
		); 

/******************* CELL 5029 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5029 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4933]),
			.N(gen[4934]),
			.NE(gen[4935]),

			.O(gen[5028]),
			.E(gen[5030]),

			.SO(gen[5123]),
			.S(gen[5124]),
			.SE(gen[5125]),

			.SELF(gen[5029]),
			.cell_state(gen[5029])
		); 

/******************* CELL 5030 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5030 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4934]),
			.N(gen[4935]),
			.NE(gen[4936]),

			.O(gen[5029]),
			.E(gen[5031]),

			.SO(gen[5124]),
			.S(gen[5125]),
			.SE(gen[5126]),

			.SELF(gen[5030]),
			.cell_state(gen[5030])
		); 

/******************* CELL 5031 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5031 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4935]),
			.N(gen[4936]),
			.NE(gen[4937]),

			.O(gen[5030]),
			.E(gen[5032]),

			.SO(gen[5125]),
			.S(gen[5126]),
			.SE(gen[5127]),

			.SELF(gen[5031]),
			.cell_state(gen[5031])
		); 

/******************* CELL 5032 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5032 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4936]),
			.N(gen[4937]),
			.NE(gen[4938]),

			.O(gen[5031]),
			.E(gen[5033]),

			.SO(gen[5126]),
			.S(gen[5127]),
			.SE(gen[5128]),

			.SELF(gen[5032]),
			.cell_state(gen[5032])
		); 

/******************* CELL 5033 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5033 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4937]),
			.N(gen[4938]),
			.NE(gen[4939]),

			.O(gen[5032]),
			.E(gen[5034]),

			.SO(gen[5127]),
			.S(gen[5128]),
			.SE(gen[5129]),

			.SELF(gen[5033]),
			.cell_state(gen[5033])
		); 

/******************* CELL 5034 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5034 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4938]),
			.N(gen[4939]),
			.NE(gen[4938]),

			.O(gen[5033]),
			.E(gen[5033]),

			.SO(gen[5128]),
			.S(gen[5129]),
			.SE(gen[5128]),

			.SELF(gen[5034]),
			.cell_state(gen[5034])
		); 

/******************* CELL 5035 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5035 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4941]),
			.N(gen[4940]),
			.NE(gen[4941]),

			.O(gen[5036]),
			.E(gen[5036]),

			.SO(gen[5131]),
			.S(gen[5130]),
			.SE(gen[5131]),

			.SELF(gen[5035]),
			.cell_state(gen[5035])
		); 

/******************* CELL 5036 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5036 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4940]),
			.N(gen[4941]),
			.NE(gen[4942]),

			.O(gen[5035]),
			.E(gen[5037]),

			.SO(gen[5130]),
			.S(gen[5131]),
			.SE(gen[5132]),

			.SELF(gen[5036]),
			.cell_state(gen[5036])
		); 

/******************* CELL 5037 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5037 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4941]),
			.N(gen[4942]),
			.NE(gen[4943]),

			.O(gen[5036]),
			.E(gen[5038]),

			.SO(gen[5131]),
			.S(gen[5132]),
			.SE(gen[5133]),

			.SELF(gen[5037]),
			.cell_state(gen[5037])
		); 

/******************* CELL 5038 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5038 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4942]),
			.N(gen[4943]),
			.NE(gen[4944]),

			.O(gen[5037]),
			.E(gen[5039]),

			.SO(gen[5132]),
			.S(gen[5133]),
			.SE(gen[5134]),

			.SELF(gen[5038]),
			.cell_state(gen[5038])
		); 

/******************* CELL 5039 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5039 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4943]),
			.N(gen[4944]),
			.NE(gen[4945]),

			.O(gen[5038]),
			.E(gen[5040]),

			.SO(gen[5133]),
			.S(gen[5134]),
			.SE(gen[5135]),

			.SELF(gen[5039]),
			.cell_state(gen[5039])
		); 

/******************* CELL 5040 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5040 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4944]),
			.N(gen[4945]),
			.NE(gen[4946]),

			.O(gen[5039]),
			.E(gen[5041]),

			.SO(gen[5134]),
			.S(gen[5135]),
			.SE(gen[5136]),

			.SELF(gen[5040]),
			.cell_state(gen[5040])
		); 

/******************* CELL 5041 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5041 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4945]),
			.N(gen[4946]),
			.NE(gen[4947]),

			.O(gen[5040]),
			.E(gen[5042]),

			.SO(gen[5135]),
			.S(gen[5136]),
			.SE(gen[5137]),

			.SELF(gen[5041]),
			.cell_state(gen[5041])
		); 

/******************* CELL 5042 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5042 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4946]),
			.N(gen[4947]),
			.NE(gen[4948]),

			.O(gen[5041]),
			.E(gen[5043]),

			.SO(gen[5136]),
			.S(gen[5137]),
			.SE(gen[5138]),

			.SELF(gen[5042]),
			.cell_state(gen[5042])
		); 

/******************* CELL 5043 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5043 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4947]),
			.N(gen[4948]),
			.NE(gen[4949]),

			.O(gen[5042]),
			.E(gen[5044]),

			.SO(gen[5137]),
			.S(gen[5138]),
			.SE(gen[5139]),

			.SELF(gen[5043]),
			.cell_state(gen[5043])
		); 

/******************* CELL 5044 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5044 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4948]),
			.N(gen[4949]),
			.NE(gen[4950]),

			.O(gen[5043]),
			.E(gen[5045]),

			.SO(gen[5138]),
			.S(gen[5139]),
			.SE(gen[5140]),

			.SELF(gen[5044]),
			.cell_state(gen[5044])
		); 

/******************* CELL 5045 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5045 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4949]),
			.N(gen[4950]),
			.NE(gen[4951]),

			.O(gen[5044]),
			.E(gen[5046]),

			.SO(gen[5139]),
			.S(gen[5140]),
			.SE(gen[5141]),

			.SELF(gen[5045]),
			.cell_state(gen[5045])
		); 

/******************* CELL 5046 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5046 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4950]),
			.N(gen[4951]),
			.NE(gen[4952]),

			.O(gen[5045]),
			.E(gen[5047]),

			.SO(gen[5140]),
			.S(gen[5141]),
			.SE(gen[5142]),

			.SELF(gen[5046]),
			.cell_state(gen[5046])
		); 

/******************* CELL 5047 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5047 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4951]),
			.N(gen[4952]),
			.NE(gen[4953]),

			.O(gen[5046]),
			.E(gen[5048]),

			.SO(gen[5141]),
			.S(gen[5142]),
			.SE(gen[5143]),

			.SELF(gen[5047]),
			.cell_state(gen[5047])
		); 

/******************* CELL 5048 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5048 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4952]),
			.N(gen[4953]),
			.NE(gen[4954]),

			.O(gen[5047]),
			.E(gen[5049]),

			.SO(gen[5142]),
			.S(gen[5143]),
			.SE(gen[5144]),

			.SELF(gen[5048]),
			.cell_state(gen[5048])
		); 

/******************* CELL 5049 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5049 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4953]),
			.N(gen[4954]),
			.NE(gen[4955]),

			.O(gen[5048]),
			.E(gen[5050]),

			.SO(gen[5143]),
			.S(gen[5144]),
			.SE(gen[5145]),

			.SELF(gen[5049]),
			.cell_state(gen[5049])
		); 

/******************* CELL 5050 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5050 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4954]),
			.N(gen[4955]),
			.NE(gen[4956]),

			.O(gen[5049]),
			.E(gen[5051]),

			.SO(gen[5144]),
			.S(gen[5145]),
			.SE(gen[5146]),

			.SELF(gen[5050]),
			.cell_state(gen[5050])
		); 

/******************* CELL 5051 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5051 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4955]),
			.N(gen[4956]),
			.NE(gen[4957]),

			.O(gen[5050]),
			.E(gen[5052]),

			.SO(gen[5145]),
			.S(gen[5146]),
			.SE(gen[5147]),

			.SELF(gen[5051]),
			.cell_state(gen[5051])
		); 

/******************* CELL 5052 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5052 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4956]),
			.N(gen[4957]),
			.NE(gen[4958]),

			.O(gen[5051]),
			.E(gen[5053]),

			.SO(gen[5146]),
			.S(gen[5147]),
			.SE(gen[5148]),

			.SELF(gen[5052]),
			.cell_state(gen[5052])
		); 

/******************* CELL 5053 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5053 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4957]),
			.N(gen[4958]),
			.NE(gen[4959]),

			.O(gen[5052]),
			.E(gen[5054]),

			.SO(gen[5147]),
			.S(gen[5148]),
			.SE(gen[5149]),

			.SELF(gen[5053]),
			.cell_state(gen[5053])
		); 

/******************* CELL 5054 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5054 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4958]),
			.N(gen[4959]),
			.NE(gen[4960]),

			.O(gen[5053]),
			.E(gen[5055]),

			.SO(gen[5148]),
			.S(gen[5149]),
			.SE(gen[5150]),

			.SELF(gen[5054]),
			.cell_state(gen[5054])
		); 

/******************* CELL 5055 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5055 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4959]),
			.N(gen[4960]),
			.NE(gen[4961]),

			.O(gen[5054]),
			.E(gen[5056]),

			.SO(gen[5149]),
			.S(gen[5150]),
			.SE(gen[5151]),

			.SELF(gen[5055]),
			.cell_state(gen[5055])
		); 

/******************* CELL 5056 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5056 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4960]),
			.N(gen[4961]),
			.NE(gen[4962]),

			.O(gen[5055]),
			.E(gen[5057]),

			.SO(gen[5150]),
			.S(gen[5151]),
			.SE(gen[5152]),

			.SELF(gen[5056]),
			.cell_state(gen[5056])
		); 

/******************* CELL 5057 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5057 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4961]),
			.N(gen[4962]),
			.NE(gen[4963]),

			.O(gen[5056]),
			.E(gen[5058]),

			.SO(gen[5151]),
			.S(gen[5152]),
			.SE(gen[5153]),

			.SELF(gen[5057]),
			.cell_state(gen[5057])
		); 

/******************* CELL 5058 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5058 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4962]),
			.N(gen[4963]),
			.NE(gen[4964]),

			.O(gen[5057]),
			.E(gen[5059]),

			.SO(gen[5152]),
			.S(gen[5153]),
			.SE(gen[5154]),

			.SELF(gen[5058]),
			.cell_state(gen[5058])
		); 

/******************* CELL 5059 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5059 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4963]),
			.N(gen[4964]),
			.NE(gen[4965]),

			.O(gen[5058]),
			.E(gen[5060]),

			.SO(gen[5153]),
			.S(gen[5154]),
			.SE(gen[5155]),

			.SELF(gen[5059]),
			.cell_state(gen[5059])
		); 

/******************* CELL 5060 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5060 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4964]),
			.N(gen[4965]),
			.NE(gen[4966]),

			.O(gen[5059]),
			.E(gen[5061]),

			.SO(gen[5154]),
			.S(gen[5155]),
			.SE(gen[5156]),

			.SELF(gen[5060]),
			.cell_state(gen[5060])
		); 

/******************* CELL 5061 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5061 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4965]),
			.N(gen[4966]),
			.NE(gen[4967]),

			.O(gen[5060]),
			.E(gen[5062]),

			.SO(gen[5155]),
			.S(gen[5156]),
			.SE(gen[5157]),

			.SELF(gen[5061]),
			.cell_state(gen[5061])
		); 

/******************* CELL 5062 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5062 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4966]),
			.N(gen[4967]),
			.NE(gen[4968]),

			.O(gen[5061]),
			.E(gen[5063]),

			.SO(gen[5156]),
			.S(gen[5157]),
			.SE(gen[5158]),

			.SELF(gen[5062]),
			.cell_state(gen[5062])
		); 

/******************* CELL 5063 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5063 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4967]),
			.N(gen[4968]),
			.NE(gen[4969]),

			.O(gen[5062]),
			.E(gen[5064]),

			.SO(gen[5157]),
			.S(gen[5158]),
			.SE(gen[5159]),

			.SELF(gen[5063]),
			.cell_state(gen[5063])
		); 

/******************* CELL 5064 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5064 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4968]),
			.N(gen[4969]),
			.NE(gen[4970]),

			.O(gen[5063]),
			.E(gen[5065]),

			.SO(gen[5158]),
			.S(gen[5159]),
			.SE(gen[5160]),

			.SELF(gen[5064]),
			.cell_state(gen[5064])
		); 

/******************* CELL 5065 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5065 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4969]),
			.N(gen[4970]),
			.NE(gen[4971]),

			.O(gen[5064]),
			.E(gen[5066]),

			.SO(gen[5159]),
			.S(gen[5160]),
			.SE(gen[5161]),

			.SELF(gen[5065]),
			.cell_state(gen[5065])
		); 

/******************* CELL 5066 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5066 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4970]),
			.N(gen[4971]),
			.NE(gen[4972]),

			.O(gen[5065]),
			.E(gen[5067]),

			.SO(gen[5160]),
			.S(gen[5161]),
			.SE(gen[5162]),

			.SELF(gen[5066]),
			.cell_state(gen[5066])
		); 

/******************* CELL 5067 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5067 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4971]),
			.N(gen[4972]),
			.NE(gen[4973]),

			.O(gen[5066]),
			.E(gen[5068]),

			.SO(gen[5161]),
			.S(gen[5162]),
			.SE(gen[5163]),

			.SELF(gen[5067]),
			.cell_state(gen[5067])
		); 

/******************* CELL 5068 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5068 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4972]),
			.N(gen[4973]),
			.NE(gen[4974]),

			.O(gen[5067]),
			.E(gen[5069]),

			.SO(gen[5162]),
			.S(gen[5163]),
			.SE(gen[5164]),

			.SELF(gen[5068]),
			.cell_state(gen[5068])
		); 

/******************* CELL 5069 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5069 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4973]),
			.N(gen[4974]),
			.NE(gen[4975]),

			.O(gen[5068]),
			.E(gen[5070]),

			.SO(gen[5163]),
			.S(gen[5164]),
			.SE(gen[5165]),

			.SELF(gen[5069]),
			.cell_state(gen[5069])
		); 

/******************* CELL 5070 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5070 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4974]),
			.N(gen[4975]),
			.NE(gen[4976]),

			.O(gen[5069]),
			.E(gen[5071]),

			.SO(gen[5164]),
			.S(gen[5165]),
			.SE(gen[5166]),

			.SELF(gen[5070]),
			.cell_state(gen[5070])
		); 

/******************* CELL 5071 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5071 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4975]),
			.N(gen[4976]),
			.NE(gen[4977]),

			.O(gen[5070]),
			.E(gen[5072]),

			.SO(gen[5165]),
			.S(gen[5166]),
			.SE(gen[5167]),

			.SELF(gen[5071]),
			.cell_state(gen[5071])
		); 

/******************* CELL 5072 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5072 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4976]),
			.N(gen[4977]),
			.NE(gen[4978]),

			.O(gen[5071]),
			.E(gen[5073]),

			.SO(gen[5166]),
			.S(gen[5167]),
			.SE(gen[5168]),

			.SELF(gen[5072]),
			.cell_state(gen[5072])
		); 

/******************* CELL 5073 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5073 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4977]),
			.N(gen[4978]),
			.NE(gen[4979]),

			.O(gen[5072]),
			.E(gen[5074]),

			.SO(gen[5167]),
			.S(gen[5168]),
			.SE(gen[5169]),

			.SELF(gen[5073]),
			.cell_state(gen[5073])
		); 

/******************* CELL 5074 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5074 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4978]),
			.N(gen[4979]),
			.NE(gen[4980]),

			.O(gen[5073]),
			.E(gen[5075]),

			.SO(gen[5168]),
			.S(gen[5169]),
			.SE(gen[5170]),

			.SELF(gen[5074]),
			.cell_state(gen[5074])
		); 

/******************* CELL 5075 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5075 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4979]),
			.N(gen[4980]),
			.NE(gen[4981]),

			.O(gen[5074]),
			.E(gen[5076]),

			.SO(gen[5169]),
			.S(gen[5170]),
			.SE(gen[5171]),

			.SELF(gen[5075]),
			.cell_state(gen[5075])
		); 

/******************* CELL 5076 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5076 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4980]),
			.N(gen[4981]),
			.NE(gen[4982]),

			.O(gen[5075]),
			.E(gen[5077]),

			.SO(gen[5170]),
			.S(gen[5171]),
			.SE(gen[5172]),

			.SELF(gen[5076]),
			.cell_state(gen[5076])
		); 

/******************* CELL 5077 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5077 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4981]),
			.N(gen[4982]),
			.NE(gen[4983]),

			.O(gen[5076]),
			.E(gen[5078]),

			.SO(gen[5171]),
			.S(gen[5172]),
			.SE(gen[5173]),

			.SELF(gen[5077]),
			.cell_state(gen[5077])
		); 

/******************* CELL 5078 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5078 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4982]),
			.N(gen[4983]),
			.NE(gen[4984]),

			.O(gen[5077]),
			.E(gen[5079]),

			.SO(gen[5172]),
			.S(gen[5173]),
			.SE(gen[5174]),

			.SELF(gen[5078]),
			.cell_state(gen[5078])
		); 

/******************* CELL 5079 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5079 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4983]),
			.N(gen[4984]),
			.NE(gen[4985]),

			.O(gen[5078]),
			.E(gen[5080]),

			.SO(gen[5173]),
			.S(gen[5174]),
			.SE(gen[5175]),

			.SELF(gen[5079]),
			.cell_state(gen[5079])
		); 

/******************* CELL 5080 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5080 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4984]),
			.N(gen[4985]),
			.NE(gen[4986]),

			.O(gen[5079]),
			.E(gen[5081]),

			.SO(gen[5174]),
			.S(gen[5175]),
			.SE(gen[5176]),

			.SELF(gen[5080]),
			.cell_state(gen[5080])
		); 

/******************* CELL 5081 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5081 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4985]),
			.N(gen[4986]),
			.NE(gen[4987]),

			.O(gen[5080]),
			.E(gen[5082]),

			.SO(gen[5175]),
			.S(gen[5176]),
			.SE(gen[5177]),

			.SELF(gen[5081]),
			.cell_state(gen[5081])
		); 

/******************* CELL 5082 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5082 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4986]),
			.N(gen[4987]),
			.NE(gen[4988]),

			.O(gen[5081]),
			.E(gen[5083]),

			.SO(gen[5176]),
			.S(gen[5177]),
			.SE(gen[5178]),

			.SELF(gen[5082]),
			.cell_state(gen[5082])
		); 

/******************* CELL 5083 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5083 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4987]),
			.N(gen[4988]),
			.NE(gen[4989]),

			.O(gen[5082]),
			.E(gen[5084]),

			.SO(gen[5177]),
			.S(gen[5178]),
			.SE(gen[5179]),

			.SELF(gen[5083]),
			.cell_state(gen[5083])
		); 

/******************* CELL 5084 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5084 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4988]),
			.N(gen[4989]),
			.NE(gen[4990]),

			.O(gen[5083]),
			.E(gen[5085]),

			.SO(gen[5178]),
			.S(gen[5179]),
			.SE(gen[5180]),

			.SELF(gen[5084]),
			.cell_state(gen[5084])
		); 

/******************* CELL 5085 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5085 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4989]),
			.N(gen[4990]),
			.NE(gen[4991]),

			.O(gen[5084]),
			.E(gen[5086]),

			.SO(gen[5179]),
			.S(gen[5180]),
			.SE(gen[5181]),

			.SELF(gen[5085]),
			.cell_state(gen[5085])
		); 

/******************* CELL 5086 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5086 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4990]),
			.N(gen[4991]),
			.NE(gen[4992]),

			.O(gen[5085]),
			.E(gen[5087]),

			.SO(gen[5180]),
			.S(gen[5181]),
			.SE(gen[5182]),

			.SELF(gen[5086]),
			.cell_state(gen[5086])
		); 

/******************* CELL 5087 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5087 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4991]),
			.N(gen[4992]),
			.NE(gen[4993]),

			.O(gen[5086]),
			.E(gen[5088]),

			.SO(gen[5181]),
			.S(gen[5182]),
			.SE(gen[5183]),

			.SELF(gen[5087]),
			.cell_state(gen[5087])
		); 

/******************* CELL 5088 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5088 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4992]),
			.N(gen[4993]),
			.NE(gen[4994]),

			.O(gen[5087]),
			.E(gen[5089]),

			.SO(gen[5182]),
			.S(gen[5183]),
			.SE(gen[5184]),

			.SELF(gen[5088]),
			.cell_state(gen[5088])
		); 

/******************* CELL 5089 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5089 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4993]),
			.N(gen[4994]),
			.NE(gen[4995]),

			.O(gen[5088]),
			.E(gen[5090]),

			.SO(gen[5183]),
			.S(gen[5184]),
			.SE(gen[5185]),

			.SELF(gen[5089]),
			.cell_state(gen[5089])
		); 

/******************* CELL 5090 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5090 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4994]),
			.N(gen[4995]),
			.NE(gen[4996]),

			.O(gen[5089]),
			.E(gen[5091]),

			.SO(gen[5184]),
			.S(gen[5185]),
			.SE(gen[5186]),

			.SELF(gen[5090]),
			.cell_state(gen[5090])
		); 

/******************* CELL 5091 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5091 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4995]),
			.N(gen[4996]),
			.NE(gen[4997]),

			.O(gen[5090]),
			.E(gen[5092]),

			.SO(gen[5185]),
			.S(gen[5186]),
			.SE(gen[5187]),

			.SELF(gen[5091]),
			.cell_state(gen[5091])
		); 

/******************* CELL 5092 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5092 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4996]),
			.N(gen[4997]),
			.NE(gen[4998]),

			.O(gen[5091]),
			.E(gen[5093]),

			.SO(gen[5186]),
			.S(gen[5187]),
			.SE(gen[5188]),

			.SELF(gen[5092]),
			.cell_state(gen[5092])
		); 

/******************* CELL 5093 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5093 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4997]),
			.N(gen[4998]),
			.NE(gen[4999]),

			.O(gen[5092]),
			.E(gen[5094]),

			.SO(gen[5187]),
			.S(gen[5188]),
			.SE(gen[5189]),

			.SELF(gen[5093]),
			.cell_state(gen[5093])
		); 

/******************* CELL 5094 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5094 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4998]),
			.N(gen[4999]),
			.NE(gen[5000]),

			.O(gen[5093]),
			.E(gen[5095]),

			.SO(gen[5188]),
			.S(gen[5189]),
			.SE(gen[5190]),

			.SELF(gen[5094]),
			.cell_state(gen[5094])
		); 

/******************* CELL 5095 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5095 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4999]),
			.N(gen[5000]),
			.NE(gen[5001]),

			.O(gen[5094]),
			.E(gen[5096]),

			.SO(gen[5189]),
			.S(gen[5190]),
			.SE(gen[5191]),

			.SELF(gen[5095]),
			.cell_state(gen[5095])
		); 

/******************* CELL 5096 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5096 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5000]),
			.N(gen[5001]),
			.NE(gen[5002]),

			.O(gen[5095]),
			.E(gen[5097]),

			.SO(gen[5190]),
			.S(gen[5191]),
			.SE(gen[5192]),

			.SELF(gen[5096]),
			.cell_state(gen[5096])
		); 

/******************* CELL 5097 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5097 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5001]),
			.N(gen[5002]),
			.NE(gen[5003]),

			.O(gen[5096]),
			.E(gen[5098]),

			.SO(gen[5191]),
			.S(gen[5192]),
			.SE(gen[5193]),

			.SELF(gen[5097]),
			.cell_state(gen[5097])
		); 

/******************* CELL 5098 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5098 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5002]),
			.N(gen[5003]),
			.NE(gen[5004]),

			.O(gen[5097]),
			.E(gen[5099]),

			.SO(gen[5192]),
			.S(gen[5193]),
			.SE(gen[5194]),

			.SELF(gen[5098]),
			.cell_state(gen[5098])
		); 

/******************* CELL 5099 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5099 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5003]),
			.N(gen[5004]),
			.NE(gen[5005]),

			.O(gen[5098]),
			.E(gen[5100]),

			.SO(gen[5193]),
			.S(gen[5194]),
			.SE(gen[5195]),

			.SELF(gen[5099]),
			.cell_state(gen[5099])
		); 

/******************* CELL 5100 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5100 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5004]),
			.N(gen[5005]),
			.NE(gen[5006]),

			.O(gen[5099]),
			.E(gen[5101]),

			.SO(gen[5194]),
			.S(gen[5195]),
			.SE(gen[5196]),

			.SELF(gen[5100]),
			.cell_state(gen[5100])
		); 

/******************* CELL 5101 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5101 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5005]),
			.N(gen[5006]),
			.NE(gen[5007]),

			.O(gen[5100]),
			.E(gen[5102]),

			.SO(gen[5195]),
			.S(gen[5196]),
			.SE(gen[5197]),

			.SELF(gen[5101]),
			.cell_state(gen[5101])
		); 

/******************* CELL 5102 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5102 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5006]),
			.N(gen[5007]),
			.NE(gen[5008]),

			.O(gen[5101]),
			.E(gen[5103]),

			.SO(gen[5196]),
			.S(gen[5197]),
			.SE(gen[5198]),

			.SELF(gen[5102]),
			.cell_state(gen[5102])
		); 

/******************* CELL 5103 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5103 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5007]),
			.N(gen[5008]),
			.NE(gen[5009]),

			.O(gen[5102]),
			.E(gen[5104]),

			.SO(gen[5197]),
			.S(gen[5198]),
			.SE(gen[5199]),

			.SELF(gen[5103]),
			.cell_state(gen[5103])
		); 

/******************* CELL 5104 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5104 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5008]),
			.N(gen[5009]),
			.NE(gen[5010]),

			.O(gen[5103]),
			.E(gen[5105]),

			.SO(gen[5198]),
			.S(gen[5199]),
			.SE(gen[5200]),

			.SELF(gen[5104]),
			.cell_state(gen[5104])
		); 

/******************* CELL 5105 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5105 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5009]),
			.N(gen[5010]),
			.NE(gen[5011]),

			.O(gen[5104]),
			.E(gen[5106]),

			.SO(gen[5199]),
			.S(gen[5200]),
			.SE(gen[5201]),

			.SELF(gen[5105]),
			.cell_state(gen[5105])
		); 

/******************* CELL 5106 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5106 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5010]),
			.N(gen[5011]),
			.NE(gen[5012]),

			.O(gen[5105]),
			.E(gen[5107]),

			.SO(gen[5200]),
			.S(gen[5201]),
			.SE(gen[5202]),

			.SELF(gen[5106]),
			.cell_state(gen[5106])
		); 

/******************* CELL 5107 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5107 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5011]),
			.N(gen[5012]),
			.NE(gen[5013]),

			.O(gen[5106]),
			.E(gen[5108]),

			.SO(gen[5201]),
			.S(gen[5202]),
			.SE(gen[5203]),

			.SELF(gen[5107]),
			.cell_state(gen[5107])
		); 

/******************* CELL 5108 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5108 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5012]),
			.N(gen[5013]),
			.NE(gen[5014]),

			.O(gen[5107]),
			.E(gen[5109]),

			.SO(gen[5202]),
			.S(gen[5203]),
			.SE(gen[5204]),

			.SELF(gen[5108]),
			.cell_state(gen[5108])
		); 

/******************* CELL 5109 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5109 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5013]),
			.N(gen[5014]),
			.NE(gen[5015]),

			.O(gen[5108]),
			.E(gen[5110]),

			.SO(gen[5203]),
			.S(gen[5204]),
			.SE(gen[5205]),

			.SELF(gen[5109]),
			.cell_state(gen[5109])
		); 

/******************* CELL 5110 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5110 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5014]),
			.N(gen[5015]),
			.NE(gen[5016]),

			.O(gen[5109]),
			.E(gen[5111]),

			.SO(gen[5204]),
			.S(gen[5205]),
			.SE(gen[5206]),

			.SELF(gen[5110]),
			.cell_state(gen[5110])
		); 

/******************* CELL 5111 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5111 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5015]),
			.N(gen[5016]),
			.NE(gen[5017]),

			.O(gen[5110]),
			.E(gen[5112]),

			.SO(gen[5205]),
			.S(gen[5206]),
			.SE(gen[5207]),

			.SELF(gen[5111]),
			.cell_state(gen[5111])
		); 

/******************* CELL 5112 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5112 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5016]),
			.N(gen[5017]),
			.NE(gen[5018]),

			.O(gen[5111]),
			.E(gen[5113]),

			.SO(gen[5206]),
			.S(gen[5207]),
			.SE(gen[5208]),

			.SELF(gen[5112]),
			.cell_state(gen[5112])
		); 

/******************* CELL 5113 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5113 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5017]),
			.N(gen[5018]),
			.NE(gen[5019]),

			.O(gen[5112]),
			.E(gen[5114]),

			.SO(gen[5207]),
			.S(gen[5208]),
			.SE(gen[5209]),

			.SELF(gen[5113]),
			.cell_state(gen[5113])
		); 

/******************* CELL 5114 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5114 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5018]),
			.N(gen[5019]),
			.NE(gen[5020]),

			.O(gen[5113]),
			.E(gen[5115]),

			.SO(gen[5208]),
			.S(gen[5209]),
			.SE(gen[5210]),

			.SELF(gen[5114]),
			.cell_state(gen[5114])
		); 

/******************* CELL 5115 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5115 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5019]),
			.N(gen[5020]),
			.NE(gen[5021]),

			.O(gen[5114]),
			.E(gen[5116]),

			.SO(gen[5209]),
			.S(gen[5210]),
			.SE(gen[5211]),

			.SELF(gen[5115]),
			.cell_state(gen[5115])
		); 

/******************* CELL 5116 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5116 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5020]),
			.N(gen[5021]),
			.NE(gen[5022]),

			.O(gen[5115]),
			.E(gen[5117]),

			.SO(gen[5210]),
			.S(gen[5211]),
			.SE(gen[5212]),

			.SELF(gen[5116]),
			.cell_state(gen[5116])
		); 

/******************* CELL 5117 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5117 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5021]),
			.N(gen[5022]),
			.NE(gen[5023]),

			.O(gen[5116]),
			.E(gen[5118]),

			.SO(gen[5211]),
			.S(gen[5212]),
			.SE(gen[5213]),

			.SELF(gen[5117]),
			.cell_state(gen[5117])
		); 

/******************* CELL 5118 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5118 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5022]),
			.N(gen[5023]),
			.NE(gen[5024]),

			.O(gen[5117]),
			.E(gen[5119]),

			.SO(gen[5212]),
			.S(gen[5213]),
			.SE(gen[5214]),

			.SELF(gen[5118]),
			.cell_state(gen[5118])
		); 

/******************* CELL 5119 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5119 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5023]),
			.N(gen[5024]),
			.NE(gen[5025]),

			.O(gen[5118]),
			.E(gen[5120]),

			.SO(gen[5213]),
			.S(gen[5214]),
			.SE(gen[5215]),

			.SELF(gen[5119]),
			.cell_state(gen[5119])
		); 

/******************* CELL 5120 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5120 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5024]),
			.N(gen[5025]),
			.NE(gen[5026]),

			.O(gen[5119]),
			.E(gen[5121]),

			.SO(gen[5214]),
			.S(gen[5215]),
			.SE(gen[5216]),

			.SELF(gen[5120]),
			.cell_state(gen[5120])
		); 

/******************* CELL 5121 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5121 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5025]),
			.N(gen[5026]),
			.NE(gen[5027]),

			.O(gen[5120]),
			.E(gen[5122]),

			.SO(gen[5215]),
			.S(gen[5216]),
			.SE(gen[5217]),

			.SELF(gen[5121]),
			.cell_state(gen[5121])
		); 

/******************* CELL 5122 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5122 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5026]),
			.N(gen[5027]),
			.NE(gen[5028]),

			.O(gen[5121]),
			.E(gen[5123]),

			.SO(gen[5216]),
			.S(gen[5217]),
			.SE(gen[5218]),

			.SELF(gen[5122]),
			.cell_state(gen[5122])
		); 

/******************* CELL 5123 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5123 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5027]),
			.N(gen[5028]),
			.NE(gen[5029]),

			.O(gen[5122]),
			.E(gen[5124]),

			.SO(gen[5217]),
			.S(gen[5218]),
			.SE(gen[5219]),

			.SELF(gen[5123]),
			.cell_state(gen[5123])
		); 

/******************* CELL 5124 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5124 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5028]),
			.N(gen[5029]),
			.NE(gen[5030]),

			.O(gen[5123]),
			.E(gen[5125]),

			.SO(gen[5218]),
			.S(gen[5219]),
			.SE(gen[5220]),

			.SELF(gen[5124]),
			.cell_state(gen[5124])
		); 

/******************* CELL 5125 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5125 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5029]),
			.N(gen[5030]),
			.NE(gen[5031]),

			.O(gen[5124]),
			.E(gen[5126]),

			.SO(gen[5219]),
			.S(gen[5220]),
			.SE(gen[5221]),

			.SELF(gen[5125]),
			.cell_state(gen[5125])
		); 

/******************* CELL 5126 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5126 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5030]),
			.N(gen[5031]),
			.NE(gen[5032]),

			.O(gen[5125]),
			.E(gen[5127]),

			.SO(gen[5220]),
			.S(gen[5221]),
			.SE(gen[5222]),

			.SELF(gen[5126]),
			.cell_state(gen[5126])
		); 

/******************* CELL 5127 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5127 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5031]),
			.N(gen[5032]),
			.NE(gen[5033]),

			.O(gen[5126]),
			.E(gen[5128]),

			.SO(gen[5221]),
			.S(gen[5222]),
			.SE(gen[5223]),

			.SELF(gen[5127]),
			.cell_state(gen[5127])
		); 

/******************* CELL 5128 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5128 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5032]),
			.N(gen[5033]),
			.NE(gen[5034]),

			.O(gen[5127]),
			.E(gen[5129]),

			.SO(gen[5222]),
			.S(gen[5223]),
			.SE(gen[5224]),

			.SELF(gen[5128]),
			.cell_state(gen[5128])
		); 

/******************* CELL 5129 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5129 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5033]),
			.N(gen[5034]),
			.NE(gen[5033]),

			.O(gen[5128]),
			.E(gen[5128]),

			.SO(gen[5223]),
			.S(gen[5224]),
			.SE(gen[5223]),

			.SELF(gen[5129]),
			.cell_state(gen[5129])
		); 

/******************* CELL 5130 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5130 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5036]),
			.N(gen[5035]),
			.NE(gen[5036]),

			.O(gen[5131]),
			.E(gen[5131]),

			.SO(gen[5226]),
			.S(gen[5225]),
			.SE(gen[5226]),

			.SELF(gen[5130]),
			.cell_state(gen[5130])
		); 

/******************* CELL 5131 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5131 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5035]),
			.N(gen[5036]),
			.NE(gen[5037]),

			.O(gen[5130]),
			.E(gen[5132]),

			.SO(gen[5225]),
			.S(gen[5226]),
			.SE(gen[5227]),

			.SELF(gen[5131]),
			.cell_state(gen[5131])
		); 

/******************* CELL 5132 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5132 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5036]),
			.N(gen[5037]),
			.NE(gen[5038]),

			.O(gen[5131]),
			.E(gen[5133]),

			.SO(gen[5226]),
			.S(gen[5227]),
			.SE(gen[5228]),

			.SELF(gen[5132]),
			.cell_state(gen[5132])
		); 

/******************* CELL 5133 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5133 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5037]),
			.N(gen[5038]),
			.NE(gen[5039]),

			.O(gen[5132]),
			.E(gen[5134]),

			.SO(gen[5227]),
			.S(gen[5228]),
			.SE(gen[5229]),

			.SELF(gen[5133]),
			.cell_state(gen[5133])
		); 

/******************* CELL 5134 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5134 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5038]),
			.N(gen[5039]),
			.NE(gen[5040]),

			.O(gen[5133]),
			.E(gen[5135]),

			.SO(gen[5228]),
			.S(gen[5229]),
			.SE(gen[5230]),

			.SELF(gen[5134]),
			.cell_state(gen[5134])
		); 

/******************* CELL 5135 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5135 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5039]),
			.N(gen[5040]),
			.NE(gen[5041]),

			.O(gen[5134]),
			.E(gen[5136]),

			.SO(gen[5229]),
			.S(gen[5230]),
			.SE(gen[5231]),

			.SELF(gen[5135]),
			.cell_state(gen[5135])
		); 

/******************* CELL 5136 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5136 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5040]),
			.N(gen[5041]),
			.NE(gen[5042]),

			.O(gen[5135]),
			.E(gen[5137]),

			.SO(gen[5230]),
			.S(gen[5231]),
			.SE(gen[5232]),

			.SELF(gen[5136]),
			.cell_state(gen[5136])
		); 

/******************* CELL 5137 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5137 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5041]),
			.N(gen[5042]),
			.NE(gen[5043]),

			.O(gen[5136]),
			.E(gen[5138]),

			.SO(gen[5231]),
			.S(gen[5232]),
			.SE(gen[5233]),

			.SELF(gen[5137]),
			.cell_state(gen[5137])
		); 

/******************* CELL 5138 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5138 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5042]),
			.N(gen[5043]),
			.NE(gen[5044]),

			.O(gen[5137]),
			.E(gen[5139]),

			.SO(gen[5232]),
			.S(gen[5233]),
			.SE(gen[5234]),

			.SELF(gen[5138]),
			.cell_state(gen[5138])
		); 

/******************* CELL 5139 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5139 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5043]),
			.N(gen[5044]),
			.NE(gen[5045]),

			.O(gen[5138]),
			.E(gen[5140]),

			.SO(gen[5233]),
			.S(gen[5234]),
			.SE(gen[5235]),

			.SELF(gen[5139]),
			.cell_state(gen[5139])
		); 

/******************* CELL 5140 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5140 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5044]),
			.N(gen[5045]),
			.NE(gen[5046]),

			.O(gen[5139]),
			.E(gen[5141]),

			.SO(gen[5234]),
			.S(gen[5235]),
			.SE(gen[5236]),

			.SELF(gen[5140]),
			.cell_state(gen[5140])
		); 

/******************* CELL 5141 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5141 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5045]),
			.N(gen[5046]),
			.NE(gen[5047]),

			.O(gen[5140]),
			.E(gen[5142]),

			.SO(gen[5235]),
			.S(gen[5236]),
			.SE(gen[5237]),

			.SELF(gen[5141]),
			.cell_state(gen[5141])
		); 

/******************* CELL 5142 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5142 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5046]),
			.N(gen[5047]),
			.NE(gen[5048]),

			.O(gen[5141]),
			.E(gen[5143]),

			.SO(gen[5236]),
			.S(gen[5237]),
			.SE(gen[5238]),

			.SELF(gen[5142]),
			.cell_state(gen[5142])
		); 

/******************* CELL 5143 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5143 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5047]),
			.N(gen[5048]),
			.NE(gen[5049]),

			.O(gen[5142]),
			.E(gen[5144]),

			.SO(gen[5237]),
			.S(gen[5238]),
			.SE(gen[5239]),

			.SELF(gen[5143]),
			.cell_state(gen[5143])
		); 

/******************* CELL 5144 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5144 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5048]),
			.N(gen[5049]),
			.NE(gen[5050]),

			.O(gen[5143]),
			.E(gen[5145]),

			.SO(gen[5238]),
			.S(gen[5239]),
			.SE(gen[5240]),

			.SELF(gen[5144]),
			.cell_state(gen[5144])
		); 

/******************* CELL 5145 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5145 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5049]),
			.N(gen[5050]),
			.NE(gen[5051]),

			.O(gen[5144]),
			.E(gen[5146]),

			.SO(gen[5239]),
			.S(gen[5240]),
			.SE(gen[5241]),

			.SELF(gen[5145]),
			.cell_state(gen[5145])
		); 

/******************* CELL 5146 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5146 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5050]),
			.N(gen[5051]),
			.NE(gen[5052]),

			.O(gen[5145]),
			.E(gen[5147]),

			.SO(gen[5240]),
			.S(gen[5241]),
			.SE(gen[5242]),

			.SELF(gen[5146]),
			.cell_state(gen[5146])
		); 

/******************* CELL 5147 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5147 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5051]),
			.N(gen[5052]),
			.NE(gen[5053]),

			.O(gen[5146]),
			.E(gen[5148]),

			.SO(gen[5241]),
			.S(gen[5242]),
			.SE(gen[5243]),

			.SELF(gen[5147]),
			.cell_state(gen[5147])
		); 

/******************* CELL 5148 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5148 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5052]),
			.N(gen[5053]),
			.NE(gen[5054]),

			.O(gen[5147]),
			.E(gen[5149]),

			.SO(gen[5242]),
			.S(gen[5243]),
			.SE(gen[5244]),

			.SELF(gen[5148]),
			.cell_state(gen[5148])
		); 

/******************* CELL 5149 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5149 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5053]),
			.N(gen[5054]),
			.NE(gen[5055]),

			.O(gen[5148]),
			.E(gen[5150]),

			.SO(gen[5243]),
			.S(gen[5244]),
			.SE(gen[5245]),

			.SELF(gen[5149]),
			.cell_state(gen[5149])
		); 

/******************* CELL 5150 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5150 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5054]),
			.N(gen[5055]),
			.NE(gen[5056]),

			.O(gen[5149]),
			.E(gen[5151]),

			.SO(gen[5244]),
			.S(gen[5245]),
			.SE(gen[5246]),

			.SELF(gen[5150]),
			.cell_state(gen[5150])
		); 

/******************* CELL 5151 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5151 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5055]),
			.N(gen[5056]),
			.NE(gen[5057]),

			.O(gen[5150]),
			.E(gen[5152]),

			.SO(gen[5245]),
			.S(gen[5246]),
			.SE(gen[5247]),

			.SELF(gen[5151]),
			.cell_state(gen[5151])
		); 

/******************* CELL 5152 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5152 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5056]),
			.N(gen[5057]),
			.NE(gen[5058]),

			.O(gen[5151]),
			.E(gen[5153]),

			.SO(gen[5246]),
			.S(gen[5247]),
			.SE(gen[5248]),

			.SELF(gen[5152]),
			.cell_state(gen[5152])
		); 

/******************* CELL 5153 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5153 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5057]),
			.N(gen[5058]),
			.NE(gen[5059]),

			.O(gen[5152]),
			.E(gen[5154]),

			.SO(gen[5247]),
			.S(gen[5248]),
			.SE(gen[5249]),

			.SELF(gen[5153]),
			.cell_state(gen[5153])
		); 

/******************* CELL 5154 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5154 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5058]),
			.N(gen[5059]),
			.NE(gen[5060]),

			.O(gen[5153]),
			.E(gen[5155]),

			.SO(gen[5248]),
			.S(gen[5249]),
			.SE(gen[5250]),

			.SELF(gen[5154]),
			.cell_state(gen[5154])
		); 

/******************* CELL 5155 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5155 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5059]),
			.N(gen[5060]),
			.NE(gen[5061]),

			.O(gen[5154]),
			.E(gen[5156]),

			.SO(gen[5249]),
			.S(gen[5250]),
			.SE(gen[5251]),

			.SELF(gen[5155]),
			.cell_state(gen[5155])
		); 

/******************* CELL 5156 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5156 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5060]),
			.N(gen[5061]),
			.NE(gen[5062]),

			.O(gen[5155]),
			.E(gen[5157]),

			.SO(gen[5250]),
			.S(gen[5251]),
			.SE(gen[5252]),

			.SELF(gen[5156]),
			.cell_state(gen[5156])
		); 

/******************* CELL 5157 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5157 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5061]),
			.N(gen[5062]),
			.NE(gen[5063]),

			.O(gen[5156]),
			.E(gen[5158]),

			.SO(gen[5251]),
			.S(gen[5252]),
			.SE(gen[5253]),

			.SELF(gen[5157]),
			.cell_state(gen[5157])
		); 

/******************* CELL 5158 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5158 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5062]),
			.N(gen[5063]),
			.NE(gen[5064]),

			.O(gen[5157]),
			.E(gen[5159]),

			.SO(gen[5252]),
			.S(gen[5253]),
			.SE(gen[5254]),

			.SELF(gen[5158]),
			.cell_state(gen[5158])
		); 

/******************* CELL 5159 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5159 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5063]),
			.N(gen[5064]),
			.NE(gen[5065]),

			.O(gen[5158]),
			.E(gen[5160]),

			.SO(gen[5253]),
			.S(gen[5254]),
			.SE(gen[5255]),

			.SELF(gen[5159]),
			.cell_state(gen[5159])
		); 

/******************* CELL 5160 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5160 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5064]),
			.N(gen[5065]),
			.NE(gen[5066]),

			.O(gen[5159]),
			.E(gen[5161]),

			.SO(gen[5254]),
			.S(gen[5255]),
			.SE(gen[5256]),

			.SELF(gen[5160]),
			.cell_state(gen[5160])
		); 

/******************* CELL 5161 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5161 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5065]),
			.N(gen[5066]),
			.NE(gen[5067]),

			.O(gen[5160]),
			.E(gen[5162]),

			.SO(gen[5255]),
			.S(gen[5256]),
			.SE(gen[5257]),

			.SELF(gen[5161]),
			.cell_state(gen[5161])
		); 

/******************* CELL 5162 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5162 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5066]),
			.N(gen[5067]),
			.NE(gen[5068]),

			.O(gen[5161]),
			.E(gen[5163]),

			.SO(gen[5256]),
			.S(gen[5257]),
			.SE(gen[5258]),

			.SELF(gen[5162]),
			.cell_state(gen[5162])
		); 

/******************* CELL 5163 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5163 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5067]),
			.N(gen[5068]),
			.NE(gen[5069]),

			.O(gen[5162]),
			.E(gen[5164]),

			.SO(gen[5257]),
			.S(gen[5258]),
			.SE(gen[5259]),

			.SELF(gen[5163]),
			.cell_state(gen[5163])
		); 

/******************* CELL 5164 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5164 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5068]),
			.N(gen[5069]),
			.NE(gen[5070]),

			.O(gen[5163]),
			.E(gen[5165]),

			.SO(gen[5258]),
			.S(gen[5259]),
			.SE(gen[5260]),

			.SELF(gen[5164]),
			.cell_state(gen[5164])
		); 

/******************* CELL 5165 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5165 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5069]),
			.N(gen[5070]),
			.NE(gen[5071]),

			.O(gen[5164]),
			.E(gen[5166]),

			.SO(gen[5259]),
			.S(gen[5260]),
			.SE(gen[5261]),

			.SELF(gen[5165]),
			.cell_state(gen[5165])
		); 

/******************* CELL 5166 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5166 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5070]),
			.N(gen[5071]),
			.NE(gen[5072]),

			.O(gen[5165]),
			.E(gen[5167]),

			.SO(gen[5260]),
			.S(gen[5261]),
			.SE(gen[5262]),

			.SELF(gen[5166]),
			.cell_state(gen[5166])
		); 

/******************* CELL 5167 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5167 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5071]),
			.N(gen[5072]),
			.NE(gen[5073]),

			.O(gen[5166]),
			.E(gen[5168]),

			.SO(gen[5261]),
			.S(gen[5262]),
			.SE(gen[5263]),

			.SELF(gen[5167]),
			.cell_state(gen[5167])
		); 

/******************* CELL 5168 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5168 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5072]),
			.N(gen[5073]),
			.NE(gen[5074]),

			.O(gen[5167]),
			.E(gen[5169]),

			.SO(gen[5262]),
			.S(gen[5263]),
			.SE(gen[5264]),

			.SELF(gen[5168]),
			.cell_state(gen[5168])
		); 

/******************* CELL 5169 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5169 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5073]),
			.N(gen[5074]),
			.NE(gen[5075]),

			.O(gen[5168]),
			.E(gen[5170]),

			.SO(gen[5263]),
			.S(gen[5264]),
			.SE(gen[5265]),

			.SELF(gen[5169]),
			.cell_state(gen[5169])
		); 

/******************* CELL 5170 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5170 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5074]),
			.N(gen[5075]),
			.NE(gen[5076]),

			.O(gen[5169]),
			.E(gen[5171]),

			.SO(gen[5264]),
			.S(gen[5265]),
			.SE(gen[5266]),

			.SELF(gen[5170]),
			.cell_state(gen[5170])
		); 

/******************* CELL 5171 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5171 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5075]),
			.N(gen[5076]),
			.NE(gen[5077]),

			.O(gen[5170]),
			.E(gen[5172]),

			.SO(gen[5265]),
			.S(gen[5266]),
			.SE(gen[5267]),

			.SELF(gen[5171]),
			.cell_state(gen[5171])
		); 

/******************* CELL 5172 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5172 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5076]),
			.N(gen[5077]),
			.NE(gen[5078]),

			.O(gen[5171]),
			.E(gen[5173]),

			.SO(gen[5266]),
			.S(gen[5267]),
			.SE(gen[5268]),

			.SELF(gen[5172]),
			.cell_state(gen[5172])
		); 

/******************* CELL 5173 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5173 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5077]),
			.N(gen[5078]),
			.NE(gen[5079]),

			.O(gen[5172]),
			.E(gen[5174]),

			.SO(gen[5267]),
			.S(gen[5268]),
			.SE(gen[5269]),

			.SELF(gen[5173]),
			.cell_state(gen[5173])
		); 

/******************* CELL 5174 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5174 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5078]),
			.N(gen[5079]),
			.NE(gen[5080]),

			.O(gen[5173]),
			.E(gen[5175]),

			.SO(gen[5268]),
			.S(gen[5269]),
			.SE(gen[5270]),

			.SELF(gen[5174]),
			.cell_state(gen[5174])
		); 

/******************* CELL 5175 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5175 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5079]),
			.N(gen[5080]),
			.NE(gen[5081]),

			.O(gen[5174]),
			.E(gen[5176]),

			.SO(gen[5269]),
			.S(gen[5270]),
			.SE(gen[5271]),

			.SELF(gen[5175]),
			.cell_state(gen[5175])
		); 

/******************* CELL 5176 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5176 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5080]),
			.N(gen[5081]),
			.NE(gen[5082]),

			.O(gen[5175]),
			.E(gen[5177]),

			.SO(gen[5270]),
			.S(gen[5271]),
			.SE(gen[5272]),

			.SELF(gen[5176]),
			.cell_state(gen[5176])
		); 

/******************* CELL 5177 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5177 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5081]),
			.N(gen[5082]),
			.NE(gen[5083]),

			.O(gen[5176]),
			.E(gen[5178]),

			.SO(gen[5271]),
			.S(gen[5272]),
			.SE(gen[5273]),

			.SELF(gen[5177]),
			.cell_state(gen[5177])
		); 

/******************* CELL 5178 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5178 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5082]),
			.N(gen[5083]),
			.NE(gen[5084]),

			.O(gen[5177]),
			.E(gen[5179]),

			.SO(gen[5272]),
			.S(gen[5273]),
			.SE(gen[5274]),

			.SELF(gen[5178]),
			.cell_state(gen[5178])
		); 

/******************* CELL 5179 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5179 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5083]),
			.N(gen[5084]),
			.NE(gen[5085]),

			.O(gen[5178]),
			.E(gen[5180]),

			.SO(gen[5273]),
			.S(gen[5274]),
			.SE(gen[5275]),

			.SELF(gen[5179]),
			.cell_state(gen[5179])
		); 

/******************* CELL 5180 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5180 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5084]),
			.N(gen[5085]),
			.NE(gen[5086]),

			.O(gen[5179]),
			.E(gen[5181]),

			.SO(gen[5274]),
			.S(gen[5275]),
			.SE(gen[5276]),

			.SELF(gen[5180]),
			.cell_state(gen[5180])
		); 

/******************* CELL 5181 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5181 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5085]),
			.N(gen[5086]),
			.NE(gen[5087]),

			.O(gen[5180]),
			.E(gen[5182]),

			.SO(gen[5275]),
			.S(gen[5276]),
			.SE(gen[5277]),

			.SELF(gen[5181]),
			.cell_state(gen[5181])
		); 

/******************* CELL 5182 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5182 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5086]),
			.N(gen[5087]),
			.NE(gen[5088]),

			.O(gen[5181]),
			.E(gen[5183]),

			.SO(gen[5276]),
			.S(gen[5277]),
			.SE(gen[5278]),

			.SELF(gen[5182]),
			.cell_state(gen[5182])
		); 

/******************* CELL 5183 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5183 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5087]),
			.N(gen[5088]),
			.NE(gen[5089]),

			.O(gen[5182]),
			.E(gen[5184]),

			.SO(gen[5277]),
			.S(gen[5278]),
			.SE(gen[5279]),

			.SELF(gen[5183]),
			.cell_state(gen[5183])
		); 

/******************* CELL 5184 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5184 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5088]),
			.N(gen[5089]),
			.NE(gen[5090]),

			.O(gen[5183]),
			.E(gen[5185]),

			.SO(gen[5278]),
			.S(gen[5279]),
			.SE(gen[5280]),

			.SELF(gen[5184]),
			.cell_state(gen[5184])
		); 

/******************* CELL 5185 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5185 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5089]),
			.N(gen[5090]),
			.NE(gen[5091]),

			.O(gen[5184]),
			.E(gen[5186]),

			.SO(gen[5279]),
			.S(gen[5280]),
			.SE(gen[5281]),

			.SELF(gen[5185]),
			.cell_state(gen[5185])
		); 

/******************* CELL 5186 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5186 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5090]),
			.N(gen[5091]),
			.NE(gen[5092]),

			.O(gen[5185]),
			.E(gen[5187]),

			.SO(gen[5280]),
			.S(gen[5281]),
			.SE(gen[5282]),

			.SELF(gen[5186]),
			.cell_state(gen[5186])
		); 

/******************* CELL 5187 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5187 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5091]),
			.N(gen[5092]),
			.NE(gen[5093]),

			.O(gen[5186]),
			.E(gen[5188]),

			.SO(gen[5281]),
			.S(gen[5282]),
			.SE(gen[5283]),

			.SELF(gen[5187]),
			.cell_state(gen[5187])
		); 

/******************* CELL 5188 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5188 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5092]),
			.N(gen[5093]),
			.NE(gen[5094]),

			.O(gen[5187]),
			.E(gen[5189]),

			.SO(gen[5282]),
			.S(gen[5283]),
			.SE(gen[5284]),

			.SELF(gen[5188]),
			.cell_state(gen[5188])
		); 

/******************* CELL 5189 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5189 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5093]),
			.N(gen[5094]),
			.NE(gen[5095]),

			.O(gen[5188]),
			.E(gen[5190]),

			.SO(gen[5283]),
			.S(gen[5284]),
			.SE(gen[5285]),

			.SELF(gen[5189]),
			.cell_state(gen[5189])
		); 

/******************* CELL 5190 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5190 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5094]),
			.N(gen[5095]),
			.NE(gen[5096]),

			.O(gen[5189]),
			.E(gen[5191]),

			.SO(gen[5284]),
			.S(gen[5285]),
			.SE(gen[5286]),

			.SELF(gen[5190]),
			.cell_state(gen[5190])
		); 

/******************* CELL 5191 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5191 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5095]),
			.N(gen[5096]),
			.NE(gen[5097]),

			.O(gen[5190]),
			.E(gen[5192]),

			.SO(gen[5285]),
			.S(gen[5286]),
			.SE(gen[5287]),

			.SELF(gen[5191]),
			.cell_state(gen[5191])
		); 

/******************* CELL 5192 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5192 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5096]),
			.N(gen[5097]),
			.NE(gen[5098]),

			.O(gen[5191]),
			.E(gen[5193]),

			.SO(gen[5286]),
			.S(gen[5287]),
			.SE(gen[5288]),

			.SELF(gen[5192]),
			.cell_state(gen[5192])
		); 

/******************* CELL 5193 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5193 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5097]),
			.N(gen[5098]),
			.NE(gen[5099]),

			.O(gen[5192]),
			.E(gen[5194]),

			.SO(gen[5287]),
			.S(gen[5288]),
			.SE(gen[5289]),

			.SELF(gen[5193]),
			.cell_state(gen[5193])
		); 

/******************* CELL 5194 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5194 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5098]),
			.N(gen[5099]),
			.NE(gen[5100]),

			.O(gen[5193]),
			.E(gen[5195]),

			.SO(gen[5288]),
			.S(gen[5289]),
			.SE(gen[5290]),

			.SELF(gen[5194]),
			.cell_state(gen[5194])
		); 

/******************* CELL 5195 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5195 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5099]),
			.N(gen[5100]),
			.NE(gen[5101]),

			.O(gen[5194]),
			.E(gen[5196]),

			.SO(gen[5289]),
			.S(gen[5290]),
			.SE(gen[5291]),

			.SELF(gen[5195]),
			.cell_state(gen[5195])
		); 

/******************* CELL 5196 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5196 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5100]),
			.N(gen[5101]),
			.NE(gen[5102]),

			.O(gen[5195]),
			.E(gen[5197]),

			.SO(gen[5290]),
			.S(gen[5291]),
			.SE(gen[5292]),

			.SELF(gen[5196]),
			.cell_state(gen[5196])
		); 

/******************* CELL 5197 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5197 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5101]),
			.N(gen[5102]),
			.NE(gen[5103]),

			.O(gen[5196]),
			.E(gen[5198]),

			.SO(gen[5291]),
			.S(gen[5292]),
			.SE(gen[5293]),

			.SELF(gen[5197]),
			.cell_state(gen[5197])
		); 

/******************* CELL 5198 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5198 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5102]),
			.N(gen[5103]),
			.NE(gen[5104]),

			.O(gen[5197]),
			.E(gen[5199]),

			.SO(gen[5292]),
			.S(gen[5293]),
			.SE(gen[5294]),

			.SELF(gen[5198]),
			.cell_state(gen[5198])
		); 

/******************* CELL 5199 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5199 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5103]),
			.N(gen[5104]),
			.NE(gen[5105]),

			.O(gen[5198]),
			.E(gen[5200]),

			.SO(gen[5293]),
			.S(gen[5294]),
			.SE(gen[5295]),

			.SELF(gen[5199]),
			.cell_state(gen[5199])
		); 

/******************* CELL 5200 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5200 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5104]),
			.N(gen[5105]),
			.NE(gen[5106]),

			.O(gen[5199]),
			.E(gen[5201]),

			.SO(gen[5294]),
			.S(gen[5295]),
			.SE(gen[5296]),

			.SELF(gen[5200]),
			.cell_state(gen[5200])
		); 

/******************* CELL 5201 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5201 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5105]),
			.N(gen[5106]),
			.NE(gen[5107]),

			.O(gen[5200]),
			.E(gen[5202]),

			.SO(gen[5295]),
			.S(gen[5296]),
			.SE(gen[5297]),

			.SELF(gen[5201]),
			.cell_state(gen[5201])
		); 

/******************* CELL 5202 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5202 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5106]),
			.N(gen[5107]),
			.NE(gen[5108]),

			.O(gen[5201]),
			.E(gen[5203]),

			.SO(gen[5296]),
			.S(gen[5297]),
			.SE(gen[5298]),

			.SELF(gen[5202]),
			.cell_state(gen[5202])
		); 

/******************* CELL 5203 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5203 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5107]),
			.N(gen[5108]),
			.NE(gen[5109]),

			.O(gen[5202]),
			.E(gen[5204]),

			.SO(gen[5297]),
			.S(gen[5298]),
			.SE(gen[5299]),

			.SELF(gen[5203]),
			.cell_state(gen[5203])
		); 

/******************* CELL 5204 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5204 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5108]),
			.N(gen[5109]),
			.NE(gen[5110]),

			.O(gen[5203]),
			.E(gen[5205]),

			.SO(gen[5298]),
			.S(gen[5299]),
			.SE(gen[5300]),

			.SELF(gen[5204]),
			.cell_state(gen[5204])
		); 

/******************* CELL 5205 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5205 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5109]),
			.N(gen[5110]),
			.NE(gen[5111]),

			.O(gen[5204]),
			.E(gen[5206]),

			.SO(gen[5299]),
			.S(gen[5300]),
			.SE(gen[5301]),

			.SELF(gen[5205]),
			.cell_state(gen[5205])
		); 

/******************* CELL 5206 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5206 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5110]),
			.N(gen[5111]),
			.NE(gen[5112]),

			.O(gen[5205]),
			.E(gen[5207]),

			.SO(gen[5300]),
			.S(gen[5301]),
			.SE(gen[5302]),

			.SELF(gen[5206]),
			.cell_state(gen[5206])
		); 

/******************* CELL 5207 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5207 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5111]),
			.N(gen[5112]),
			.NE(gen[5113]),

			.O(gen[5206]),
			.E(gen[5208]),

			.SO(gen[5301]),
			.S(gen[5302]),
			.SE(gen[5303]),

			.SELF(gen[5207]),
			.cell_state(gen[5207])
		); 

/******************* CELL 5208 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5208 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5112]),
			.N(gen[5113]),
			.NE(gen[5114]),

			.O(gen[5207]),
			.E(gen[5209]),

			.SO(gen[5302]),
			.S(gen[5303]),
			.SE(gen[5304]),

			.SELF(gen[5208]),
			.cell_state(gen[5208])
		); 

/******************* CELL 5209 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5209 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5113]),
			.N(gen[5114]),
			.NE(gen[5115]),

			.O(gen[5208]),
			.E(gen[5210]),

			.SO(gen[5303]),
			.S(gen[5304]),
			.SE(gen[5305]),

			.SELF(gen[5209]),
			.cell_state(gen[5209])
		); 

/******************* CELL 5210 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5210 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5114]),
			.N(gen[5115]),
			.NE(gen[5116]),

			.O(gen[5209]),
			.E(gen[5211]),

			.SO(gen[5304]),
			.S(gen[5305]),
			.SE(gen[5306]),

			.SELF(gen[5210]),
			.cell_state(gen[5210])
		); 

/******************* CELL 5211 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5211 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5115]),
			.N(gen[5116]),
			.NE(gen[5117]),

			.O(gen[5210]),
			.E(gen[5212]),

			.SO(gen[5305]),
			.S(gen[5306]),
			.SE(gen[5307]),

			.SELF(gen[5211]),
			.cell_state(gen[5211])
		); 

/******************* CELL 5212 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5212 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5116]),
			.N(gen[5117]),
			.NE(gen[5118]),

			.O(gen[5211]),
			.E(gen[5213]),

			.SO(gen[5306]),
			.S(gen[5307]),
			.SE(gen[5308]),

			.SELF(gen[5212]),
			.cell_state(gen[5212])
		); 

/******************* CELL 5213 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5213 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5117]),
			.N(gen[5118]),
			.NE(gen[5119]),

			.O(gen[5212]),
			.E(gen[5214]),

			.SO(gen[5307]),
			.S(gen[5308]),
			.SE(gen[5309]),

			.SELF(gen[5213]),
			.cell_state(gen[5213])
		); 

/******************* CELL 5214 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5214 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5118]),
			.N(gen[5119]),
			.NE(gen[5120]),

			.O(gen[5213]),
			.E(gen[5215]),

			.SO(gen[5308]),
			.S(gen[5309]),
			.SE(gen[5310]),

			.SELF(gen[5214]),
			.cell_state(gen[5214])
		); 

/******************* CELL 5215 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5215 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5119]),
			.N(gen[5120]),
			.NE(gen[5121]),

			.O(gen[5214]),
			.E(gen[5216]),

			.SO(gen[5309]),
			.S(gen[5310]),
			.SE(gen[5311]),

			.SELF(gen[5215]),
			.cell_state(gen[5215])
		); 

/******************* CELL 5216 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5216 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5120]),
			.N(gen[5121]),
			.NE(gen[5122]),

			.O(gen[5215]),
			.E(gen[5217]),

			.SO(gen[5310]),
			.S(gen[5311]),
			.SE(gen[5312]),

			.SELF(gen[5216]),
			.cell_state(gen[5216])
		); 

/******************* CELL 5217 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5217 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5121]),
			.N(gen[5122]),
			.NE(gen[5123]),

			.O(gen[5216]),
			.E(gen[5218]),

			.SO(gen[5311]),
			.S(gen[5312]),
			.SE(gen[5313]),

			.SELF(gen[5217]),
			.cell_state(gen[5217])
		); 

/******************* CELL 5218 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5218 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5122]),
			.N(gen[5123]),
			.NE(gen[5124]),

			.O(gen[5217]),
			.E(gen[5219]),

			.SO(gen[5312]),
			.S(gen[5313]),
			.SE(gen[5314]),

			.SELF(gen[5218]),
			.cell_state(gen[5218])
		); 

/******************* CELL 5219 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5219 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5123]),
			.N(gen[5124]),
			.NE(gen[5125]),

			.O(gen[5218]),
			.E(gen[5220]),

			.SO(gen[5313]),
			.S(gen[5314]),
			.SE(gen[5315]),

			.SELF(gen[5219]),
			.cell_state(gen[5219])
		); 

/******************* CELL 5220 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5220 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5124]),
			.N(gen[5125]),
			.NE(gen[5126]),

			.O(gen[5219]),
			.E(gen[5221]),

			.SO(gen[5314]),
			.S(gen[5315]),
			.SE(gen[5316]),

			.SELF(gen[5220]),
			.cell_state(gen[5220])
		); 

/******************* CELL 5221 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5221 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5125]),
			.N(gen[5126]),
			.NE(gen[5127]),

			.O(gen[5220]),
			.E(gen[5222]),

			.SO(gen[5315]),
			.S(gen[5316]),
			.SE(gen[5317]),

			.SELF(gen[5221]),
			.cell_state(gen[5221])
		); 

/******************* CELL 5222 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5222 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5126]),
			.N(gen[5127]),
			.NE(gen[5128]),

			.O(gen[5221]),
			.E(gen[5223]),

			.SO(gen[5316]),
			.S(gen[5317]),
			.SE(gen[5318]),

			.SELF(gen[5222]),
			.cell_state(gen[5222])
		); 

/******************* CELL 5223 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5223 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5127]),
			.N(gen[5128]),
			.NE(gen[5129]),

			.O(gen[5222]),
			.E(gen[5224]),

			.SO(gen[5317]),
			.S(gen[5318]),
			.SE(gen[5319]),

			.SELF(gen[5223]),
			.cell_state(gen[5223])
		); 

/******************* CELL 5224 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5224 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5128]),
			.N(gen[5129]),
			.NE(gen[5128]),

			.O(gen[5223]),
			.E(gen[5223]),

			.SO(gen[5318]),
			.S(gen[5319]),
			.SE(gen[5318]),

			.SELF(gen[5224]),
			.cell_state(gen[5224])
		); 

/******************* CELL 5225 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5225 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5131]),
			.N(gen[5130]),
			.NE(gen[5131]),

			.O(gen[5226]),
			.E(gen[5226]),

			.SO(gen[5321]),
			.S(gen[5320]),
			.SE(gen[5321]),

			.SELF(gen[5225]),
			.cell_state(gen[5225])
		); 

/******************* CELL 5226 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5226 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5130]),
			.N(gen[5131]),
			.NE(gen[5132]),

			.O(gen[5225]),
			.E(gen[5227]),

			.SO(gen[5320]),
			.S(gen[5321]),
			.SE(gen[5322]),

			.SELF(gen[5226]),
			.cell_state(gen[5226])
		); 

/******************* CELL 5227 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5227 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5131]),
			.N(gen[5132]),
			.NE(gen[5133]),

			.O(gen[5226]),
			.E(gen[5228]),

			.SO(gen[5321]),
			.S(gen[5322]),
			.SE(gen[5323]),

			.SELF(gen[5227]),
			.cell_state(gen[5227])
		); 

/******************* CELL 5228 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5228 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5132]),
			.N(gen[5133]),
			.NE(gen[5134]),

			.O(gen[5227]),
			.E(gen[5229]),

			.SO(gen[5322]),
			.S(gen[5323]),
			.SE(gen[5324]),

			.SELF(gen[5228]),
			.cell_state(gen[5228])
		); 

/******************* CELL 5229 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5229 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5133]),
			.N(gen[5134]),
			.NE(gen[5135]),

			.O(gen[5228]),
			.E(gen[5230]),

			.SO(gen[5323]),
			.S(gen[5324]),
			.SE(gen[5325]),

			.SELF(gen[5229]),
			.cell_state(gen[5229])
		); 

/******************* CELL 5230 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5230 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5134]),
			.N(gen[5135]),
			.NE(gen[5136]),

			.O(gen[5229]),
			.E(gen[5231]),

			.SO(gen[5324]),
			.S(gen[5325]),
			.SE(gen[5326]),

			.SELF(gen[5230]),
			.cell_state(gen[5230])
		); 

/******************* CELL 5231 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5231 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5135]),
			.N(gen[5136]),
			.NE(gen[5137]),

			.O(gen[5230]),
			.E(gen[5232]),

			.SO(gen[5325]),
			.S(gen[5326]),
			.SE(gen[5327]),

			.SELF(gen[5231]),
			.cell_state(gen[5231])
		); 

/******************* CELL 5232 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5232 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5136]),
			.N(gen[5137]),
			.NE(gen[5138]),

			.O(gen[5231]),
			.E(gen[5233]),

			.SO(gen[5326]),
			.S(gen[5327]),
			.SE(gen[5328]),

			.SELF(gen[5232]),
			.cell_state(gen[5232])
		); 

/******************* CELL 5233 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5233 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5137]),
			.N(gen[5138]),
			.NE(gen[5139]),

			.O(gen[5232]),
			.E(gen[5234]),

			.SO(gen[5327]),
			.S(gen[5328]),
			.SE(gen[5329]),

			.SELF(gen[5233]),
			.cell_state(gen[5233])
		); 

/******************* CELL 5234 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5234 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5138]),
			.N(gen[5139]),
			.NE(gen[5140]),

			.O(gen[5233]),
			.E(gen[5235]),

			.SO(gen[5328]),
			.S(gen[5329]),
			.SE(gen[5330]),

			.SELF(gen[5234]),
			.cell_state(gen[5234])
		); 

/******************* CELL 5235 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5235 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5139]),
			.N(gen[5140]),
			.NE(gen[5141]),

			.O(gen[5234]),
			.E(gen[5236]),

			.SO(gen[5329]),
			.S(gen[5330]),
			.SE(gen[5331]),

			.SELF(gen[5235]),
			.cell_state(gen[5235])
		); 

/******************* CELL 5236 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5236 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5140]),
			.N(gen[5141]),
			.NE(gen[5142]),

			.O(gen[5235]),
			.E(gen[5237]),

			.SO(gen[5330]),
			.S(gen[5331]),
			.SE(gen[5332]),

			.SELF(gen[5236]),
			.cell_state(gen[5236])
		); 

/******************* CELL 5237 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5237 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5141]),
			.N(gen[5142]),
			.NE(gen[5143]),

			.O(gen[5236]),
			.E(gen[5238]),

			.SO(gen[5331]),
			.S(gen[5332]),
			.SE(gen[5333]),

			.SELF(gen[5237]),
			.cell_state(gen[5237])
		); 

/******************* CELL 5238 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5238 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5142]),
			.N(gen[5143]),
			.NE(gen[5144]),

			.O(gen[5237]),
			.E(gen[5239]),

			.SO(gen[5332]),
			.S(gen[5333]),
			.SE(gen[5334]),

			.SELF(gen[5238]),
			.cell_state(gen[5238])
		); 

/******************* CELL 5239 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5239 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5143]),
			.N(gen[5144]),
			.NE(gen[5145]),

			.O(gen[5238]),
			.E(gen[5240]),

			.SO(gen[5333]),
			.S(gen[5334]),
			.SE(gen[5335]),

			.SELF(gen[5239]),
			.cell_state(gen[5239])
		); 

/******************* CELL 5240 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5240 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5144]),
			.N(gen[5145]),
			.NE(gen[5146]),

			.O(gen[5239]),
			.E(gen[5241]),

			.SO(gen[5334]),
			.S(gen[5335]),
			.SE(gen[5336]),

			.SELF(gen[5240]),
			.cell_state(gen[5240])
		); 

/******************* CELL 5241 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5241 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5145]),
			.N(gen[5146]),
			.NE(gen[5147]),

			.O(gen[5240]),
			.E(gen[5242]),

			.SO(gen[5335]),
			.S(gen[5336]),
			.SE(gen[5337]),

			.SELF(gen[5241]),
			.cell_state(gen[5241])
		); 

/******************* CELL 5242 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5242 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5146]),
			.N(gen[5147]),
			.NE(gen[5148]),

			.O(gen[5241]),
			.E(gen[5243]),

			.SO(gen[5336]),
			.S(gen[5337]),
			.SE(gen[5338]),

			.SELF(gen[5242]),
			.cell_state(gen[5242])
		); 

/******************* CELL 5243 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5243 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5147]),
			.N(gen[5148]),
			.NE(gen[5149]),

			.O(gen[5242]),
			.E(gen[5244]),

			.SO(gen[5337]),
			.S(gen[5338]),
			.SE(gen[5339]),

			.SELF(gen[5243]),
			.cell_state(gen[5243])
		); 

/******************* CELL 5244 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5244 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5148]),
			.N(gen[5149]),
			.NE(gen[5150]),

			.O(gen[5243]),
			.E(gen[5245]),

			.SO(gen[5338]),
			.S(gen[5339]),
			.SE(gen[5340]),

			.SELF(gen[5244]),
			.cell_state(gen[5244])
		); 

/******************* CELL 5245 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5245 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5149]),
			.N(gen[5150]),
			.NE(gen[5151]),

			.O(gen[5244]),
			.E(gen[5246]),

			.SO(gen[5339]),
			.S(gen[5340]),
			.SE(gen[5341]),

			.SELF(gen[5245]),
			.cell_state(gen[5245])
		); 

/******************* CELL 5246 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5246 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5150]),
			.N(gen[5151]),
			.NE(gen[5152]),

			.O(gen[5245]),
			.E(gen[5247]),

			.SO(gen[5340]),
			.S(gen[5341]),
			.SE(gen[5342]),

			.SELF(gen[5246]),
			.cell_state(gen[5246])
		); 

/******************* CELL 5247 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5247 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5151]),
			.N(gen[5152]),
			.NE(gen[5153]),

			.O(gen[5246]),
			.E(gen[5248]),

			.SO(gen[5341]),
			.S(gen[5342]),
			.SE(gen[5343]),

			.SELF(gen[5247]),
			.cell_state(gen[5247])
		); 

/******************* CELL 5248 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5248 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5152]),
			.N(gen[5153]),
			.NE(gen[5154]),

			.O(gen[5247]),
			.E(gen[5249]),

			.SO(gen[5342]),
			.S(gen[5343]),
			.SE(gen[5344]),

			.SELF(gen[5248]),
			.cell_state(gen[5248])
		); 

/******************* CELL 5249 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5249 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5153]),
			.N(gen[5154]),
			.NE(gen[5155]),

			.O(gen[5248]),
			.E(gen[5250]),

			.SO(gen[5343]),
			.S(gen[5344]),
			.SE(gen[5345]),

			.SELF(gen[5249]),
			.cell_state(gen[5249])
		); 

/******************* CELL 5250 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5250 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5154]),
			.N(gen[5155]),
			.NE(gen[5156]),

			.O(gen[5249]),
			.E(gen[5251]),

			.SO(gen[5344]),
			.S(gen[5345]),
			.SE(gen[5346]),

			.SELF(gen[5250]),
			.cell_state(gen[5250])
		); 

/******************* CELL 5251 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5251 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5155]),
			.N(gen[5156]),
			.NE(gen[5157]),

			.O(gen[5250]),
			.E(gen[5252]),

			.SO(gen[5345]),
			.S(gen[5346]),
			.SE(gen[5347]),

			.SELF(gen[5251]),
			.cell_state(gen[5251])
		); 

/******************* CELL 5252 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5252 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5156]),
			.N(gen[5157]),
			.NE(gen[5158]),

			.O(gen[5251]),
			.E(gen[5253]),

			.SO(gen[5346]),
			.S(gen[5347]),
			.SE(gen[5348]),

			.SELF(gen[5252]),
			.cell_state(gen[5252])
		); 

/******************* CELL 5253 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5253 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5157]),
			.N(gen[5158]),
			.NE(gen[5159]),

			.O(gen[5252]),
			.E(gen[5254]),

			.SO(gen[5347]),
			.S(gen[5348]),
			.SE(gen[5349]),

			.SELF(gen[5253]),
			.cell_state(gen[5253])
		); 

/******************* CELL 5254 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5254 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5158]),
			.N(gen[5159]),
			.NE(gen[5160]),

			.O(gen[5253]),
			.E(gen[5255]),

			.SO(gen[5348]),
			.S(gen[5349]),
			.SE(gen[5350]),

			.SELF(gen[5254]),
			.cell_state(gen[5254])
		); 

/******************* CELL 5255 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5255 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5159]),
			.N(gen[5160]),
			.NE(gen[5161]),

			.O(gen[5254]),
			.E(gen[5256]),

			.SO(gen[5349]),
			.S(gen[5350]),
			.SE(gen[5351]),

			.SELF(gen[5255]),
			.cell_state(gen[5255])
		); 

/******************* CELL 5256 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5256 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5160]),
			.N(gen[5161]),
			.NE(gen[5162]),

			.O(gen[5255]),
			.E(gen[5257]),

			.SO(gen[5350]),
			.S(gen[5351]),
			.SE(gen[5352]),

			.SELF(gen[5256]),
			.cell_state(gen[5256])
		); 

/******************* CELL 5257 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5257 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5161]),
			.N(gen[5162]),
			.NE(gen[5163]),

			.O(gen[5256]),
			.E(gen[5258]),

			.SO(gen[5351]),
			.S(gen[5352]),
			.SE(gen[5353]),

			.SELF(gen[5257]),
			.cell_state(gen[5257])
		); 

/******************* CELL 5258 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5258 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5162]),
			.N(gen[5163]),
			.NE(gen[5164]),

			.O(gen[5257]),
			.E(gen[5259]),

			.SO(gen[5352]),
			.S(gen[5353]),
			.SE(gen[5354]),

			.SELF(gen[5258]),
			.cell_state(gen[5258])
		); 

/******************* CELL 5259 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5259 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5163]),
			.N(gen[5164]),
			.NE(gen[5165]),

			.O(gen[5258]),
			.E(gen[5260]),

			.SO(gen[5353]),
			.S(gen[5354]),
			.SE(gen[5355]),

			.SELF(gen[5259]),
			.cell_state(gen[5259])
		); 

/******************* CELL 5260 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5260 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5164]),
			.N(gen[5165]),
			.NE(gen[5166]),

			.O(gen[5259]),
			.E(gen[5261]),

			.SO(gen[5354]),
			.S(gen[5355]),
			.SE(gen[5356]),

			.SELF(gen[5260]),
			.cell_state(gen[5260])
		); 

/******************* CELL 5261 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5261 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5165]),
			.N(gen[5166]),
			.NE(gen[5167]),

			.O(gen[5260]),
			.E(gen[5262]),

			.SO(gen[5355]),
			.S(gen[5356]),
			.SE(gen[5357]),

			.SELF(gen[5261]),
			.cell_state(gen[5261])
		); 

/******************* CELL 5262 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5262 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5166]),
			.N(gen[5167]),
			.NE(gen[5168]),

			.O(gen[5261]),
			.E(gen[5263]),

			.SO(gen[5356]),
			.S(gen[5357]),
			.SE(gen[5358]),

			.SELF(gen[5262]),
			.cell_state(gen[5262])
		); 

/******************* CELL 5263 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5263 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5167]),
			.N(gen[5168]),
			.NE(gen[5169]),

			.O(gen[5262]),
			.E(gen[5264]),

			.SO(gen[5357]),
			.S(gen[5358]),
			.SE(gen[5359]),

			.SELF(gen[5263]),
			.cell_state(gen[5263])
		); 

/******************* CELL 5264 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5264 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5168]),
			.N(gen[5169]),
			.NE(gen[5170]),

			.O(gen[5263]),
			.E(gen[5265]),

			.SO(gen[5358]),
			.S(gen[5359]),
			.SE(gen[5360]),

			.SELF(gen[5264]),
			.cell_state(gen[5264])
		); 

/******************* CELL 5265 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5265 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5169]),
			.N(gen[5170]),
			.NE(gen[5171]),

			.O(gen[5264]),
			.E(gen[5266]),

			.SO(gen[5359]),
			.S(gen[5360]),
			.SE(gen[5361]),

			.SELF(gen[5265]),
			.cell_state(gen[5265])
		); 

/******************* CELL 5266 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5266 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5170]),
			.N(gen[5171]),
			.NE(gen[5172]),

			.O(gen[5265]),
			.E(gen[5267]),

			.SO(gen[5360]),
			.S(gen[5361]),
			.SE(gen[5362]),

			.SELF(gen[5266]),
			.cell_state(gen[5266])
		); 

/******************* CELL 5267 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5267 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5171]),
			.N(gen[5172]),
			.NE(gen[5173]),

			.O(gen[5266]),
			.E(gen[5268]),

			.SO(gen[5361]),
			.S(gen[5362]),
			.SE(gen[5363]),

			.SELF(gen[5267]),
			.cell_state(gen[5267])
		); 

/******************* CELL 5268 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5268 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5172]),
			.N(gen[5173]),
			.NE(gen[5174]),

			.O(gen[5267]),
			.E(gen[5269]),

			.SO(gen[5362]),
			.S(gen[5363]),
			.SE(gen[5364]),

			.SELF(gen[5268]),
			.cell_state(gen[5268])
		); 

/******************* CELL 5269 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5269 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5173]),
			.N(gen[5174]),
			.NE(gen[5175]),

			.O(gen[5268]),
			.E(gen[5270]),

			.SO(gen[5363]),
			.S(gen[5364]),
			.SE(gen[5365]),

			.SELF(gen[5269]),
			.cell_state(gen[5269])
		); 

/******************* CELL 5270 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5270 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5174]),
			.N(gen[5175]),
			.NE(gen[5176]),

			.O(gen[5269]),
			.E(gen[5271]),

			.SO(gen[5364]),
			.S(gen[5365]),
			.SE(gen[5366]),

			.SELF(gen[5270]),
			.cell_state(gen[5270])
		); 

/******************* CELL 5271 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5271 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5175]),
			.N(gen[5176]),
			.NE(gen[5177]),

			.O(gen[5270]),
			.E(gen[5272]),

			.SO(gen[5365]),
			.S(gen[5366]),
			.SE(gen[5367]),

			.SELF(gen[5271]),
			.cell_state(gen[5271])
		); 

/******************* CELL 5272 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5272 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5176]),
			.N(gen[5177]),
			.NE(gen[5178]),

			.O(gen[5271]),
			.E(gen[5273]),

			.SO(gen[5366]),
			.S(gen[5367]),
			.SE(gen[5368]),

			.SELF(gen[5272]),
			.cell_state(gen[5272])
		); 

/******************* CELL 5273 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5273 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5177]),
			.N(gen[5178]),
			.NE(gen[5179]),

			.O(gen[5272]),
			.E(gen[5274]),

			.SO(gen[5367]),
			.S(gen[5368]),
			.SE(gen[5369]),

			.SELF(gen[5273]),
			.cell_state(gen[5273])
		); 

/******************* CELL 5274 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5274 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5178]),
			.N(gen[5179]),
			.NE(gen[5180]),

			.O(gen[5273]),
			.E(gen[5275]),

			.SO(gen[5368]),
			.S(gen[5369]),
			.SE(gen[5370]),

			.SELF(gen[5274]),
			.cell_state(gen[5274])
		); 

/******************* CELL 5275 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5275 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5179]),
			.N(gen[5180]),
			.NE(gen[5181]),

			.O(gen[5274]),
			.E(gen[5276]),

			.SO(gen[5369]),
			.S(gen[5370]),
			.SE(gen[5371]),

			.SELF(gen[5275]),
			.cell_state(gen[5275])
		); 

/******************* CELL 5276 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5276 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5180]),
			.N(gen[5181]),
			.NE(gen[5182]),

			.O(gen[5275]),
			.E(gen[5277]),

			.SO(gen[5370]),
			.S(gen[5371]),
			.SE(gen[5372]),

			.SELF(gen[5276]),
			.cell_state(gen[5276])
		); 

/******************* CELL 5277 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5277 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5181]),
			.N(gen[5182]),
			.NE(gen[5183]),

			.O(gen[5276]),
			.E(gen[5278]),

			.SO(gen[5371]),
			.S(gen[5372]),
			.SE(gen[5373]),

			.SELF(gen[5277]),
			.cell_state(gen[5277])
		); 

/******************* CELL 5278 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5278 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5182]),
			.N(gen[5183]),
			.NE(gen[5184]),

			.O(gen[5277]),
			.E(gen[5279]),

			.SO(gen[5372]),
			.S(gen[5373]),
			.SE(gen[5374]),

			.SELF(gen[5278]),
			.cell_state(gen[5278])
		); 

/******************* CELL 5279 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5279 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5183]),
			.N(gen[5184]),
			.NE(gen[5185]),

			.O(gen[5278]),
			.E(gen[5280]),

			.SO(gen[5373]),
			.S(gen[5374]),
			.SE(gen[5375]),

			.SELF(gen[5279]),
			.cell_state(gen[5279])
		); 

/******************* CELL 5280 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5280 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5184]),
			.N(gen[5185]),
			.NE(gen[5186]),

			.O(gen[5279]),
			.E(gen[5281]),

			.SO(gen[5374]),
			.S(gen[5375]),
			.SE(gen[5376]),

			.SELF(gen[5280]),
			.cell_state(gen[5280])
		); 

/******************* CELL 5281 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5281 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5185]),
			.N(gen[5186]),
			.NE(gen[5187]),

			.O(gen[5280]),
			.E(gen[5282]),

			.SO(gen[5375]),
			.S(gen[5376]),
			.SE(gen[5377]),

			.SELF(gen[5281]),
			.cell_state(gen[5281])
		); 

/******************* CELL 5282 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5282 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5186]),
			.N(gen[5187]),
			.NE(gen[5188]),

			.O(gen[5281]),
			.E(gen[5283]),

			.SO(gen[5376]),
			.S(gen[5377]),
			.SE(gen[5378]),

			.SELF(gen[5282]),
			.cell_state(gen[5282])
		); 

/******************* CELL 5283 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5283 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5187]),
			.N(gen[5188]),
			.NE(gen[5189]),

			.O(gen[5282]),
			.E(gen[5284]),

			.SO(gen[5377]),
			.S(gen[5378]),
			.SE(gen[5379]),

			.SELF(gen[5283]),
			.cell_state(gen[5283])
		); 

/******************* CELL 5284 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5284 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5188]),
			.N(gen[5189]),
			.NE(gen[5190]),

			.O(gen[5283]),
			.E(gen[5285]),

			.SO(gen[5378]),
			.S(gen[5379]),
			.SE(gen[5380]),

			.SELF(gen[5284]),
			.cell_state(gen[5284])
		); 

/******************* CELL 5285 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5285 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5189]),
			.N(gen[5190]),
			.NE(gen[5191]),

			.O(gen[5284]),
			.E(gen[5286]),

			.SO(gen[5379]),
			.S(gen[5380]),
			.SE(gen[5381]),

			.SELF(gen[5285]),
			.cell_state(gen[5285])
		); 

/******************* CELL 5286 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5286 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5190]),
			.N(gen[5191]),
			.NE(gen[5192]),

			.O(gen[5285]),
			.E(gen[5287]),

			.SO(gen[5380]),
			.S(gen[5381]),
			.SE(gen[5382]),

			.SELF(gen[5286]),
			.cell_state(gen[5286])
		); 

/******************* CELL 5287 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5287 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5191]),
			.N(gen[5192]),
			.NE(gen[5193]),

			.O(gen[5286]),
			.E(gen[5288]),

			.SO(gen[5381]),
			.S(gen[5382]),
			.SE(gen[5383]),

			.SELF(gen[5287]),
			.cell_state(gen[5287])
		); 

/******************* CELL 5288 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5288 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5192]),
			.N(gen[5193]),
			.NE(gen[5194]),

			.O(gen[5287]),
			.E(gen[5289]),

			.SO(gen[5382]),
			.S(gen[5383]),
			.SE(gen[5384]),

			.SELF(gen[5288]),
			.cell_state(gen[5288])
		); 

/******************* CELL 5289 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5289 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5193]),
			.N(gen[5194]),
			.NE(gen[5195]),

			.O(gen[5288]),
			.E(gen[5290]),

			.SO(gen[5383]),
			.S(gen[5384]),
			.SE(gen[5385]),

			.SELF(gen[5289]),
			.cell_state(gen[5289])
		); 

/******************* CELL 5290 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5290 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5194]),
			.N(gen[5195]),
			.NE(gen[5196]),

			.O(gen[5289]),
			.E(gen[5291]),

			.SO(gen[5384]),
			.S(gen[5385]),
			.SE(gen[5386]),

			.SELF(gen[5290]),
			.cell_state(gen[5290])
		); 

/******************* CELL 5291 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5291 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5195]),
			.N(gen[5196]),
			.NE(gen[5197]),

			.O(gen[5290]),
			.E(gen[5292]),

			.SO(gen[5385]),
			.S(gen[5386]),
			.SE(gen[5387]),

			.SELF(gen[5291]),
			.cell_state(gen[5291])
		); 

/******************* CELL 5292 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5292 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5196]),
			.N(gen[5197]),
			.NE(gen[5198]),

			.O(gen[5291]),
			.E(gen[5293]),

			.SO(gen[5386]),
			.S(gen[5387]),
			.SE(gen[5388]),

			.SELF(gen[5292]),
			.cell_state(gen[5292])
		); 

/******************* CELL 5293 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5293 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5197]),
			.N(gen[5198]),
			.NE(gen[5199]),

			.O(gen[5292]),
			.E(gen[5294]),

			.SO(gen[5387]),
			.S(gen[5388]),
			.SE(gen[5389]),

			.SELF(gen[5293]),
			.cell_state(gen[5293])
		); 

/******************* CELL 5294 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5294 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5198]),
			.N(gen[5199]),
			.NE(gen[5200]),

			.O(gen[5293]),
			.E(gen[5295]),

			.SO(gen[5388]),
			.S(gen[5389]),
			.SE(gen[5390]),

			.SELF(gen[5294]),
			.cell_state(gen[5294])
		); 

/******************* CELL 5295 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5295 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5199]),
			.N(gen[5200]),
			.NE(gen[5201]),

			.O(gen[5294]),
			.E(gen[5296]),

			.SO(gen[5389]),
			.S(gen[5390]),
			.SE(gen[5391]),

			.SELF(gen[5295]),
			.cell_state(gen[5295])
		); 

/******************* CELL 5296 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5296 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5200]),
			.N(gen[5201]),
			.NE(gen[5202]),

			.O(gen[5295]),
			.E(gen[5297]),

			.SO(gen[5390]),
			.S(gen[5391]),
			.SE(gen[5392]),

			.SELF(gen[5296]),
			.cell_state(gen[5296])
		); 

/******************* CELL 5297 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5297 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5201]),
			.N(gen[5202]),
			.NE(gen[5203]),

			.O(gen[5296]),
			.E(gen[5298]),

			.SO(gen[5391]),
			.S(gen[5392]),
			.SE(gen[5393]),

			.SELF(gen[5297]),
			.cell_state(gen[5297])
		); 

/******************* CELL 5298 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5298 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5202]),
			.N(gen[5203]),
			.NE(gen[5204]),

			.O(gen[5297]),
			.E(gen[5299]),

			.SO(gen[5392]),
			.S(gen[5393]),
			.SE(gen[5394]),

			.SELF(gen[5298]),
			.cell_state(gen[5298])
		); 

/******************* CELL 5299 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5299 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5203]),
			.N(gen[5204]),
			.NE(gen[5205]),

			.O(gen[5298]),
			.E(gen[5300]),

			.SO(gen[5393]),
			.S(gen[5394]),
			.SE(gen[5395]),

			.SELF(gen[5299]),
			.cell_state(gen[5299])
		); 

/******************* CELL 5300 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5300 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5204]),
			.N(gen[5205]),
			.NE(gen[5206]),

			.O(gen[5299]),
			.E(gen[5301]),

			.SO(gen[5394]),
			.S(gen[5395]),
			.SE(gen[5396]),

			.SELF(gen[5300]),
			.cell_state(gen[5300])
		); 

/******************* CELL 5301 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5301 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5205]),
			.N(gen[5206]),
			.NE(gen[5207]),

			.O(gen[5300]),
			.E(gen[5302]),

			.SO(gen[5395]),
			.S(gen[5396]),
			.SE(gen[5397]),

			.SELF(gen[5301]),
			.cell_state(gen[5301])
		); 

/******************* CELL 5302 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5302 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5206]),
			.N(gen[5207]),
			.NE(gen[5208]),

			.O(gen[5301]),
			.E(gen[5303]),

			.SO(gen[5396]),
			.S(gen[5397]),
			.SE(gen[5398]),

			.SELF(gen[5302]),
			.cell_state(gen[5302])
		); 

/******************* CELL 5303 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5303 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5207]),
			.N(gen[5208]),
			.NE(gen[5209]),

			.O(gen[5302]),
			.E(gen[5304]),

			.SO(gen[5397]),
			.S(gen[5398]),
			.SE(gen[5399]),

			.SELF(gen[5303]),
			.cell_state(gen[5303])
		); 

/******************* CELL 5304 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5304 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5208]),
			.N(gen[5209]),
			.NE(gen[5210]),

			.O(gen[5303]),
			.E(gen[5305]),

			.SO(gen[5398]),
			.S(gen[5399]),
			.SE(gen[5400]),

			.SELF(gen[5304]),
			.cell_state(gen[5304])
		); 

/******************* CELL 5305 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5305 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5209]),
			.N(gen[5210]),
			.NE(gen[5211]),

			.O(gen[5304]),
			.E(gen[5306]),

			.SO(gen[5399]),
			.S(gen[5400]),
			.SE(gen[5401]),

			.SELF(gen[5305]),
			.cell_state(gen[5305])
		); 

/******************* CELL 5306 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5306 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5210]),
			.N(gen[5211]),
			.NE(gen[5212]),

			.O(gen[5305]),
			.E(gen[5307]),

			.SO(gen[5400]),
			.S(gen[5401]),
			.SE(gen[5402]),

			.SELF(gen[5306]),
			.cell_state(gen[5306])
		); 

/******************* CELL 5307 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5307 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5211]),
			.N(gen[5212]),
			.NE(gen[5213]),

			.O(gen[5306]),
			.E(gen[5308]),

			.SO(gen[5401]),
			.S(gen[5402]),
			.SE(gen[5403]),

			.SELF(gen[5307]),
			.cell_state(gen[5307])
		); 

/******************* CELL 5308 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5308 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5212]),
			.N(gen[5213]),
			.NE(gen[5214]),

			.O(gen[5307]),
			.E(gen[5309]),

			.SO(gen[5402]),
			.S(gen[5403]),
			.SE(gen[5404]),

			.SELF(gen[5308]),
			.cell_state(gen[5308])
		); 

/******************* CELL 5309 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5309 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5213]),
			.N(gen[5214]),
			.NE(gen[5215]),

			.O(gen[5308]),
			.E(gen[5310]),

			.SO(gen[5403]),
			.S(gen[5404]),
			.SE(gen[5405]),

			.SELF(gen[5309]),
			.cell_state(gen[5309])
		); 

/******************* CELL 5310 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5310 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5214]),
			.N(gen[5215]),
			.NE(gen[5216]),

			.O(gen[5309]),
			.E(gen[5311]),

			.SO(gen[5404]),
			.S(gen[5405]),
			.SE(gen[5406]),

			.SELF(gen[5310]),
			.cell_state(gen[5310])
		); 

/******************* CELL 5311 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5311 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5215]),
			.N(gen[5216]),
			.NE(gen[5217]),

			.O(gen[5310]),
			.E(gen[5312]),

			.SO(gen[5405]),
			.S(gen[5406]),
			.SE(gen[5407]),

			.SELF(gen[5311]),
			.cell_state(gen[5311])
		); 

/******************* CELL 5312 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5312 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5216]),
			.N(gen[5217]),
			.NE(gen[5218]),

			.O(gen[5311]),
			.E(gen[5313]),

			.SO(gen[5406]),
			.S(gen[5407]),
			.SE(gen[5408]),

			.SELF(gen[5312]),
			.cell_state(gen[5312])
		); 

/******************* CELL 5313 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5313 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5217]),
			.N(gen[5218]),
			.NE(gen[5219]),

			.O(gen[5312]),
			.E(gen[5314]),

			.SO(gen[5407]),
			.S(gen[5408]),
			.SE(gen[5409]),

			.SELF(gen[5313]),
			.cell_state(gen[5313])
		); 

/******************* CELL 5314 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5314 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5218]),
			.N(gen[5219]),
			.NE(gen[5220]),

			.O(gen[5313]),
			.E(gen[5315]),

			.SO(gen[5408]),
			.S(gen[5409]),
			.SE(gen[5410]),

			.SELF(gen[5314]),
			.cell_state(gen[5314])
		); 

/******************* CELL 5315 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5315 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5219]),
			.N(gen[5220]),
			.NE(gen[5221]),

			.O(gen[5314]),
			.E(gen[5316]),

			.SO(gen[5409]),
			.S(gen[5410]),
			.SE(gen[5411]),

			.SELF(gen[5315]),
			.cell_state(gen[5315])
		); 

/******************* CELL 5316 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5316 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5220]),
			.N(gen[5221]),
			.NE(gen[5222]),

			.O(gen[5315]),
			.E(gen[5317]),

			.SO(gen[5410]),
			.S(gen[5411]),
			.SE(gen[5412]),

			.SELF(gen[5316]),
			.cell_state(gen[5316])
		); 

/******************* CELL 5317 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5317 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5221]),
			.N(gen[5222]),
			.NE(gen[5223]),

			.O(gen[5316]),
			.E(gen[5318]),

			.SO(gen[5411]),
			.S(gen[5412]),
			.SE(gen[5413]),

			.SELF(gen[5317]),
			.cell_state(gen[5317])
		); 

/******************* CELL 5318 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5318 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5222]),
			.N(gen[5223]),
			.NE(gen[5224]),

			.O(gen[5317]),
			.E(gen[5319]),

			.SO(gen[5412]),
			.S(gen[5413]),
			.SE(gen[5414]),

			.SELF(gen[5318]),
			.cell_state(gen[5318])
		); 

/******************* CELL 5319 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5319 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5223]),
			.N(gen[5224]),
			.NE(gen[5223]),

			.O(gen[5318]),
			.E(gen[5318]),

			.SO(gen[5413]),
			.S(gen[5414]),
			.SE(gen[5413]),

			.SELF(gen[5319]),
			.cell_state(gen[5319])
		); 

/******************* CELL 5320 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5320 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5226]),
			.N(gen[5225]),
			.NE(gen[5226]),

			.O(gen[5321]),
			.E(gen[5321]),

			.SO(gen[5416]),
			.S(gen[5415]),
			.SE(gen[5416]),

			.SELF(gen[5320]),
			.cell_state(gen[5320])
		); 

/******************* CELL 5321 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5321 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5225]),
			.N(gen[5226]),
			.NE(gen[5227]),

			.O(gen[5320]),
			.E(gen[5322]),

			.SO(gen[5415]),
			.S(gen[5416]),
			.SE(gen[5417]),

			.SELF(gen[5321]),
			.cell_state(gen[5321])
		); 

/******************* CELL 5322 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5322 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5226]),
			.N(gen[5227]),
			.NE(gen[5228]),

			.O(gen[5321]),
			.E(gen[5323]),

			.SO(gen[5416]),
			.S(gen[5417]),
			.SE(gen[5418]),

			.SELF(gen[5322]),
			.cell_state(gen[5322])
		); 

/******************* CELL 5323 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5323 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5227]),
			.N(gen[5228]),
			.NE(gen[5229]),

			.O(gen[5322]),
			.E(gen[5324]),

			.SO(gen[5417]),
			.S(gen[5418]),
			.SE(gen[5419]),

			.SELF(gen[5323]),
			.cell_state(gen[5323])
		); 

/******************* CELL 5324 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5324 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5228]),
			.N(gen[5229]),
			.NE(gen[5230]),

			.O(gen[5323]),
			.E(gen[5325]),

			.SO(gen[5418]),
			.S(gen[5419]),
			.SE(gen[5420]),

			.SELF(gen[5324]),
			.cell_state(gen[5324])
		); 

/******************* CELL 5325 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5325 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5229]),
			.N(gen[5230]),
			.NE(gen[5231]),

			.O(gen[5324]),
			.E(gen[5326]),

			.SO(gen[5419]),
			.S(gen[5420]),
			.SE(gen[5421]),

			.SELF(gen[5325]),
			.cell_state(gen[5325])
		); 

/******************* CELL 5326 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5326 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5230]),
			.N(gen[5231]),
			.NE(gen[5232]),

			.O(gen[5325]),
			.E(gen[5327]),

			.SO(gen[5420]),
			.S(gen[5421]),
			.SE(gen[5422]),

			.SELF(gen[5326]),
			.cell_state(gen[5326])
		); 

/******************* CELL 5327 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5327 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5231]),
			.N(gen[5232]),
			.NE(gen[5233]),

			.O(gen[5326]),
			.E(gen[5328]),

			.SO(gen[5421]),
			.S(gen[5422]),
			.SE(gen[5423]),

			.SELF(gen[5327]),
			.cell_state(gen[5327])
		); 

/******************* CELL 5328 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5328 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5232]),
			.N(gen[5233]),
			.NE(gen[5234]),

			.O(gen[5327]),
			.E(gen[5329]),

			.SO(gen[5422]),
			.S(gen[5423]),
			.SE(gen[5424]),

			.SELF(gen[5328]),
			.cell_state(gen[5328])
		); 

/******************* CELL 5329 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5329 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5233]),
			.N(gen[5234]),
			.NE(gen[5235]),

			.O(gen[5328]),
			.E(gen[5330]),

			.SO(gen[5423]),
			.S(gen[5424]),
			.SE(gen[5425]),

			.SELF(gen[5329]),
			.cell_state(gen[5329])
		); 

/******************* CELL 5330 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5330 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5234]),
			.N(gen[5235]),
			.NE(gen[5236]),

			.O(gen[5329]),
			.E(gen[5331]),

			.SO(gen[5424]),
			.S(gen[5425]),
			.SE(gen[5426]),

			.SELF(gen[5330]),
			.cell_state(gen[5330])
		); 

/******************* CELL 5331 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5331 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5235]),
			.N(gen[5236]),
			.NE(gen[5237]),

			.O(gen[5330]),
			.E(gen[5332]),

			.SO(gen[5425]),
			.S(gen[5426]),
			.SE(gen[5427]),

			.SELF(gen[5331]),
			.cell_state(gen[5331])
		); 

/******************* CELL 5332 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5332 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5236]),
			.N(gen[5237]),
			.NE(gen[5238]),

			.O(gen[5331]),
			.E(gen[5333]),

			.SO(gen[5426]),
			.S(gen[5427]),
			.SE(gen[5428]),

			.SELF(gen[5332]),
			.cell_state(gen[5332])
		); 

/******************* CELL 5333 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5333 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5237]),
			.N(gen[5238]),
			.NE(gen[5239]),

			.O(gen[5332]),
			.E(gen[5334]),

			.SO(gen[5427]),
			.S(gen[5428]),
			.SE(gen[5429]),

			.SELF(gen[5333]),
			.cell_state(gen[5333])
		); 

/******************* CELL 5334 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5334 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5238]),
			.N(gen[5239]),
			.NE(gen[5240]),

			.O(gen[5333]),
			.E(gen[5335]),

			.SO(gen[5428]),
			.S(gen[5429]),
			.SE(gen[5430]),

			.SELF(gen[5334]),
			.cell_state(gen[5334])
		); 

/******************* CELL 5335 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5335 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5239]),
			.N(gen[5240]),
			.NE(gen[5241]),

			.O(gen[5334]),
			.E(gen[5336]),

			.SO(gen[5429]),
			.S(gen[5430]),
			.SE(gen[5431]),

			.SELF(gen[5335]),
			.cell_state(gen[5335])
		); 

/******************* CELL 5336 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5336 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5240]),
			.N(gen[5241]),
			.NE(gen[5242]),

			.O(gen[5335]),
			.E(gen[5337]),

			.SO(gen[5430]),
			.S(gen[5431]),
			.SE(gen[5432]),

			.SELF(gen[5336]),
			.cell_state(gen[5336])
		); 

/******************* CELL 5337 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5337 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5241]),
			.N(gen[5242]),
			.NE(gen[5243]),

			.O(gen[5336]),
			.E(gen[5338]),

			.SO(gen[5431]),
			.S(gen[5432]),
			.SE(gen[5433]),

			.SELF(gen[5337]),
			.cell_state(gen[5337])
		); 

/******************* CELL 5338 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5338 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5242]),
			.N(gen[5243]),
			.NE(gen[5244]),

			.O(gen[5337]),
			.E(gen[5339]),

			.SO(gen[5432]),
			.S(gen[5433]),
			.SE(gen[5434]),

			.SELF(gen[5338]),
			.cell_state(gen[5338])
		); 

/******************* CELL 5339 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5339 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5243]),
			.N(gen[5244]),
			.NE(gen[5245]),

			.O(gen[5338]),
			.E(gen[5340]),

			.SO(gen[5433]),
			.S(gen[5434]),
			.SE(gen[5435]),

			.SELF(gen[5339]),
			.cell_state(gen[5339])
		); 

/******************* CELL 5340 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5340 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5244]),
			.N(gen[5245]),
			.NE(gen[5246]),

			.O(gen[5339]),
			.E(gen[5341]),

			.SO(gen[5434]),
			.S(gen[5435]),
			.SE(gen[5436]),

			.SELF(gen[5340]),
			.cell_state(gen[5340])
		); 

/******************* CELL 5341 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5341 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5245]),
			.N(gen[5246]),
			.NE(gen[5247]),

			.O(gen[5340]),
			.E(gen[5342]),

			.SO(gen[5435]),
			.S(gen[5436]),
			.SE(gen[5437]),

			.SELF(gen[5341]),
			.cell_state(gen[5341])
		); 

/******************* CELL 5342 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5342 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5246]),
			.N(gen[5247]),
			.NE(gen[5248]),

			.O(gen[5341]),
			.E(gen[5343]),

			.SO(gen[5436]),
			.S(gen[5437]),
			.SE(gen[5438]),

			.SELF(gen[5342]),
			.cell_state(gen[5342])
		); 

/******************* CELL 5343 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5343 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5247]),
			.N(gen[5248]),
			.NE(gen[5249]),

			.O(gen[5342]),
			.E(gen[5344]),

			.SO(gen[5437]),
			.S(gen[5438]),
			.SE(gen[5439]),

			.SELF(gen[5343]),
			.cell_state(gen[5343])
		); 

/******************* CELL 5344 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5344 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5248]),
			.N(gen[5249]),
			.NE(gen[5250]),

			.O(gen[5343]),
			.E(gen[5345]),

			.SO(gen[5438]),
			.S(gen[5439]),
			.SE(gen[5440]),

			.SELF(gen[5344]),
			.cell_state(gen[5344])
		); 

/******************* CELL 5345 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5345 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5249]),
			.N(gen[5250]),
			.NE(gen[5251]),

			.O(gen[5344]),
			.E(gen[5346]),

			.SO(gen[5439]),
			.S(gen[5440]),
			.SE(gen[5441]),

			.SELF(gen[5345]),
			.cell_state(gen[5345])
		); 

/******************* CELL 5346 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5346 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5250]),
			.N(gen[5251]),
			.NE(gen[5252]),

			.O(gen[5345]),
			.E(gen[5347]),

			.SO(gen[5440]),
			.S(gen[5441]),
			.SE(gen[5442]),

			.SELF(gen[5346]),
			.cell_state(gen[5346])
		); 

/******************* CELL 5347 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5347 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5251]),
			.N(gen[5252]),
			.NE(gen[5253]),

			.O(gen[5346]),
			.E(gen[5348]),

			.SO(gen[5441]),
			.S(gen[5442]),
			.SE(gen[5443]),

			.SELF(gen[5347]),
			.cell_state(gen[5347])
		); 

/******************* CELL 5348 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5348 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5252]),
			.N(gen[5253]),
			.NE(gen[5254]),

			.O(gen[5347]),
			.E(gen[5349]),

			.SO(gen[5442]),
			.S(gen[5443]),
			.SE(gen[5444]),

			.SELF(gen[5348]),
			.cell_state(gen[5348])
		); 

/******************* CELL 5349 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5349 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5253]),
			.N(gen[5254]),
			.NE(gen[5255]),

			.O(gen[5348]),
			.E(gen[5350]),

			.SO(gen[5443]),
			.S(gen[5444]),
			.SE(gen[5445]),

			.SELF(gen[5349]),
			.cell_state(gen[5349])
		); 

/******************* CELL 5350 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5350 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5254]),
			.N(gen[5255]),
			.NE(gen[5256]),

			.O(gen[5349]),
			.E(gen[5351]),

			.SO(gen[5444]),
			.S(gen[5445]),
			.SE(gen[5446]),

			.SELF(gen[5350]),
			.cell_state(gen[5350])
		); 

/******************* CELL 5351 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5351 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5255]),
			.N(gen[5256]),
			.NE(gen[5257]),

			.O(gen[5350]),
			.E(gen[5352]),

			.SO(gen[5445]),
			.S(gen[5446]),
			.SE(gen[5447]),

			.SELF(gen[5351]),
			.cell_state(gen[5351])
		); 

/******************* CELL 5352 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5352 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5256]),
			.N(gen[5257]),
			.NE(gen[5258]),

			.O(gen[5351]),
			.E(gen[5353]),

			.SO(gen[5446]),
			.S(gen[5447]),
			.SE(gen[5448]),

			.SELF(gen[5352]),
			.cell_state(gen[5352])
		); 

/******************* CELL 5353 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5353 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5257]),
			.N(gen[5258]),
			.NE(gen[5259]),

			.O(gen[5352]),
			.E(gen[5354]),

			.SO(gen[5447]),
			.S(gen[5448]),
			.SE(gen[5449]),

			.SELF(gen[5353]),
			.cell_state(gen[5353])
		); 

/******************* CELL 5354 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5354 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5258]),
			.N(gen[5259]),
			.NE(gen[5260]),

			.O(gen[5353]),
			.E(gen[5355]),

			.SO(gen[5448]),
			.S(gen[5449]),
			.SE(gen[5450]),

			.SELF(gen[5354]),
			.cell_state(gen[5354])
		); 

/******************* CELL 5355 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5355 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5259]),
			.N(gen[5260]),
			.NE(gen[5261]),

			.O(gen[5354]),
			.E(gen[5356]),

			.SO(gen[5449]),
			.S(gen[5450]),
			.SE(gen[5451]),

			.SELF(gen[5355]),
			.cell_state(gen[5355])
		); 

/******************* CELL 5356 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5356 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5260]),
			.N(gen[5261]),
			.NE(gen[5262]),

			.O(gen[5355]),
			.E(gen[5357]),

			.SO(gen[5450]),
			.S(gen[5451]),
			.SE(gen[5452]),

			.SELF(gen[5356]),
			.cell_state(gen[5356])
		); 

/******************* CELL 5357 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5357 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5261]),
			.N(gen[5262]),
			.NE(gen[5263]),

			.O(gen[5356]),
			.E(gen[5358]),

			.SO(gen[5451]),
			.S(gen[5452]),
			.SE(gen[5453]),

			.SELF(gen[5357]),
			.cell_state(gen[5357])
		); 

/******************* CELL 5358 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5358 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5262]),
			.N(gen[5263]),
			.NE(gen[5264]),

			.O(gen[5357]),
			.E(gen[5359]),

			.SO(gen[5452]),
			.S(gen[5453]),
			.SE(gen[5454]),

			.SELF(gen[5358]),
			.cell_state(gen[5358])
		); 

/******************* CELL 5359 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5359 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5263]),
			.N(gen[5264]),
			.NE(gen[5265]),

			.O(gen[5358]),
			.E(gen[5360]),

			.SO(gen[5453]),
			.S(gen[5454]),
			.SE(gen[5455]),

			.SELF(gen[5359]),
			.cell_state(gen[5359])
		); 

/******************* CELL 5360 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5360 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5264]),
			.N(gen[5265]),
			.NE(gen[5266]),

			.O(gen[5359]),
			.E(gen[5361]),

			.SO(gen[5454]),
			.S(gen[5455]),
			.SE(gen[5456]),

			.SELF(gen[5360]),
			.cell_state(gen[5360])
		); 

/******************* CELL 5361 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5361 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5265]),
			.N(gen[5266]),
			.NE(gen[5267]),

			.O(gen[5360]),
			.E(gen[5362]),

			.SO(gen[5455]),
			.S(gen[5456]),
			.SE(gen[5457]),

			.SELF(gen[5361]),
			.cell_state(gen[5361])
		); 

/******************* CELL 5362 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5362 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5266]),
			.N(gen[5267]),
			.NE(gen[5268]),

			.O(gen[5361]),
			.E(gen[5363]),

			.SO(gen[5456]),
			.S(gen[5457]),
			.SE(gen[5458]),

			.SELF(gen[5362]),
			.cell_state(gen[5362])
		); 

/******************* CELL 5363 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5363 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5267]),
			.N(gen[5268]),
			.NE(gen[5269]),

			.O(gen[5362]),
			.E(gen[5364]),

			.SO(gen[5457]),
			.S(gen[5458]),
			.SE(gen[5459]),

			.SELF(gen[5363]),
			.cell_state(gen[5363])
		); 

/******************* CELL 5364 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5364 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5268]),
			.N(gen[5269]),
			.NE(gen[5270]),

			.O(gen[5363]),
			.E(gen[5365]),

			.SO(gen[5458]),
			.S(gen[5459]),
			.SE(gen[5460]),

			.SELF(gen[5364]),
			.cell_state(gen[5364])
		); 

/******************* CELL 5365 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5365 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5269]),
			.N(gen[5270]),
			.NE(gen[5271]),

			.O(gen[5364]),
			.E(gen[5366]),

			.SO(gen[5459]),
			.S(gen[5460]),
			.SE(gen[5461]),

			.SELF(gen[5365]),
			.cell_state(gen[5365])
		); 

/******************* CELL 5366 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5366 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5270]),
			.N(gen[5271]),
			.NE(gen[5272]),

			.O(gen[5365]),
			.E(gen[5367]),

			.SO(gen[5460]),
			.S(gen[5461]),
			.SE(gen[5462]),

			.SELF(gen[5366]),
			.cell_state(gen[5366])
		); 

/******************* CELL 5367 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5367 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5271]),
			.N(gen[5272]),
			.NE(gen[5273]),

			.O(gen[5366]),
			.E(gen[5368]),

			.SO(gen[5461]),
			.S(gen[5462]),
			.SE(gen[5463]),

			.SELF(gen[5367]),
			.cell_state(gen[5367])
		); 

/******************* CELL 5368 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5368 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5272]),
			.N(gen[5273]),
			.NE(gen[5274]),

			.O(gen[5367]),
			.E(gen[5369]),

			.SO(gen[5462]),
			.S(gen[5463]),
			.SE(gen[5464]),

			.SELF(gen[5368]),
			.cell_state(gen[5368])
		); 

/******************* CELL 5369 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5369 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5273]),
			.N(gen[5274]),
			.NE(gen[5275]),

			.O(gen[5368]),
			.E(gen[5370]),

			.SO(gen[5463]),
			.S(gen[5464]),
			.SE(gen[5465]),

			.SELF(gen[5369]),
			.cell_state(gen[5369])
		); 

/******************* CELL 5370 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5370 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5274]),
			.N(gen[5275]),
			.NE(gen[5276]),

			.O(gen[5369]),
			.E(gen[5371]),

			.SO(gen[5464]),
			.S(gen[5465]),
			.SE(gen[5466]),

			.SELF(gen[5370]),
			.cell_state(gen[5370])
		); 

/******************* CELL 5371 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5371 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5275]),
			.N(gen[5276]),
			.NE(gen[5277]),

			.O(gen[5370]),
			.E(gen[5372]),

			.SO(gen[5465]),
			.S(gen[5466]),
			.SE(gen[5467]),

			.SELF(gen[5371]),
			.cell_state(gen[5371])
		); 

/******************* CELL 5372 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5372 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5276]),
			.N(gen[5277]),
			.NE(gen[5278]),

			.O(gen[5371]),
			.E(gen[5373]),

			.SO(gen[5466]),
			.S(gen[5467]),
			.SE(gen[5468]),

			.SELF(gen[5372]),
			.cell_state(gen[5372])
		); 

/******************* CELL 5373 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5373 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5277]),
			.N(gen[5278]),
			.NE(gen[5279]),

			.O(gen[5372]),
			.E(gen[5374]),

			.SO(gen[5467]),
			.S(gen[5468]),
			.SE(gen[5469]),

			.SELF(gen[5373]),
			.cell_state(gen[5373])
		); 

/******************* CELL 5374 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5374 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5278]),
			.N(gen[5279]),
			.NE(gen[5280]),

			.O(gen[5373]),
			.E(gen[5375]),

			.SO(gen[5468]),
			.S(gen[5469]),
			.SE(gen[5470]),

			.SELF(gen[5374]),
			.cell_state(gen[5374])
		); 

/******************* CELL 5375 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5375 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5279]),
			.N(gen[5280]),
			.NE(gen[5281]),

			.O(gen[5374]),
			.E(gen[5376]),

			.SO(gen[5469]),
			.S(gen[5470]),
			.SE(gen[5471]),

			.SELF(gen[5375]),
			.cell_state(gen[5375])
		); 

/******************* CELL 5376 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5376 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5280]),
			.N(gen[5281]),
			.NE(gen[5282]),

			.O(gen[5375]),
			.E(gen[5377]),

			.SO(gen[5470]),
			.S(gen[5471]),
			.SE(gen[5472]),

			.SELF(gen[5376]),
			.cell_state(gen[5376])
		); 

/******************* CELL 5377 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5377 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5281]),
			.N(gen[5282]),
			.NE(gen[5283]),

			.O(gen[5376]),
			.E(gen[5378]),

			.SO(gen[5471]),
			.S(gen[5472]),
			.SE(gen[5473]),

			.SELF(gen[5377]),
			.cell_state(gen[5377])
		); 

/******************* CELL 5378 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5378 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5282]),
			.N(gen[5283]),
			.NE(gen[5284]),

			.O(gen[5377]),
			.E(gen[5379]),

			.SO(gen[5472]),
			.S(gen[5473]),
			.SE(gen[5474]),

			.SELF(gen[5378]),
			.cell_state(gen[5378])
		); 

/******************* CELL 5379 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5379 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5283]),
			.N(gen[5284]),
			.NE(gen[5285]),

			.O(gen[5378]),
			.E(gen[5380]),

			.SO(gen[5473]),
			.S(gen[5474]),
			.SE(gen[5475]),

			.SELF(gen[5379]),
			.cell_state(gen[5379])
		); 

/******************* CELL 5380 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5380 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5284]),
			.N(gen[5285]),
			.NE(gen[5286]),

			.O(gen[5379]),
			.E(gen[5381]),

			.SO(gen[5474]),
			.S(gen[5475]),
			.SE(gen[5476]),

			.SELF(gen[5380]),
			.cell_state(gen[5380])
		); 

/******************* CELL 5381 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5381 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5285]),
			.N(gen[5286]),
			.NE(gen[5287]),

			.O(gen[5380]),
			.E(gen[5382]),

			.SO(gen[5475]),
			.S(gen[5476]),
			.SE(gen[5477]),

			.SELF(gen[5381]),
			.cell_state(gen[5381])
		); 

/******************* CELL 5382 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5382 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5286]),
			.N(gen[5287]),
			.NE(gen[5288]),

			.O(gen[5381]),
			.E(gen[5383]),

			.SO(gen[5476]),
			.S(gen[5477]),
			.SE(gen[5478]),

			.SELF(gen[5382]),
			.cell_state(gen[5382])
		); 

/******************* CELL 5383 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5383 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5287]),
			.N(gen[5288]),
			.NE(gen[5289]),

			.O(gen[5382]),
			.E(gen[5384]),

			.SO(gen[5477]),
			.S(gen[5478]),
			.SE(gen[5479]),

			.SELF(gen[5383]),
			.cell_state(gen[5383])
		); 

/******************* CELL 5384 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5384 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5288]),
			.N(gen[5289]),
			.NE(gen[5290]),

			.O(gen[5383]),
			.E(gen[5385]),

			.SO(gen[5478]),
			.S(gen[5479]),
			.SE(gen[5480]),

			.SELF(gen[5384]),
			.cell_state(gen[5384])
		); 

/******************* CELL 5385 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5385 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5289]),
			.N(gen[5290]),
			.NE(gen[5291]),

			.O(gen[5384]),
			.E(gen[5386]),

			.SO(gen[5479]),
			.S(gen[5480]),
			.SE(gen[5481]),

			.SELF(gen[5385]),
			.cell_state(gen[5385])
		); 

/******************* CELL 5386 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5386 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5290]),
			.N(gen[5291]),
			.NE(gen[5292]),

			.O(gen[5385]),
			.E(gen[5387]),

			.SO(gen[5480]),
			.S(gen[5481]),
			.SE(gen[5482]),

			.SELF(gen[5386]),
			.cell_state(gen[5386])
		); 

/******************* CELL 5387 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5387 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5291]),
			.N(gen[5292]),
			.NE(gen[5293]),

			.O(gen[5386]),
			.E(gen[5388]),

			.SO(gen[5481]),
			.S(gen[5482]),
			.SE(gen[5483]),

			.SELF(gen[5387]),
			.cell_state(gen[5387])
		); 

/******************* CELL 5388 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5388 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5292]),
			.N(gen[5293]),
			.NE(gen[5294]),

			.O(gen[5387]),
			.E(gen[5389]),

			.SO(gen[5482]),
			.S(gen[5483]),
			.SE(gen[5484]),

			.SELF(gen[5388]),
			.cell_state(gen[5388])
		); 

/******************* CELL 5389 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5389 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5293]),
			.N(gen[5294]),
			.NE(gen[5295]),

			.O(gen[5388]),
			.E(gen[5390]),

			.SO(gen[5483]),
			.S(gen[5484]),
			.SE(gen[5485]),

			.SELF(gen[5389]),
			.cell_state(gen[5389])
		); 

/******************* CELL 5390 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5390 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5294]),
			.N(gen[5295]),
			.NE(gen[5296]),

			.O(gen[5389]),
			.E(gen[5391]),

			.SO(gen[5484]),
			.S(gen[5485]),
			.SE(gen[5486]),

			.SELF(gen[5390]),
			.cell_state(gen[5390])
		); 

/******************* CELL 5391 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5391 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5295]),
			.N(gen[5296]),
			.NE(gen[5297]),

			.O(gen[5390]),
			.E(gen[5392]),

			.SO(gen[5485]),
			.S(gen[5486]),
			.SE(gen[5487]),

			.SELF(gen[5391]),
			.cell_state(gen[5391])
		); 

/******************* CELL 5392 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5392 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5296]),
			.N(gen[5297]),
			.NE(gen[5298]),

			.O(gen[5391]),
			.E(gen[5393]),

			.SO(gen[5486]),
			.S(gen[5487]),
			.SE(gen[5488]),

			.SELF(gen[5392]),
			.cell_state(gen[5392])
		); 

/******************* CELL 5393 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5393 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5297]),
			.N(gen[5298]),
			.NE(gen[5299]),

			.O(gen[5392]),
			.E(gen[5394]),

			.SO(gen[5487]),
			.S(gen[5488]),
			.SE(gen[5489]),

			.SELF(gen[5393]),
			.cell_state(gen[5393])
		); 

/******************* CELL 5394 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5394 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5298]),
			.N(gen[5299]),
			.NE(gen[5300]),

			.O(gen[5393]),
			.E(gen[5395]),

			.SO(gen[5488]),
			.S(gen[5489]),
			.SE(gen[5490]),

			.SELF(gen[5394]),
			.cell_state(gen[5394])
		); 

/******************* CELL 5395 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5395 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5299]),
			.N(gen[5300]),
			.NE(gen[5301]),

			.O(gen[5394]),
			.E(gen[5396]),

			.SO(gen[5489]),
			.S(gen[5490]),
			.SE(gen[5491]),

			.SELF(gen[5395]),
			.cell_state(gen[5395])
		); 

/******************* CELL 5396 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5396 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5300]),
			.N(gen[5301]),
			.NE(gen[5302]),

			.O(gen[5395]),
			.E(gen[5397]),

			.SO(gen[5490]),
			.S(gen[5491]),
			.SE(gen[5492]),

			.SELF(gen[5396]),
			.cell_state(gen[5396])
		); 

/******************* CELL 5397 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5397 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5301]),
			.N(gen[5302]),
			.NE(gen[5303]),

			.O(gen[5396]),
			.E(gen[5398]),

			.SO(gen[5491]),
			.S(gen[5492]),
			.SE(gen[5493]),

			.SELF(gen[5397]),
			.cell_state(gen[5397])
		); 

/******************* CELL 5398 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5398 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5302]),
			.N(gen[5303]),
			.NE(gen[5304]),

			.O(gen[5397]),
			.E(gen[5399]),

			.SO(gen[5492]),
			.S(gen[5493]),
			.SE(gen[5494]),

			.SELF(gen[5398]),
			.cell_state(gen[5398])
		); 

/******************* CELL 5399 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5399 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5303]),
			.N(gen[5304]),
			.NE(gen[5305]),

			.O(gen[5398]),
			.E(gen[5400]),

			.SO(gen[5493]),
			.S(gen[5494]),
			.SE(gen[5495]),

			.SELF(gen[5399]),
			.cell_state(gen[5399])
		); 

/******************* CELL 5400 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5400 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5304]),
			.N(gen[5305]),
			.NE(gen[5306]),

			.O(gen[5399]),
			.E(gen[5401]),

			.SO(gen[5494]),
			.S(gen[5495]),
			.SE(gen[5496]),

			.SELF(gen[5400]),
			.cell_state(gen[5400])
		); 

/******************* CELL 5401 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5401 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5305]),
			.N(gen[5306]),
			.NE(gen[5307]),

			.O(gen[5400]),
			.E(gen[5402]),

			.SO(gen[5495]),
			.S(gen[5496]),
			.SE(gen[5497]),

			.SELF(gen[5401]),
			.cell_state(gen[5401])
		); 

/******************* CELL 5402 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5402 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5306]),
			.N(gen[5307]),
			.NE(gen[5308]),

			.O(gen[5401]),
			.E(gen[5403]),

			.SO(gen[5496]),
			.S(gen[5497]),
			.SE(gen[5498]),

			.SELF(gen[5402]),
			.cell_state(gen[5402])
		); 

/******************* CELL 5403 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5403 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5307]),
			.N(gen[5308]),
			.NE(gen[5309]),

			.O(gen[5402]),
			.E(gen[5404]),

			.SO(gen[5497]),
			.S(gen[5498]),
			.SE(gen[5499]),

			.SELF(gen[5403]),
			.cell_state(gen[5403])
		); 

/******************* CELL 5404 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5404 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5308]),
			.N(gen[5309]),
			.NE(gen[5310]),

			.O(gen[5403]),
			.E(gen[5405]),

			.SO(gen[5498]),
			.S(gen[5499]),
			.SE(gen[5500]),

			.SELF(gen[5404]),
			.cell_state(gen[5404])
		); 

/******************* CELL 5405 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5405 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5309]),
			.N(gen[5310]),
			.NE(gen[5311]),

			.O(gen[5404]),
			.E(gen[5406]),

			.SO(gen[5499]),
			.S(gen[5500]),
			.SE(gen[5501]),

			.SELF(gen[5405]),
			.cell_state(gen[5405])
		); 

/******************* CELL 5406 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5406 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5310]),
			.N(gen[5311]),
			.NE(gen[5312]),

			.O(gen[5405]),
			.E(gen[5407]),

			.SO(gen[5500]),
			.S(gen[5501]),
			.SE(gen[5502]),

			.SELF(gen[5406]),
			.cell_state(gen[5406])
		); 

/******************* CELL 5407 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5407 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5311]),
			.N(gen[5312]),
			.NE(gen[5313]),

			.O(gen[5406]),
			.E(gen[5408]),

			.SO(gen[5501]),
			.S(gen[5502]),
			.SE(gen[5503]),

			.SELF(gen[5407]),
			.cell_state(gen[5407])
		); 

/******************* CELL 5408 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5408 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5312]),
			.N(gen[5313]),
			.NE(gen[5314]),

			.O(gen[5407]),
			.E(gen[5409]),

			.SO(gen[5502]),
			.S(gen[5503]),
			.SE(gen[5504]),

			.SELF(gen[5408]),
			.cell_state(gen[5408])
		); 

/******************* CELL 5409 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5409 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5313]),
			.N(gen[5314]),
			.NE(gen[5315]),

			.O(gen[5408]),
			.E(gen[5410]),

			.SO(gen[5503]),
			.S(gen[5504]),
			.SE(gen[5505]),

			.SELF(gen[5409]),
			.cell_state(gen[5409])
		); 

/******************* CELL 5410 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5410 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5314]),
			.N(gen[5315]),
			.NE(gen[5316]),

			.O(gen[5409]),
			.E(gen[5411]),

			.SO(gen[5504]),
			.S(gen[5505]),
			.SE(gen[5506]),

			.SELF(gen[5410]),
			.cell_state(gen[5410])
		); 

/******************* CELL 5411 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5411 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5315]),
			.N(gen[5316]),
			.NE(gen[5317]),

			.O(gen[5410]),
			.E(gen[5412]),

			.SO(gen[5505]),
			.S(gen[5506]),
			.SE(gen[5507]),

			.SELF(gen[5411]),
			.cell_state(gen[5411])
		); 

/******************* CELL 5412 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5412 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5316]),
			.N(gen[5317]),
			.NE(gen[5318]),

			.O(gen[5411]),
			.E(gen[5413]),

			.SO(gen[5506]),
			.S(gen[5507]),
			.SE(gen[5508]),

			.SELF(gen[5412]),
			.cell_state(gen[5412])
		); 

/******************* CELL 5413 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5413 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5317]),
			.N(gen[5318]),
			.NE(gen[5319]),

			.O(gen[5412]),
			.E(gen[5414]),

			.SO(gen[5507]),
			.S(gen[5508]),
			.SE(gen[5509]),

			.SELF(gen[5413]),
			.cell_state(gen[5413])
		); 

/******************* CELL 5414 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5414 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5318]),
			.N(gen[5319]),
			.NE(gen[5318]),

			.O(gen[5413]),
			.E(gen[5413]),

			.SO(gen[5508]),
			.S(gen[5509]),
			.SE(gen[5508]),

			.SELF(gen[5414]),
			.cell_state(gen[5414])
		); 

/******************* CELL 5415 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5415 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5321]),
			.N(gen[5320]),
			.NE(gen[5321]),

			.O(gen[5416]),
			.E(gen[5416]),

			.SO(gen[5511]),
			.S(gen[5510]),
			.SE(gen[5511]),

			.SELF(gen[5415]),
			.cell_state(gen[5415])
		); 

/******************* CELL 5416 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5416 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5320]),
			.N(gen[5321]),
			.NE(gen[5322]),

			.O(gen[5415]),
			.E(gen[5417]),

			.SO(gen[5510]),
			.S(gen[5511]),
			.SE(gen[5512]),

			.SELF(gen[5416]),
			.cell_state(gen[5416])
		); 

/******************* CELL 5417 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5417 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5321]),
			.N(gen[5322]),
			.NE(gen[5323]),

			.O(gen[5416]),
			.E(gen[5418]),

			.SO(gen[5511]),
			.S(gen[5512]),
			.SE(gen[5513]),

			.SELF(gen[5417]),
			.cell_state(gen[5417])
		); 

/******************* CELL 5418 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5418 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5322]),
			.N(gen[5323]),
			.NE(gen[5324]),

			.O(gen[5417]),
			.E(gen[5419]),

			.SO(gen[5512]),
			.S(gen[5513]),
			.SE(gen[5514]),

			.SELF(gen[5418]),
			.cell_state(gen[5418])
		); 

/******************* CELL 5419 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5419 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5323]),
			.N(gen[5324]),
			.NE(gen[5325]),

			.O(gen[5418]),
			.E(gen[5420]),

			.SO(gen[5513]),
			.S(gen[5514]),
			.SE(gen[5515]),

			.SELF(gen[5419]),
			.cell_state(gen[5419])
		); 

/******************* CELL 5420 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5420 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5324]),
			.N(gen[5325]),
			.NE(gen[5326]),

			.O(gen[5419]),
			.E(gen[5421]),

			.SO(gen[5514]),
			.S(gen[5515]),
			.SE(gen[5516]),

			.SELF(gen[5420]),
			.cell_state(gen[5420])
		); 

/******************* CELL 5421 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5421 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5325]),
			.N(gen[5326]),
			.NE(gen[5327]),

			.O(gen[5420]),
			.E(gen[5422]),

			.SO(gen[5515]),
			.S(gen[5516]),
			.SE(gen[5517]),

			.SELF(gen[5421]),
			.cell_state(gen[5421])
		); 

/******************* CELL 5422 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5422 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5326]),
			.N(gen[5327]),
			.NE(gen[5328]),

			.O(gen[5421]),
			.E(gen[5423]),

			.SO(gen[5516]),
			.S(gen[5517]),
			.SE(gen[5518]),

			.SELF(gen[5422]),
			.cell_state(gen[5422])
		); 

/******************* CELL 5423 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5423 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5327]),
			.N(gen[5328]),
			.NE(gen[5329]),

			.O(gen[5422]),
			.E(gen[5424]),

			.SO(gen[5517]),
			.S(gen[5518]),
			.SE(gen[5519]),

			.SELF(gen[5423]),
			.cell_state(gen[5423])
		); 

/******************* CELL 5424 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5424 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5328]),
			.N(gen[5329]),
			.NE(gen[5330]),

			.O(gen[5423]),
			.E(gen[5425]),

			.SO(gen[5518]),
			.S(gen[5519]),
			.SE(gen[5520]),

			.SELF(gen[5424]),
			.cell_state(gen[5424])
		); 

/******************* CELL 5425 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5425 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5329]),
			.N(gen[5330]),
			.NE(gen[5331]),

			.O(gen[5424]),
			.E(gen[5426]),

			.SO(gen[5519]),
			.S(gen[5520]),
			.SE(gen[5521]),

			.SELF(gen[5425]),
			.cell_state(gen[5425])
		); 

/******************* CELL 5426 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5426 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5330]),
			.N(gen[5331]),
			.NE(gen[5332]),

			.O(gen[5425]),
			.E(gen[5427]),

			.SO(gen[5520]),
			.S(gen[5521]),
			.SE(gen[5522]),

			.SELF(gen[5426]),
			.cell_state(gen[5426])
		); 

/******************* CELL 5427 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5427 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5331]),
			.N(gen[5332]),
			.NE(gen[5333]),

			.O(gen[5426]),
			.E(gen[5428]),

			.SO(gen[5521]),
			.S(gen[5522]),
			.SE(gen[5523]),

			.SELF(gen[5427]),
			.cell_state(gen[5427])
		); 

/******************* CELL 5428 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5428 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5332]),
			.N(gen[5333]),
			.NE(gen[5334]),

			.O(gen[5427]),
			.E(gen[5429]),

			.SO(gen[5522]),
			.S(gen[5523]),
			.SE(gen[5524]),

			.SELF(gen[5428]),
			.cell_state(gen[5428])
		); 

/******************* CELL 5429 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5429 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5333]),
			.N(gen[5334]),
			.NE(gen[5335]),

			.O(gen[5428]),
			.E(gen[5430]),

			.SO(gen[5523]),
			.S(gen[5524]),
			.SE(gen[5525]),

			.SELF(gen[5429]),
			.cell_state(gen[5429])
		); 

/******************* CELL 5430 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5430 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5334]),
			.N(gen[5335]),
			.NE(gen[5336]),

			.O(gen[5429]),
			.E(gen[5431]),

			.SO(gen[5524]),
			.S(gen[5525]),
			.SE(gen[5526]),

			.SELF(gen[5430]),
			.cell_state(gen[5430])
		); 

/******************* CELL 5431 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5431 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5335]),
			.N(gen[5336]),
			.NE(gen[5337]),

			.O(gen[5430]),
			.E(gen[5432]),

			.SO(gen[5525]),
			.S(gen[5526]),
			.SE(gen[5527]),

			.SELF(gen[5431]),
			.cell_state(gen[5431])
		); 

/******************* CELL 5432 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5432 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5336]),
			.N(gen[5337]),
			.NE(gen[5338]),

			.O(gen[5431]),
			.E(gen[5433]),

			.SO(gen[5526]),
			.S(gen[5527]),
			.SE(gen[5528]),

			.SELF(gen[5432]),
			.cell_state(gen[5432])
		); 

/******************* CELL 5433 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5433 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5337]),
			.N(gen[5338]),
			.NE(gen[5339]),

			.O(gen[5432]),
			.E(gen[5434]),

			.SO(gen[5527]),
			.S(gen[5528]),
			.SE(gen[5529]),

			.SELF(gen[5433]),
			.cell_state(gen[5433])
		); 

/******************* CELL 5434 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5434 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5338]),
			.N(gen[5339]),
			.NE(gen[5340]),

			.O(gen[5433]),
			.E(gen[5435]),

			.SO(gen[5528]),
			.S(gen[5529]),
			.SE(gen[5530]),

			.SELF(gen[5434]),
			.cell_state(gen[5434])
		); 

/******************* CELL 5435 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5435 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5339]),
			.N(gen[5340]),
			.NE(gen[5341]),

			.O(gen[5434]),
			.E(gen[5436]),

			.SO(gen[5529]),
			.S(gen[5530]),
			.SE(gen[5531]),

			.SELF(gen[5435]),
			.cell_state(gen[5435])
		); 

/******************* CELL 5436 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5436 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5340]),
			.N(gen[5341]),
			.NE(gen[5342]),

			.O(gen[5435]),
			.E(gen[5437]),

			.SO(gen[5530]),
			.S(gen[5531]),
			.SE(gen[5532]),

			.SELF(gen[5436]),
			.cell_state(gen[5436])
		); 

/******************* CELL 5437 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5437 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5341]),
			.N(gen[5342]),
			.NE(gen[5343]),

			.O(gen[5436]),
			.E(gen[5438]),

			.SO(gen[5531]),
			.S(gen[5532]),
			.SE(gen[5533]),

			.SELF(gen[5437]),
			.cell_state(gen[5437])
		); 

/******************* CELL 5438 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5438 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5342]),
			.N(gen[5343]),
			.NE(gen[5344]),

			.O(gen[5437]),
			.E(gen[5439]),

			.SO(gen[5532]),
			.S(gen[5533]),
			.SE(gen[5534]),

			.SELF(gen[5438]),
			.cell_state(gen[5438])
		); 

/******************* CELL 5439 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5439 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5343]),
			.N(gen[5344]),
			.NE(gen[5345]),

			.O(gen[5438]),
			.E(gen[5440]),

			.SO(gen[5533]),
			.S(gen[5534]),
			.SE(gen[5535]),

			.SELF(gen[5439]),
			.cell_state(gen[5439])
		); 

/******************* CELL 5440 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5440 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5344]),
			.N(gen[5345]),
			.NE(gen[5346]),

			.O(gen[5439]),
			.E(gen[5441]),

			.SO(gen[5534]),
			.S(gen[5535]),
			.SE(gen[5536]),

			.SELF(gen[5440]),
			.cell_state(gen[5440])
		); 

/******************* CELL 5441 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5441 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5345]),
			.N(gen[5346]),
			.NE(gen[5347]),

			.O(gen[5440]),
			.E(gen[5442]),

			.SO(gen[5535]),
			.S(gen[5536]),
			.SE(gen[5537]),

			.SELF(gen[5441]),
			.cell_state(gen[5441])
		); 

/******************* CELL 5442 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5442 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5346]),
			.N(gen[5347]),
			.NE(gen[5348]),

			.O(gen[5441]),
			.E(gen[5443]),

			.SO(gen[5536]),
			.S(gen[5537]),
			.SE(gen[5538]),

			.SELF(gen[5442]),
			.cell_state(gen[5442])
		); 

/******************* CELL 5443 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5443 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5347]),
			.N(gen[5348]),
			.NE(gen[5349]),

			.O(gen[5442]),
			.E(gen[5444]),

			.SO(gen[5537]),
			.S(gen[5538]),
			.SE(gen[5539]),

			.SELF(gen[5443]),
			.cell_state(gen[5443])
		); 

/******************* CELL 5444 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5444 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5348]),
			.N(gen[5349]),
			.NE(gen[5350]),

			.O(gen[5443]),
			.E(gen[5445]),

			.SO(gen[5538]),
			.S(gen[5539]),
			.SE(gen[5540]),

			.SELF(gen[5444]),
			.cell_state(gen[5444])
		); 

/******************* CELL 5445 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5445 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5349]),
			.N(gen[5350]),
			.NE(gen[5351]),

			.O(gen[5444]),
			.E(gen[5446]),

			.SO(gen[5539]),
			.S(gen[5540]),
			.SE(gen[5541]),

			.SELF(gen[5445]),
			.cell_state(gen[5445])
		); 

/******************* CELL 5446 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5446 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5350]),
			.N(gen[5351]),
			.NE(gen[5352]),

			.O(gen[5445]),
			.E(gen[5447]),

			.SO(gen[5540]),
			.S(gen[5541]),
			.SE(gen[5542]),

			.SELF(gen[5446]),
			.cell_state(gen[5446])
		); 

/******************* CELL 5447 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5447 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5351]),
			.N(gen[5352]),
			.NE(gen[5353]),

			.O(gen[5446]),
			.E(gen[5448]),

			.SO(gen[5541]),
			.S(gen[5542]),
			.SE(gen[5543]),

			.SELF(gen[5447]),
			.cell_state(gen[5447])
		); 

/******************* CELL 5448 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5448 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5352]),
			.N(gen[5353]),
			.NE(gen[5354]),

			.O(gen[5447]),
			.E(gen[5449]),

			.SO(gen[5542]),
			.S(gen[5543]),
			.SE(gen[5544]),

			.SELF(gen[5448]),
			.cell_state(gen[5448])
		); 

/******************* CELL 5449 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5449 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5353]),
			.N(gen[5354]),
			.NE(gen[5355]),

			.O(gen[5448]),
			.E(gen[5450]),

			.SO(gen[5543]),
			.S(gen[5544]),
			.SE(gen[5545]),

			.SELF(gen[5449]),
			.cell_state(gen[5449])
		); 

/******************* CELL 5450 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5450 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5354]),
			.N(gen[5355]),
			.NE(gen[5356]),

			.O(gen[5449]),
			.E(gen[5451]),

			.SO(gen[5544]),
			.S(gen[5545]),
			.SE(gen[5546]),

			.SELF(gen[5450]),
			.cell_state(gen[5450])
		); 

/******************* CELL 5451 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5451 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5355]),
			.N(gen[5356]),
			.NE(gen[5357]),

			.O(gen[5450]),
			.E(gen[5452]),

			.SO(gen[5545]),
			.S(gen[5546]),
			.SE(gen[5547]),

			.SELF(gen[5451]),
			.cell_state(gen[5451])
		); 

/******************* CELL 5452 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5452 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5356]),
			.N(gen[5357]),
			.NE(gen[5358]),

			.O(gen[5451]),
			.E(gen[5453]),

			.SO(gen[5546]),
			.S(gen[5547]),
			.SE(gen[5548]),

			.SELF(gen[5452]),
			.cell_state(gen[5452])
		); 

/******************* CELL 5453 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5453 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5357]),
			.N(gen[5358]),
			.NE(gen[5359]),

			.O(gen[5452]),
			.E(gen[5454]),

			.SO(gen[5547]),
			.S(gen[5548]),
			.SE(gen[5549]),

			.SELF(gen[5453]),
			.cell_state(gen[5453])
		); 

/******************* CELL 5454 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5454 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5358]),
			.N(gen[5359]),
			.NE(gen[5360]),

			.O(gen[5453]),
			.E(gen[5455]),

			.SO(gen[5548]),
			.S(gen[5549]),
			.SE(gen[5550]),

			.SELF(gen[5454]),
			.cell_state(gen[5454])
		); 

/******************* CELL 5455 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5455 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5359]),
			.N(gen[5360]),
			.NE(gen[5361]),

			.O(gen[5454]),
			.E(gen[5456]),

			.SO(gen[5549]),
			.S(gen[5550]),
			.SE(gen[5551]),

			.SELF(gen[5455]),
			.cell_state(gen[5455])
		); 

/******************* CELL 5456 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5456 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5360]),
			.N(gen[5361]),
			.NE(gen[5362]),

			.O(gen[5455]),
			.E(gen[5457]),

			.SO(gen[5550]),
			.S(gen[5551]),
			.SE(gen[5552]),

			.SELF(gen[5456]),
			.cell_state(gen[5456])
		); 

/******************* CELL 5457 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5457 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5361]),
			.N(gen[5362]),
			.NE(gen[5363]),

			.O(gen[5456]),
			.E(gen[5458]),

			.SO(gen[5551]),
			.S(gen[5552]),
			.SE(gen[5553]),

			.SELF(gen[5457]),
			.cell_state(gen[5457])
		); 

/******************* CELL 5458 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5458 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5362]),
			.N(gen[5363]),
			.NE(gen[5364]),

			.O(gen[5457]),
			.E(gen[5459]),

			.SO(gen[5552]),
			.S(gen[5553]),
			.SE(gen[5554]),

			.SELF(gen[5458]),
			.cell_state(gen[5458])
		); 

/******************* CELL 5459 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5459 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5363]),
			.N(gen[5364]),
			.NE(gen[5365]),

			.O(gen[5458]),
			.E(gen[5460]),

			.SO(gen[5553]),
			.S(gen[5554]),
			.SE(gen[5555]),

			.SELF(gen[5459]),
			.cell_state(gen[5459])
		); 

/******************* CELL 5460 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5460 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5364]),
			.N(gen[5365]),
			.NE(gen[5366]),

			.O(gen[5459]),
			.E(gen[5461]),

			.SO(gen[5554]),
			.S(gen[5555]),
			.SE(gen[5556]),

			.SELF(gen[5460]),
			.cell_state(gen[5460])
		); 

/******************* CELL 5461 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5461 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5365]),
			.N(gen[5366]),
			.NE(gen[5367]),

			.O(gen[5460]),
			.E(gen[5462]),

			.SO(gen[5555]),
			.S(gen[5556]),
			.SE(gen[5557]),

			.SELF(gen[5461]),
			.cell_state(gen[5461])
		); 

/******************* CELL 5462 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5462 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5366]),
			.N(gen[5367]),
			.NE(gen[5368]),

			.O(gen[5461]),
			.E(gen[5463]),

			.SO(gen[5556]),
			.S(gen[5557]),
			.SE(gen[5558]),

			.SELF(gen[5462]),
			.cell_state(gen[5462])
		); 

/******************* CELL 5463 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5463 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5367]),
			.N(gen[5368]),
			.NE(gen[5369]),

			.O(gen[5462]),
			.E(gen[5464]),

			.SO(gen[5557]),
			.S(gen[5558]),
			.SE(gen[5559]),

			.SELF(gen[5463]),
			.cell_state(gen[5463])
		); 

/******************* CELL 5464 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5464 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5368]),
			.N(gen[5369]),
			.NE(gen[5370]),

			.O(gen[5463]),
			.E(gen[5465]),

			.SO(gen[5558]),
			.S(gen[5559]),
			.SE(gen[5560]),

			.SELF(gen[5464]),
			.cell_state(gen[5464])
		); 

/******************* CELL 5465 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5465 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5369]),
			.N(gen[5370]),
			.NE(gen[5371]),

			.O(gen[5464]),
			.E(gen[5466]),

			.SO(gen[5559]),
			.S(gen[5560]),
			.SE(gen[5561]),

			.SELF(gen[5465]),
			.cell_state(gen[5465])
		); 

/******************* CELL 5466 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5466 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5370]),
			.N(gen[5371]),
			.NE(gen[5372]),

			.O(gen[5465]),
			.E(gen[5467]),

			.SO(gen[5560]),
			.S(gen[5561]),
			.SE(gen[5562]),

			.SELF(gen[5466]),
			.cell_state(gen[5466])
		); 

/******************* CELL 5467 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5467 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5371]),
			.N(gen[5372]),
			.NE(gen[5373]),

			.O(gen[5466]),
			.E(gen[5468]),

			.SO(gen[5561]),
			.S(gen[5562]),
			.SE(gen[5563]),

			.SELF(gen[5467]),
			.cell_state(gen[5467])
		); 

/******************* CELL 5468 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5468 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5372]),
			.N(gen[5373]),
			.NE(gen[5374]),

			.O(gen[5467]),
			.E(gen[5469]),

			.SO(gen[5562]),
			.S(gen[5563]),
			.SE(gen[5564]),

			.SELF(gen[5468]),
			.cell_state(gen[5468])
		); 

/******************* CELL 5469 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5469 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5373]),
			.N(gen[5374]),
			.NE(gen[5375]),

			.O(gen[5468]),
			.E(gen[5470]),

			.SO(gen[5563]),
			.S(gen[5564]),
			.SE(gen[5565]),

			.SELF(gen[5469]),
			.cell_state(gen[5469])
		); 

/******************* CELL 5470 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5470 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5374]),
			.N(gen[5375]),
			.NE(gen[5376]),

			.O(gen[5469]),
			.E(gen[5471]),

			.SO(gen[5564]),
			.S(gen[5565]),
			.SE(gen[5566]),

			.SELF(gen[5470]),
			.cell_state(gen[5470])
		); 

/******************* CELL 5471 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5471 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5375]),
			.N(gen[5376]),
			.NE(gen[5377]),

			.O(gen[5470]),
			.E(gen[5472]),

			.SO(gen[5565]),
			.S(gen[5566]),
			.SE(gen[5567]),

			.SELF(gen[5471]),
			.cell_state(gen[5471])
		); 

/******************* CELL 5472 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5472 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5376]),
			.N(gen[5377]),
			.NE(gen[5378]),

			.O(gen[5471]),
			.E(gen[5473]),

			.SO(gen[5566]),
			.S(gen[5567]),
			.SE(gen[5568]),

			.SELF(gen[5472]),
			.cell_state(gen[5472])
		); 

/******************* CELL 5473 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5473 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5377]),
			.N(gen[5378]),
			.NE(gen[5379]),

			.O(gen[5472]),
			.E(gen[5474]),

			.SO(gen[5567]),
			.S(gen[5568]),
			.SE(gen[5569]),

			.SELF(gen[5473]),
			.cell_state(gen[5473])
		); 

/******************* CELL 5474 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5474 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5378]),
			.N(gen[5379]),
			.NE(gen[5380]),

			.O(gen[5473]),
			.E(gen[5475]),

			.SO(gen[5568]),
			.S(gen[5569]),
			.SE(gen[5570]),

			.SELF(gen[5474]),
			.cell_state(gen[5474])
		); 

/******************* CELL 5475 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5475 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5379]),
			.N(gen[5380]),
			.NE(gen[5381]),

			.O(gen[5474]),
			.E(gen[5476]),

			.SO(gen[5569]),
			.S(gen[5570]),
			.SE(gen[5571]),

			.SELF(gen[5475]),
			.cell_state(gen[5475])
		); 

/******************* CELL 5476 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5476 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5380]),
			.N(gen[5381]),
			.NE(gen[5382]),

			.O(gen[5475]),
			.E(gen[5477]),

			.SO(gen[5570]),
			.S(gen[5571]),
			.SE(gen[5572]),

			.SELF(gen[5476]),
			.cell_state(gen[5476])
		); 

/******************* CELL 5477 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5477 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5381]),
			.N(gen[5382]),
			.NE(gen[5383]),

			.O(gen[5476]),
			.E(gen[5478]),

			.SO(gen[5571]),
			.S(gen[5572]),
			.SE(gen[5573]),

			.SELF(gen[5477]),
			.cell_state(gen[5477])
		); 

/******************* CELL 5478 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5478 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5382]),
			.N(gen[5383]),
			.NE(gen[5384]),

			.O(gen[5477]),
			.E(gen[5479]),

			.SO(gen[5572]),
			.S(gen[5573]),
			.SE(gen[5574]),

			.SELF(gen[5478]),
			.cell_state(gen[5478])
		); 

/******************* CELL 5479 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5479 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5383]),
			.N(gen[5384]),
			.NE(gen[5385]),

			.O(gen[5478]),
			.E(gen[5480]),

			.SO(gen[5573]),
			.S(gen[5574]),
			.SE(gen[5575]),

			.SELF(gen[5479]),
			.cell_state(gen[5479])
		); 

/******************* CELL 5480 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5480 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5384]),
			.N(gen[5385]),
			.NE(gen[5386]),

			.O(gen[5479]),
			.E(gen[5481]),

			.SO(gen[5574]),
			.S(gen[5575]),
			.SE(gen[5576]),

			.SELF(gen[5480]),
			.cell_state(gen[5480])
		); 

/******************* CELL 5481 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5481 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5385]),
			.N(gen[5386]),
			.NE(gen[5387]),

			.O(gen[5480]),
			.E(gen[5482]),

			.SO(gen[5575]),
			.S(gen[5576]),
			.SE(gen[5577]),

			.SELF(gen[5481]),
			.cell_state(gen[5481])
		); 

/******************* CELL 5482 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5482 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5386]),
			.N(gen[5387]),
			.NE(gen[5388]),

			.O(gen[5481]),
			.E(gen[5483]),

			.SO(gen[5576]),
			.S(gen[5577]),
			.SE(gen[5578]),

			.SELF(gen[5482]),
			.cell_state(gen[5482])
		); 

/******************* CELL 5483 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5483 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5387]),
			.N(gen[5388]),
			.NE(gen[5389]),

			.O(gen[5482]),
			.E(gen[5484]),

			.SO(gen[5577]),
			.S(gen[5578]),
			.SE(gen[5579]),

			.SELF(gen[5483]),
			.cell_state(gen[5483])
		); 

/******************* CELL 5484 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5484 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5388]),
			.N(gen[5389]),
			.NE(gen[5390]),

			.O(gen[5483]),
			.E(gen[5485]),

			.SO(gen[5578]),
			.S(gen[5579]),
			.SE(gen[5580]),

			.SELF(gen[5484]),
			.cell_state(gen[5484])
		); 

/******************* CELL 5485 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5485 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5389]),
			.N(gen[5390]),
			.NE(gen[5391]),

			.O(gen[5484]),
			.E(gen[5486]),

			.SO(gen[5579]),
			.S(gen[5580]),
			.SE(gen[5581]),

			.SELF(gen[5485]),
			.cell_state(gen[5485])
		); 

/******************* CELL 5486 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5486 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5390]),
			.N(gen[5391]),
			.NE(gen[5392]),

			.O(gen[5485]),
			.E(gen[5487]),

			.SO(gen[5580]),
			.S(gen[5581]),
			.SE(gen[5582]),

			.SELF(gen[5486]),
			.cell_state(gen[5486])
		); 

/******************* CELL 5487 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5487 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5391]),
			.N(gen[5392]),
			.NE(gen[5393]),

			.O(gen[5486]),
			.E(gen[5488]),

			.SO(gen[5581]),
			.S(gen[5582]),
			.SE(gen[5583]),

			.SELF(gen[5487]),
			.cell_state(gen[5487])
		); 

/******************* CELL 5488 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5488 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5392]),
			.N(gen[5393]),
			.NE(gen[5394]),

			.O(gen[5487]),
			.E(gen[5489]),

			.SO(gen[5582]),
			.S(gen[5583]),
			.SE(gen[5584]),

			.SELF(gen[5488]),
			.cell_state(gen[5488])
		); 

/******************* CELL 5489 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5489 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5393]),
			.N(gen[5394]),
			.NE(gen[5395]),

			.O(gen[5488]),
			.E(gen[5490]),

			.SO(gen[5583]),
			.S(gen[5584]),
			.SE(gen[5585]),

			.SELF(gen[5489]),
			.cell_state(gen[5489])
		); 

/******************* CELL 5490 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5490 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5394]),
			.N(gen[5395]),
			.NE(gen[5396]),

			.O(gen[5489]),
			.E(gen[5491]),

			.SO(gen[5584]),
			.S(gen[5585]),
			.SE(gen[5586]),

			.SELF(gen[5490]),
			.cell_state(gen[5490])
		); 

/******************* CELL 5491 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5491 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5395]),
			.N(gen[5396]),
			.NE(gen[5397]),

			.O(gen[5490]),
			.E(gen[5492]),

			.SO(gen[5585]),
			.S(gen[5586]),
			.SE(gen[5587]),

			.SELF(gen[5491]),
			.cell_state(gen[5491])
		); 

/******************* CELL 5492 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5492 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5396]),
			.N(gen[5397]),
			.NE(gen[5398]),

			.O(gen[5491]),
			.E(gen[5493]),

			.SO(gen[5586]),
			.S(gen[5587]),
			.SE(gen[5588]),

			.SELF(gen[5492]),
			.cell_state(gen[5492])
		); 

/******************* CELL 5493 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5493 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5397]),
			.N(gen[5398]),
			.NE(gen[5399]),

			.O(gen[5492]),
			.E(gen[5494]),

			.SO(gen[5587]),
			.S(gen[5588]),
			.SE(gen[5589]),

			.SELF(gen[5493]),
			.cell_state(gen[5493])
		); 

/******************* CELL 5494 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5494 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5398]),
			.N(gen[5399]),
			.NE(gen[5400]),

			.O(gen[5493]),
			.E(gen[5495]),

			.SO(gen[5588]),
			.S(gen[5589]),
			.SE(gen[5590]),

			.SELF(gen[5494]),
			.cell_state(gen[5494])
		); 

/******************* CELL 5495 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5495 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5399]),
			.N(gen[5400]),
			.NE(gen[5401]),

			.O(gen[5494]),
			.E(gen[5496]),

			.SO(gen[5589]),
			.S(gen[5590]),
			.SE(gen[5591]),

			.SELF(gen[5495]),
			.cell_state(gen[5495])
		); 

/******************* CELL 5496 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5496 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5400]),
			.N(gen[5401]),
			.NE(gen[5402]),

			.O(gen[5495]),
			.E(gen[5497]),

			.SO(gen[5590]),
			.S(gen[5591]),
			.SE(gen[5592]),

			.SELF(gen[5496]),
			.cell_state(gen[5496])
		); 

/******************* CELL 5497 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5497 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5401]),
			.N(gen[5402]),
			.NE(gen[5403]),

			.O(gen[5496]),
			.E(gen[5498]),

			.SO(gen[5591]),
			.S(gen[5592]),
			.SE(gen[5593]),

			.SELF(gen[5497]),
			.cell_state(gen[5497])
		); 

/******************* CELL 5498 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5498 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5402]),
			.N(gen[5403]),
			.NE(gen[5404]),

			.O(gen[5497]),
			.E(gen[5499]),

			.SO(gen[5592]),
			.S(gen[5593]),
			.SE(gen[5594]),

			.SELF(gen[5498]),
			.cell_state(gen[5498])
		); 

/******************* CELL 5499 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5499 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5403]),
			.N(gen[5404]),
			.NE(gen[5405]),

			.O(gen[5498]),
			.E(gen[5500]),

			.SO(gen[5593]),
			.S(gen[5594]),
			.SE(gen[5595]),

			.SELF(gen[5499]),
			.cell_state(gen[5499])
		); 

/******************* CELL 5500 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5500 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5404]),
			.N(gen[5405]),
			.NE(gen[5406]),

			.O(gen[5499]),
			.E(gen[5501]),

			.SO(gen[5594]),
			.S(gen[5595]),
			.SE(gen[5596]),

			.SELF(gen[5500]),
			.cell_state(gen[5500])
		); 

/******************* CELL 5501 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5501 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5405]),
			.N(gen[5406]),
			.NE(gen[5407]),

			.O(gen[5500]),
			.E(gen[5502]),

			.SO(gen[5595]),
			.S(gen[5596]),
			.SE(gen[5597]),

			.SELF(gen[5501]),
			.cell_state(gen[5501])
		); 

/******************* CELL 5502 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5502 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5406]),
			.N(gen[5407]),
			.NE(gen[5408]),

			.O(gen[5501]),
			.E(gen[5503]),

			.SO(gen[5596]),
			.S(gen[5597]),
			.SE(gen[5598]),

			.SELF(gen[5502]),
			.cell_state(gen[5502])
		); 

/******************* CELL 5503 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5503 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5407]),
			.N(gen[5408]),
			.NE(gen[5409]),

			.O(gen[5502]),
			.E(gen[5504]),

			.SO(gen[5597]),
			.S(gen[5598]),
			.SE(gen[5599]),

			.SELF(gen[5503]),
			.cell_state(gen[5503])
		); 

/******************* CELL 5504 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5504 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5408]),
			.N(gen[5409]),
			.NE(gen[5410]),

			.O(gen[5503]),
			.E(gen[5505]),

			.SO(gen[5598]),
			.S(gen[5599]),
			.SE(gen[5600]),

			.SELF(gen[5504]),
			.cell_state(gen[5504])
		); 

/******************* CELL 5505 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5505 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5409]),
			.N(gen[5410]),
			.NE(gen[5411]),

			.O(gen[5504]),
			.E(gen[5506]),

			.SO(gen[5599]),
			.S(gen[5600]),
			.SE(gen[5601]),

			.SELF(gen[5505]),
			.cell_state(gen[5505])
		); 

/******************* CELL 5506 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5506 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5410]),
			.N(gen[5411]),
			.NE(gen[5412]),

			.O(gen[5505]),
			.E(gen[5507]),

			.SO(gen[5600]),
			.S(gen[5601]),
			.SE(gen[5602]),

			.SELF(gen[5506]),
			.cell_state(gen[5506])
		); 

/******************* CELL 5507 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5507 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5411]),
			.N(gen[5412]),
			.NE(gen[5413]),

			.O(gen[5506]),
			.E(gen[5508]),

			.SO(gen[5601]),
			.S(gen[5602]),
			.SE(gen[5603]),

			.SELF(gen[5507]),
			.cell_state(gen[5507])
		); 

/******************* CELL 5508 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5508 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5412]),
			.N(gen[5413]),
			.NE(gen[5414]),

			.O(gen[5507]),
			.E(gen[5509]),

			.SO(gen[5602]),
			.S(gen[5603]),
			.SE(gen[5604]),

			.SELF(gen[5508]),
			.cell_state(gen[5508])
		); 

/******************* CELL 5509 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5509 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5413]),
			.N(gen[5414]),
			.NE(gen[5413]),

			.O(gen[5508]),
			.E(gen[5508]),

			.SO(gen[5603]),
			.S(gen[5604]),
			.SE(gen[5603]),

			.SELF(gen[5509]),
			.cell_state(gen[5509])
		); 

/******************* CELL 5510 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5510 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5416]),
			.N(gen[5415]),
			.NE(gen[5416]),

			.O(gen[5511]),
			.E(gen[5511]),

			.SO(gen[5606]),
			.S(gen[5605]),
			.SE(gen[5606]),

			.SELF(gen[5510]),
			.cell_state(gen[5510])
		); 

/******************* CELL 5511 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5511 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5415]),
			.N(gen[5416]),
			.NE(gen[5417]),

			.O(gen[5510]),
			.E(gen[5512]),

			.SO(gen[5605]),
			.S(gen[5606]),
			.SE(gen[5607]),

			.SELF(gen[5511]),
			.cell_state(gen[5511])
		); 

/******************* CELL 5512 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5512 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5416]),
			.N(gen[5417]),
			.NE(gen[5418]),

			.O(gen[5511]),
			.E(gen[5513]),

			.SO(gen[5606]),
			.S(gen[5607]),
			.SE(gen[5608]),

			.SELF(gen[5512]),
			.cell_state(gen[5512])
		); 

/******************* CELL 5513 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5513 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5417]),
			.N(gen[5418]),
			.NE(gen[5419]),

			.O(gen[5512]),
			.E(gen[5514]),

			.SO(gen[5607]),
			.S(gen[5608]),
			.SE(gen[5609]),

			.SELF(gen[5513]),
			.cell_state(gen[5513])
		); 

/******************* CELL 5514 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5514 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5418]),
			.N(gen[5419]),
			.NE(gen[5420]),

			.O(gen[5513]),
			.E(gen[5515]),

			.SO(gen[5608]),
			.S(gen[5609]),
			.SE(gen[5610]),

			.SELF(gen[5514]),
			.cell_state(gen[5514])
		); 

/******************* CELL 5515 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5515 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5419]),
			.N(gen[5420]),
			.NE(gen[5421]),

			.O(gen[5514]),
			.E(gen[5516]),

			.SO(gen[5609]),
			.S(gen[5610]),
			.SE(gen[5611]),

			.SELF(gen[5515]),
			.cell_state(gen[5515])
		); 

/******************* CELL 5516 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5516 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5420]),
			.N(gen[5421]),
			.NE(gen[5422]),

			.O(gen[5515]),
			.E(gen[5517]),

			.SO(gen[5610]),
			.S(gen[5611]),
			.SE(gen[5612]),

			.SELF(gen[5516]),
			.cell_state(gen[5516])
		); 

/******************* CELL 5517 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5517 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5421]),
			.N(gen[5422]),
			.NE(gen[5423]),

			.O(gen[5516]),
			.E(gen[5518]),

			.SO(gen[5611]),
			.S(gen[5612]),
			.SE(gen[5613]),

			.SELF(gen[5517]),
			.cell_state(gen[5517])
		); 

/******************* CELL 5518 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5518 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5422]),
			.N(gen[5423]),
			.NE(gen[5424]),

			.O(gen[5517]),
			.E(gen[5519]),

			.SO(gen[5612]),
			.S(gen[5613]),
			.SE(gen[5614]),

			.SELF(gen[5518]),
			.cell_state(gen[5518])
		); 

/******************* CELL 5519 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5519 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5423]),
			.N(gen[5424]),
			.NE(gen[5425]),

			.O(gen[5518]),
			.E(gen[5520]),

			.SO(gen[5613]),
			.S(gen[5614]),
			.SE(gen[5615]),

			.SELF(gen[5519]),
			.cell_state(gen[5519])
		); 

/******************* CELL 5520 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5520 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5424]),
			.N(gen[5425]),
			.NE(gen[5426]),

			.O(gen[5519]),
			.E(gen[5521]),

			.SO(gen[5614]),
			.S(gen[5615]),
			.SE(gen[5616]),

			.SELF(gen[5520]),
			.cell_state(gen[5520])
		); 

/******************* CELL 5521 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5521 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5425]),
			.N(gen[5426]),
			.NE(gen[5427]),

			.O(gen[5520]),
			.E(gen[5522]),

			.SO(gen[5615]),
			.S(gen[5616]),
			.SE(gen[5617]),

			.SELF(gen[5521]),
			.cell_state(gen[5521])
		); 

/******************* CELL 5522 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5522 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5426]),
			.N(gen[5427]),
			.NE(gen[5428]),

			.O(gen[5521]),
			.E(gen[5523]),

			.SO(gen[5616]),
			.S(gen[5617]),
			.SE(gen[5618]),

			.SELF(gen[5522]),
			.cell_state(gen[5522])
		); 

/******************* CELL 5523 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5523 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5427]),
			.N(gen[5428]),
			.NE(gen[5429]),

			.O(gen[5522]),
			.E(gen[5524]),

			.SO(gen[5617]),
			.S(gen[5618]),
			.SE(gen[5619]),

			.SELF(gen[5523]),
			.cell_state(gen[5523])
		); 

/******************* CELL 5524 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5524 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5428]),
			.N(gen[5429]),
			.NE(gen[5430]),

			.O(gen[5523]),
			.E(gen[5525]),

			.SO(gen[5618]),
			.S(gen[5619]),
			.SE(gen[5620]),

			.SELF(gen[5524]),
			.cell_state(gen[5524])
		); 

/******************* CELL 5525 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5525 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5429]),
			.N(gen[5430]),
			.NE(gen[5431]),

			.O(gen[5524]),
			.E(gen[5526]),

			.SO(gen[5619]),
			.S(gen[5620]),
			.SE(gen[5621]),

			.SELF(gen[5525]),
			.cell_state(gen[5525])
		); 

/******************* CELL 5526 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5526 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5430]),
			.N(gen[5431]),
			.NE(gen[5432]),

			.O(gen[5525]),
			.E(gen[5527]),

			.SO(gen[5620]),
			.S(gen[5621]),
			.SE(gen[5622]),

			.SELF(gen[5526]),
			.cell_state(gen[5526])
		); 

/******************* CELL 5527 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5527 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5431]),
			.N(gen[5432]),
			.NE(gen[5433]),

			.O(gen[5526]),
			.E(gen[5528]),

			.SO(gen[5621]),
			.S(gen[5622]),
			.SE(gen[5623]),

			.SELF(gen[5527]),
			.cell_state(gen[5527])
		); 

/******************* CELL 5528 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5528 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5432]),
			.N(gen[5433]),
			.NE(gen[5434]),

			.O(gen[5527]),
			.E(gen[5529]),

			.SO(gen[5622]),
			.S(gen[5623]),
			.SE(gen[5624]),

			.SELF(gen[5528]),
			.cell_state(gen[5528])
		); 

/******************* CELL 5529 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5529 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5433]),
			.N(gen[5434]),
			.NE(gen[5435]),

			.O(gen[5528]),
			.E(gen[5530]),

			.SO(gen[5623]),
			.S(gen[5624]),
			.SE(gen[5625]),

			.SELF(gen[5529]),
			.cell_state(gen[5529])
		); 

/******************* CELL 5530 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5530 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5434]),
			.N(gen[5435]),
			.NE(gen[5436]),

			.O(gen[5529]),
			.E(gen[5531]),

			.SO(gen[5624]),
			.S(gen[5625]),
			.SE(gen[5626]),

			.SELF(gen[5530]),
			.cell_state(gen[5530])
		); 

/******************* CELL 5531 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5531 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5435]),
			.N(gen[5436]),
			.NE(gen[5437]),

			.O(gen[5530]),
			.E(gen[5532]),

			.SO(gen[5625]),
			.S(gen[5626]),
			.SE(gen[5627]),

			.SELF(gen[5531]),
			.cell_state(gen[5531])
		); 

/******************* CELL 5532 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5532 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5436]),
			.N(gen[5437]),
			.NE(gen[5438]),

			.O(gen[5531]),
			.E(gen[5533]),

			.SO(gen[5626]),
			.S(gen[5627]),
			.SE(gen[5628]),

			.SELF(gen[5532]),
			.cell_state(gen[5532])
		); 

/******************* CELL 5533 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5533 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5437]),
			.N(gen[5438]),
			.NE(gen[5439]),

			.O(gen[5532]),
			.E(gen[5534]),

			.SO(gen[5627]),
			.S(gen[5628]),
			.SE(gen[5629]),

			.SELF(gen[5533]),
			.cell_state(gen[5533])
		); 

/******************* CELL 5534 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5534 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5438]),
			.N(gen[5439]),
			.NE(gen[5440]),

			.O(gen[5533]),
			.E(gen[5535]),

			.SO(gen[5628]),
			.S(gen[5629]),
			.SE(gen[5630]),

			.SELF(gen[5534]),
			.cell_state(gen[5534])
		); 

/******************* CELL 5535 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5535 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5439]),
			.N(gen[5440]),
			.NE(gen[5441]),

			.O(gen[5534]),
			.E(gen[5536]),

			.SO(gen[5629]),
			.S(gen[5630]),
			.SE(gen[5631]),

			.SELF(gen[5535]),
			.cell_state(gen[5535])
		); 

/******************* CELL 5536 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5536 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5440]),
			.N(gen[5441]),
			.NE(gen[5442]),

			.O(gen[5535]),
			.E(gen[5537]),

			.SO(gen[5630]),
			.S(gen[5631]),
			.SE(gen[5632]),

			.SELF(gen[5536]),
			.cell_state(gen[5536])
		); 

/******************* CELL 5537 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5537 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5441]),
			.N(gen[5442]),
			.NE(gen[5443]),

			.O(gen[5536]),
			.E(gen[5538]),

			.SO(gen[5631]),
			.S(gen[5632]),
			.SE(gen[5633]),

			.SELF(gen[5537]),
			.cell_state(gen[5537])
		); 

/******************* CELL 5538 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5538 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5442]),
			.N(gen[5443]),
			.NE(gen[5444]),

			.O(gen[5537]),
			.E(gen[5539]),

			.SO(gen[5632]),
			.S(gen[5633]),
			.SE(gen[5634]),

			.SELF(gen[5538]),
			.cell_state(gen[5538])
		); 

/******************* CELL 5539 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5539 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5443]),
			.N(gen[5444]),
			.NE(gen[5445]),

			.O(gen[5538]),
			.E(gen[5540]),

			.SO(gen[5633]),
			.S(gen[5634]),
			.SE(gen[5635]),

			.SELF(gen[5539]),
			.cell_state(gen[5539])
		); 

/******************* CELL 5540 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5540 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5444]),
			.N(gen[5445]),
			.NE(gen[5446]),

			.O(gen[5539]),
			.E(gen[5541]),

			.SO(gen[5634]),
			.S(gen[5635]),
			.SE(gen[5636]),

			.SELF(gen[5540]),
			.cell_state(gen[5540])
		); 

/******************* CELL 5541 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5541 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5445]),
			.N(gen[5446]),
			.NE(gen[5447]),

			.O(gen[5540]),
			.E(gen[5542]),

			.SO(gen[5635]),
			.S(gen[5636]),
			.SE(gen[5637]),

			.SELF(gen[5541]),
			.cell_state(gen[5541])
		); 

/******************* CELL 5542 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5542 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5446]),
			.N(gen[5447]),
			.NE(gen[5448]),

			.O(gen[5541]),
			.E(gen[5543]),

			.SO(gen[5636]),
			.S(gen[5637]),
			.SE(gen[5638]),

			.SELF(gen[5542]),
			.cell_state(gen[5542])
		); 

/******************* CELL 5543 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5543 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5447]),
			.N(gen[5448]),
			.NE(gen[5449]),

			.O(gen[5542]),
			.E(gen[5544]),

			.SO(gen[5637]),
			.S(gen[5638]),
			.SE(gen[5639]),

			.SELF(gen[5543]),
			.cell_state(gen[5543])
		); 

/******************* CELL 5544 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5544 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5448]),
			.N(gen[5449]),
			.NE(gen[5450]),

			.O(gen[5543]),
			.E(gen[5545]),

			.SO(gen[5638]),
			.S(gen[5639]),
			.SE(gen[5640]),

			.SELF(gen[5544]),
			.cell_state(gen[5544])
		); 

/******************* CELL 5545 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5545 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5449]),
			.N(gen[5450]),
			.NE(gen[5451]),

			.O(gen[5544]),
			.E(gen[5546]),

			.SO(gen[5639]),
			.S(gen[5640]),
			.SE(gen[5641]),

			.SELF(gen[5545]),
			.cell_state(gen[5545])
		); 

/******************* CELL 5546 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5546 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5450]),
			.N(gen[5451]),
			.NE(gen[5452]),

			.O(gen[5545]),
			.E(gen[5547]),

			.SO(gen[5640]),
			.S(gen[5641]),
			.SE(gen[5642]),

			.SELF(gen[5546]),
			.cell_state(gen[5546])
		); 

/******************* CELL 5547 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5547 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5451]),
			.N(gen[5452]),
			.NE(gen[5453]),

			.O(gen[5546]),
			.E(gen[5548]),

			.SO(gen[5641]),
			.S(gen[5642]),
			.SE(gen[5643]),

			.SELF(gen[5547]),
			.cell_state(gen[5547])
		); 

/******************* CELL 5548 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5548 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5452]),
			.N(gen[5453]),
			.NE(gen[5454]),

			.O(gen[5547]),
			.E(gen[5549]),

			.SO(gen[5642]),
			.S(gen[5643]),
			.SE(gen[5644]),

			.SELF(gen[5548]),
			.cell_state(gen[5548])
		); 

/******************* CELL 5549 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5549 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5453]),
			.N(gen[5454]),
			.NE(gen[5455]),

			.O(gen[5548]),
			.E(gen[5550]),

			.SO(gen[5643]),
			.S(gen[5644]),
			.SE(gen[5645]),

			.SELF(gen[5549]),
			.cell_state(gen[5549])
		); 

/******************* CELL 5550 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5550 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5454]),
			.N(gen[5455]),
			.NE(gen[5456]),

			.O(gen[5549]),
			.E(gen[5551]),

			.SO(gen[5644]),
			.S(gen[5645]),
			.SE(gen[5646]),

			.SELF(gen[5550]),
			.cell_state(gen[5550])
		); 

/******************* CELL 5551 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5551 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5455]),
			.N(gen[5456]),
			.NE(gen[5457]),

			.O(gen[5550]),
			.E(gen[5552]),

			.SO(gen[5645]),
			.S(gen[5646]),
			.SE(gen[5647]),

			.SELF(gen[5551]),
			.cell_state(gen[5551])
		); 

/******************* CELL 5552 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5552 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5456]),
			.N(gen[5457]),
			.NE(gen[5458]),

			.O(gen[5551]),
			.E(gen[5553]),

			.SO(gen[5646]),
			.S(gen[5647]),
			.SE(gen[5648]),

			.SELF(gen[5552]),
			.cell_state(gen[5552])
		); 

/******************* CELL 5553 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5553 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5457]),
			.N(gen[5458]),
			.NE(gen[5459]),

			.O(gen[5552]),
			.E(gen[5554]),

			.SO(gen[5647]),
			.S(gen[5648]),
			.SE(gen[5649]),

			.SELF(gen[5553]),
			.cell_state(gen[5553])
		); 

/******************* CELL 5554 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5554 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5458]),
			.N(gen[5459]),
			.NE(gen[5460]),

			.O(gen[5553]),
			.E(gen[5555]),

			.SO(gen[5648]),
			.S(gen[5649]),
			.SE(gen[5650]),

			.SELF(gen[5554]),
			.cell_state(gen[5554])
		); 

/******************* CELL 5555 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5555 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5459]),
			.N(gen[5460]),
			.NE(gen[5461]),

			.O(gen[5554]),
			.E(gen[5556]),

			.SO(gen[5649]),
			.S(gen[5650]),
			.SE(gen[5651]),

			.SELF(gen[5555]),
			.cell_state(gen[5555])
		); 

/******************* CELL 5556 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5556 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5460]),
			.N(gen[5461]),
			.NE(gen[5462]),

			.O(gen[5555]),
			.E(gen[5557]),

			.SO(gen[5650]),
			.S(gen[5651]),
			.SE(gen[5652]),

			.SELF(gen[5556]),
			.cell_state(gen[5556])
		); 

/******************* CELL 5557 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5557 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5461]),
			.N(gen[5462]),
			.NE(gen[5463]),

			.O(gen[5556]),
			.E(gen[5558]),

			.SO(gen[5651]),
			.S(gen[5652]),
			.SE(gen[5653]),

			.SELF(gen[5557]),
			.cell_state(gen[5557])
		); 

/******************* CELL 5558 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5558 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5462]),
			.N(gen[5463]),
			.NE(gen[5464]),

			.O(gen[5557]),
			.E(gen[5559]),

			.SO(gen[5652]),
			.S(gen[5653]),
			.SE(gen[5654]),

			.SELF(gen[5558]),
			.cell_state(gen[5558])
		); 

/******************* CELL 5559 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5559 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5463]),
			.N(gen[5464]),
			.NE(gen[5465]),

			.O(gen[5558]),
			.E(gen[5560]),

			.SO(gen[5653]),
			.S(gen[5654]),
			.SE(gen[5655]),

			.SELF(gen[5559]),
			.cell_state(gen[5559])
		); 

/******************* CELL 5560 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5560 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5464]),
			.N(gen[5465]),
			.NE(gen[5466]),

			.O(gen[5559]),
			.E(gen[5561]),

			.SO(gen[5654]),
			.S(gen[5655]),
			.SE(gen[5656]),

			.SELF(gen[5560]),
			.cell_state(gen[5560])
		); 

/******************* CELL 5561 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5561 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5465]),
			.N(gen[5466]),
			.NE(gen[5467]),

			.O(gen[5560]),
			.E(gen[5562]),

			.SO(gen[5655]),
			.S(gen[5656]),
			.SE(gen[5657]),

			.SELF(gen[5561]),
			.cell_state(gen[5561])
		); 

/******************* CELL 5562 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5562 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5466]),
			.N(gen[5467]),
			.NE(gen[5468]),

			.O(gen[5561]),
			.E(gen[5563]),

			.SO(gen[5656]),
			.S(gen[5657]),
			.SE(gen[5658]),

			.SELF(gen[5562]),
			.cell_state(gen[5562])
		); 

/******************* CELL 5563 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5563 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5467]),
			.N(gen[5468]),
			.NE(gen[5469]),

			.O(gen[5562]),
			.E(gen[5564]),

			.SO(gen[5657]),
			.S(gen[5658]),
			.SE(gen[5659]),

			.SELF(gen[5563]),
			.cell_state(gen[5563])
		); 

/******************* CELL 5564 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5564 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5468]),
			.N(gen[5469]),
			.NE(gen[5470]),

			.O(gen[5563]),
			.E(gen[5565]),

			.SO(gen[5658]),
			.S(gen[5659]),
			.SE(gen[5660]),

			.SELF(gen[5564]),
			.cell_state(gen[5564])
		); 

/******************* CELL 5565 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5565 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5469]),
			.N(gen[5470]),
			.NE(gen[5471]),

			.O(gen[5564]),
			.E(gen[5566]),

			.SO(gen[5659]),
			.S(gen[5660]),
			.SE(gen[5661]),

			.SELF(gen[5565]),
			.cell_state(gen[5565])
		); 

/******************* CELL 5566 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5566 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5470]),
			.N(gen[5471]),
			.NE(gen[5472]),

			.O(gen[5565]),
			.E(gen[5567]),

			.SO(gen[5660]),
			.S(gen[5661]),
			.SE(gen[5662]),

			.SELF(gen[5566]),
			.cell_state(gen[5566])
		); 

/******************* CELL 5567 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5567 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5471]),
			.N(gen[5472]),
			.NE(gen[5473]),

			.O(gen[5566]),
			.E(gen[5568]),

			.SO(gen[5661]),
			.S(gen[5662]),
			.SE(gen[5663]),

			.SELF(gen[5567]),
			.cell_state(gen[5567])
		); 

/******************* CELL 5568 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5568 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5472]),
			.N(gen[5473]),
			.NE(gen[5474]),

			.O(gen[5567]),
			.E(gen[5569]),

			.SO(gen[5662]),
			.S(gen[5663]),
			.SE(gen[5664]),

			.SELF(gen[5568]),
			.cell_state(gen[5568])
		); 

/******************* CELL 5569 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5569 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5473]),
			.N(gen[5474]),
			.NE(gen[5475]),

			.O(gen[5568]),
			.E(gen[5570]),

			.SO(gen[5663]),
			.S(gen[5664]),
			.SE(gen[5665]),

			.SELF(gen[5569]),
			.cell_state(gen[5569])
		); 

/******************* CELL 5570 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5570 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5474]),
			.N(gen[5475]),
			.NE(gen[5476]),

			.O(gen[5569]),
			.E(gen[5571]),

			.SO(gen[5664]),
			.S(gen[5665]),
			.SE(gen[5666]),

			.SELF(gen[5570]),
			.cell_state(gen[5570])
		); 

/******************* CELL 5571 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5571 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5475]),
			.N(gen[5476]),
			.NE(gen[5477]),

			.O(gen[5570]),
			.E(gen[5572]),

			.SO(gen[5665]),
			.S(gen[5666]),
			.SE(gen[5667]),

			.SELF(gen[5571]),
			.cell_state(gen[5571])
		); 

/******************* CELL 5572 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5572 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5476]),
			.N(gen[5477]),
			.NE(gen[5478]),

			.O(gen[5571]),
			.E(gen[5573]),

			.SO(gen[5666]),
			.S(gen[5667]),
			.SE(gen[5668]),

			.SELF(gen[5572]),
			.cell_state(gen[5572])
		); 

/******************* CELL 5573 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5573 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5477]),
			.N(gen[5478]),
			.NE(gen[5479]),

			.O(gen[5572]),
			.E(gen[5574]),

			.SO(gen[5667]),
			.S(gen[5668]),
			.SE(gen[5669]),

			.SELF(gen[5573]),
			.cell_state(gen[5573])
		); 

/******************* CELL 5574 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5574 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5478]),
			.N(gen[5479]),
			.NE(gen[5480]),

			.O(gen[5573]),
			.E(gen[5575]),

			.SO(gen[5668]),
			.S(gen[5669]),
			.SE(gen[5670]),

			.SELF(gen[5574]),
			.cell_state(gen[5574])
		); 

/******************* CELL 5575 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5575 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5479]),
			.N(gen[5480]),
			.NE(gen[5481]),

			.O(gen[5574]),
			.E(gen[5576]),

			.SO(gen[5669]),
			.S(gen[5670]),
			.SE(gen[5671]),

			.SELF(gen[5575]),
			.cell_state(gen[5575])
		); 

/******************* CELL 5576 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5576 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5480]),
			.N(gen[5481]),
			.NE(gen[5482]),

			.O(gen[5575]),
			.E(gen[5577]),

			.SO(gen[5670]),
			.S(gen[5671]),
			.SE(gen[5672]),

			.SELF(gen[5576]),
			.cell_state(gen[5576])
		); 

/******************* CELL 5577 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5577 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5481]),
			.N(gen[5482]),
			.NE(gen[5483]),

			.O(gen[5576]),
			.E(gen[5578]),

			.SO(gen[5671]),
			.S(gen[5672]),
			.SE(gen[5673]),

			.SELF(gen[5577]),
			.cell_state(gen[5577])
		); 

/******************* CELL 5578 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5578 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5482]),
			.N(gen[5483]),
			.NE(gen[5484]),

			.O(gen[5577]),
			.E(gen[5579]),

			.SO(gen[5672]),
			.S(gen[5673]),
			.SE(gen[5674]),

			.SELF(gen[5578]),
			.cell_state(gen[5578])
		); 

/******************* CELL 5579 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5579 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5483]),
			.N(gen[5484]),
			.NE(gen[5485]),

			.O(gen[5578]),
			.E(gen[5580]),

			.SO(gen[5673]),
			.S(gen[5674]),
			.SE(gen[5675]),

			.SELF(gen[5579]),
			.cell_state(gen[5579])
		); 

/******************* CELL 5580 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5580 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5484]),
			.N(gen[5485]),
			.NE(gen[5486]),

			.O(gen[5579]),
			.E(gen[5581]),

			.SO(gen[5674]),
			.S(gen[5675]),
			.SE(gen[5676]),

			.SELF(gen[5580]),
			.cell_state(gen[5580])
		); 

/******************* CELL 5581 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5581 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5485]),
			.N(gen[5486]),
			.NE(gen[5487]),

			.O(gen[5580]),
			.E(gen[5582]),

			.SO(gen[5675]),
			.S(gen[5676]),
			.SE(gen[5677]),

			.SELF(gen[5581]),
			.cell_state(gen[5581])
		); 

/******************* CELL 5582 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5582 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5486]),
			.N(gen[5487]),
			.NE(gen[5488]),

			.O(gen[5581]),
			.E(gen[5583]),

			.SO(gen[5676]),
			.S(gen[5677]),
			.SE(gen[5678]),

			.SELF(gen[5582]),
			.cell_state(gen[5582])
		); 

/******************* CELL 5583 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5583 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5487]),
			.N(gen[5488]),
			.NE(gen[5489]),

			.O(gen[5582]),
			.E(gen[5584]),

			.SO(gen[5677]),
			.S(gen[5678]),
			.SE(gen[5679]),

			.SELF(gen[5583]),
			.cell_state(gen[5583])
		); 

/******************* CELL 5584 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5584 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5488]),
			.N(gen[5489]),
			.NE(gen[5490]),

			.O(gen[5583]),
			.E(gen[5585]),

			.SO(gen[5678]),
			.S(gen[5679]),
			.SE(gen[5680]),

			.SELF(gen[5584]),
			.cell_state(gen[5584])
		); 

/******************* CELL 5585 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5585 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5489]),
			.N(gen[5490]),
			.NE(gen[5491]),

			.O(gen[5584]),
			.E(gen[5586]),

			.SO(gen[5679]),
			.S(gen[5680]),
			.SE(gen[5681]),

			.SELF(gen[5585]),
			.cell_state(gen[5585])
		); 

/******************* CELL 5586 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5586 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5490]),
			.N(gen[5491]),
			.NE(gen[5492]),

			.O(gen[5585]),
			.E(gen[5587]),

			.SO(gen[5680]),
			.S(gen[5681]),
			.SE(gen[5682]),

			.SELF(gen[5586]),
			.cell_state(gen[5586])
		); 

/******************* CELL 5587 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5587 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5491]),
			.N(gen[5492]),
			.NE(gen[5493]),

			.O(gen[5586]),
			.E(gen[5588]),

			.SO(gen[5681]),
			.S(gen[5682]),
			.SE(gen[5683]),

			.SELF(gen[5587]),
			.cell_state(gen[5587])
		); 

/******************* CELL 5588 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5588 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5492]),
			.N(gen[5493]),
			.NE(gen[5494]),

			.O(gen[5587]),
			.E(gen[5589]),

			.SO(gen[5682]),
			.S(gen[5683]),
			.SE(gen[5684]),

			.SELF(gen[5588]),
			.cell_state(gen[5588])
		); 

/******************* CELL 5589 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5589 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5493]),
			.N(gen[5494]),
			.NE(gen[5495]),

			.O(gen[5588]),
			.E(gen[5590]),

			.SO(gen[5683]),
			.S(gen[5684]),
			.SE(gen[5685]),

			.SELF(gen[5589]),
			.cell_state(gen[5589])
		); 

/******************* CELL 5590 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5590 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5494]),
			.N(gen[5495]),
			.NE(gen[5496]),

			.O(gen[5589]),
			.E(gen[5591]),

			.SO(gen[5684]),
			.S(gen[5685]),
			.SE(gen[5686]),

			.SELF(gen[5590]),
			.cell_state(gen[5590])
		); 

/******************* CELL 5591 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5591 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5495]),
			.N(gen[5496]),
			.NE(gen[5497]),

			.O(gen[5590]),
			.E(gen[5592]),

			.SO(gen[5685]),
			.S(gen[5686]),
			.SE(gen[5687]),

			.SELF(gen[5591]),
			.cell_state(gen[5591])
		); 

/******************* CELL 5592 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5592 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5496]),
			.N(gen[5497]),
			.NE(gen[5498]),

			.O(gen[5591]),
			.E(gen[5593]),

			.SO(gen[5686]),
			.S(gen[5687]),
			.SE(gen[5688]),

			.SELF(gen[5592]),
			.cell_state(gen[5592])
		); 

/******************* CELL 5593 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5593 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5497]),
			.N(gen[5498]),
			.NE(gen[5499]),

			.O(gen[5592]),
			.E(gen[5594]),

			.SO(gen[5687]),
			.S(gen[5688]),
			.SE(gen[5689]),

			.SELF(gen[5593]),
			.cell_state(gen[5593])
		); 

/******************* CELL 5594 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5594 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5498]),
			.N(gen[5499]),
			.NE(gen[5500]),

			.O(gen[5593]),
			.E(gen[5595]),

			.SO(gen[5688]),
			.S(gen[5689]),
			.SE(gen[5690]),

			.SELF(gen[5594]),
			.cell_state(gen[5594])
		); 

/******************* CELL 5595 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5595 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5499]),
			.N(gen[5500]),
			.NE(gen[5501]),

			.O(gen[5594]),
			.E(gen[5596]),

			.SO(gen[5689]),
			.S(gen[5690]),
			.SE(gen[5691]),

			.SELF(gen[5595]),
			.cell_state(gen[5595])
		); 

/******************* CELL 5596 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5596 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5500]),
			.N(gen[5501]),
			.NE(gen[5502]),

			.O(gen[5595]),
			.E(gen[5597]),

			.SO(gen[5690]),
			.S(gen[5691]),
			.SE(gen[5692]),

			.SELF(gen[5596]),
			.cell_state(gen[5596])
		); 

/******************* CELL 5597 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5597 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5501]),
			.N(gen[5502]),
			.NE(gen[5503]),

			.O(gen[5596]),
			.E(gen[5598]),

			.SO(gen[5691]),
			.S(gen[5692]),
			.SE(gen[5693]),

			.SELF(gen[5597]),
			.cell_state(gen[5597])
		); 

/******************* CELL 5598 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5598 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5502]),
			.N(gen[5503]),
			.NE(gen[5504]),

			.O(gen[5597]),
			.E(gen[5599]),

			.SO(gen[5692]),
			.S(gen[5693]),
			.SE(gen[5694]),

			.SELF(gen[5598]),
			.cell_state(gen[5598])
		); 

/******************* CELL 5599 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5599 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5503]),
			.N(gen[5504]),
			.NE(gen[5505]),

			.O(gen[5598]),
			.E(gen[5600]),

			.SO(gen[5693]),
			.S(gen[5694]),
			.SE(gen[5695]),

			.SELF(gen[5599]),
			.cell_state(gen[5599])
		); 

/******************* CELL 5600 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5600 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5504]),
			.N(gen[5505]),
			.NE(gen[5506]),

			.O(gen[5599]),
			.E(gen[5601]),

			.SO(gen[5694]),
			.S(gen[5695]),
			.SE(gen[5696]),

			.SELF(gen[5600]),
			.cell_state(gen[5600])
		); 

/******************* CELL 5601 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5601 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5505]),
			.N(gen[5506]),
			.NE(gen[5507]),

			.O(gen[5600]),
			.E(gen[5602]),

			.SO(gen[5695]),
			.S(gen[5696]),
			.SE(gen[5697]),

			.SELF(gen[5601]),
			.cell_state(gen[5601])
		); 

/******************* CELL 5602 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5602 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5506]),
			.N(gen[5507]),
			.NE(gen[5508]),

			.O(gen[5601]),
			.E(gen[5603]),

			.SO(gen[5696]),
			.S(gen[5697]),
			.SE(gen[5698]),

			.SELF(gen[5602]),
			.cell_state(gen[5602])
		); 

/******************* CELL 5603 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5603 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5507]),
			.N(gen[5508]),
			.NE(gen[5509]),

			.O(gen[5602]),
			.E(gen[5604]),

			.SO(gen[5697]),
			.S(gen[5698]),
			.SE(gen[5699]),

			.SELF(gen[5603]),
			.cell_state(gen[5603])
		); 

/******************* CELL 5604 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5604 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5508]),
			.N(gen[5509]),
			.NE(gen[5508]),

			.O(gen[5603]),
			.E(gen[5603]),

			.SO(gen[5698]),
			.S(gen[5699]),
			.SE(gen[5698]),

			.SELF(gen[5604]),
			.cell_state(gen[5604])
		); 

/******************* CELL 5605 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5605 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5511]),
			.N(gen[5510]),
			.NE(gen[5511]),

			.O(gen[5606]),
			.E(gen[5606]),

			.SO(gen[5701]),
			.S(gen[5700]),
			.SE(gen[5701]),

			.SELF(gen[5605]),
			.cell_state(gen[5605])
		); 

/******************* CELL 5606 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5606 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5510]),
			.N(gen[5511]),
			.NE(gen[5512]),

			.O(gen[5605]),
			.E(gen[5607]),

			.SO(gen[5700]),
			.S(gen[5701]),
			.SE(gen[5702]),

			.SELF(gen[5606]),
			.cell_state(gen[5606])
		); 

/******************* CELL 5607 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5607 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5511]),
			.N(gen[5512]),
			.NE(gen[5513]),

			.O(gen[5606]),
			.E(gen[5608]),

			.SO(gen[5701]),
			.S(gen[5702]),
			.SE(gen[5703]),

			.SELF(gen[5607]),
			.cell_state(gen[5607])
		); 

/******************* CELL 5608 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5608 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5512]),
			.N(gen[5513]),
			.NE(gen[5514]),

			.O(gen[5607]),
			.E(gen[5609]),

			.SO(gen[5702]),
			.S(gen[5703]),
			.SE(gen[5704]),

			.SELF(gen[5608]),
			.cell_state(gen[5608])
		); 

/******************* CELL 5609 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5609 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5513]),
			.N(gen[5514]),
			.NE(gen[5515]),

			.O(gen[5608]),
			.E(gen[5610]),

			.SO(gen[5703]),
			.S(gen[5704]),
			.SE(gen[5705]),

			.SELF(gen[5609]),
			.cell_state(gen[5609])
		); 

/******************* CELL 5610 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5610 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5514]),
			.N(gen[5515]),
			.NE(gen[5516]),

			.O(gen[5609]),
			.E(gen[5611]),

			.SO(gen[5704]),
			.S(gen[5705]),
			.SE(gen[5706]),

			.SELF(gen[5610]),
			.cell_state(gen[5610])
		); 

/******************* CELL 5611 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5611 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5515]),
			.N(gen[5516]),
			.NE(gen[5517]),

			.O(gen[5610]),
			.E(gen[5612]),

			.SO(gen[5705]),
			.S(gen[5706]),
			.SE(gen[5707]),

			.SELF(gen[5611]),
			.cell_state(gen[5611])
		); 

/******************* CELL 5612 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5612 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5516]),
			.N(gen[5517]),
			.NE(gen[5518]),

			.O(gen[5611]),
			.E(gen[5613]),

			.SO(gen[5706]),
			.S(gen[5707]),
			.SE(gen[5708]),

			.SELF(gen[5612]),
			.cell_state(gen[5612])
		); 

/******************* CELL 5613 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5613 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5517]),
			.N(gen[5518]),
			.NE(gen[5519]),

			.O(gen[5612]),
			.E(gen[5614]),

			.SO(gen[5707]),
			.S(gen[5708]),
			.SE(gen[5709]),

			.SELF(gen[5613]),
			.cell_state(gen[5613])
		); 

/******************* CELL 5614 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5614 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5518]),
			.N(gen[5519]),
			.NE(gen[5520]),

			.O(gen[5613]),
			.E(gen[5615]),

			.SO(gen[5708]),
			.S(gen[5709]),
			.SE(gen[5710]),

			.SELF(gen[5614]),
			.cell_state(gen[5614])
		); 

/******************* CELL 5615 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5615 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5519]),
			.N(gen[5520]),
			.NE(gen[5521]),

			.O(gen[5614]),
			.E(gen[5616]),

			.SO(gen[5709]),
			.S(gen[5710]),
			.SE(gen[5711]),

			.SELF(gen[5615]),
			.cell_state(gen[5615])
		); 

/******************* CELL 5616 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5616 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5520]),
			.N(gen[5521]),
			.NE(gen[5522]),

			.O(gen[5615]),
			.E(gen[5617]),

			.SO(gen[5710]),
			.S(gen[5711]),
			.SE(gen[5712]),

			.SELF(gen[5616]),
			.cell_state(gen[5616])
		); 

/******************* CELL 5617 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5617 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5521]),
			.N(gen[5522]),
			.NE(gen[5523]),

			.O(gen[5616]),
			.E(gen[5618]),

			.SO(gen[5711]),
			.S(gen[5712]),
			.SE(gen[5713]),

			.SELF(gen[5617]),
			.cell_state(gen[5617])
		); 

/******************* CELL 5618 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5618 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5522]),
			.N(gen[5523]),
			.NE(gen[5524]),

			.O(gen[5617]),
			.E(gen[5619]),

			.SO(gen[5712]),
			.S(gen[5713]),
			.SE(gen[5714]),

			.SELF(gen[5618]),
			.cell_state(gen[5618])
		); 

/******************* CELL 5619 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5619 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5523]),
			.N(gen[5524]),
			.NE(gen[5525]),

			.O(gen[5618]),
			.E(gen[5620]),

			.SO(gen[5713]),
			.S(gen[5714]),
			.SE(gen[5715]),

			.SELF(gen[5619]),
			.cell_state(gen[5619])
		); 

/******************* CELL 5620 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5620 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5524]),
			.N(gen[5525]),
			.NE(gen[5526]),

			.O(gen[5619]),
			.E(gen[5621]),

			.SO(gen[5714]),
			.S(gen[5715]),
			.SE(gen[5716]),

			.SELF(gen[5620]),
			.cell_state(gen[5620])
		); 

/******************* CELL 5621 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5621 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5525]),
			.N(gen[5526]),
			.NE(gen[5527]),

			.O(gen[5620]),
			.E(gen[5622]),

			.SO(gen[5715]),
			.S(gen[5716]),
			.SE(gen[5717]),

			.SELF(gen[5621]),
			.cell_state(gen[5621])
		); 

/******************* CELL 5622 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5622 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5526]),
			.N(gen[5527]),
			.NE(gen[5528]),

			.O(gen[5621]),
			.E(gen[5623]),

			.SO(gen[5716]),
			.S(gen[5717]),
			.SE(gen[5718]),

			.SELF(gen[5622]),
			.cell_state(gen[5622])
		); 

/******************* CELL 5623 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5623 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5527]),
			.N(gen[5528]),
			.NE(gen[5529]),

			.O(gen[5622]),
			.E(gen[5624]),

			.SO(gen[5717]),
			.S(gen[5718]),
			.SE(gen[5719]),

			.SELF(gen[5623]),
			.cell_state(gen[5623])
		); 

/******************* CELL 5624 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5624 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5528]),
			.N(gen[5529]),
			.NE(gen[5530]),

			.O(gen[5623]),
			.E(gen[5625]),

			.SO(gen[5718]),
			.S(gen[5719]),
			.SE(gen[5720]),

			.SELF(gen[5624]),
			.cell_state(gen[5624])
		); 

/******************* CELL 5625 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5625 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5529]),
			.N(gen[5530]),
			.NE(gen[5531]),

			.O(gen[5624]),
			.E(gen[5626]),

			.SO(gen[5719]),
			.S(gen[5720]),
			.SE(gen[5721]),

			.SELF(gen[5625]),
			.cell_state(gen[5625])
		); 

/******************* CELL 5626 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5626 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5530]),
			.N(gen[5531]),
			.NE(gen[5532]),

			.O(gen[5625]),
			.E(gen[5627]),

			.SO(gen[5720]),
			.S(gen[5721]),
			.SE(gen[5722]),

			.SELF(gen[5626]),
			.cell_state(gen[5626])
		); 

/******************* CELL 5627 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5627 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5531]),
			.N(gen[5532]),
			.NE(gen[5533]),

			.O(gen[5626]),
			.E(gen[5628]),

			.SO(gen[5721]),
			.S(gen[5722]),
			.SE(gen[5723]),

			.SELF(gen[5627]),
			.cell_state(gen[5627])
		); 

/******************* CELL 5628 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5628 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5532]),
			.N(gen[5533]),
			.NE(gen[5534]),

			.O(gen[5627]),
			.E(gen[5629]),

			.SO(gen[5722]),
			.S(gen[5723]),
			.SE(gen[5724]),

			.SELF(gen[5628]),
			.cell_state(gen[5628])
		); 

/******************* CELL 5629 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5629 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5533]),
			.N(gen[5534]),
			.NE(gen[5535]),

			.O(gen[5628]),
			.E(gen[5630]),

			.SO(gen[5723]),
			.S(gen[5724]),
			.SE(gen[5725]),

			.SELF(gen[5629]),
			.cell_state(gen[5629])
		); 

/******************* CELL 5630 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5630 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5534]),
			.N(gen[5535]),
			.NE(gen[5536]),

			.O(gen[5629]),
			.E(gen[5631]),

			.SO(gen[5724]),
			.S(gen[5725]),
			.SE(gen[5726]),

			.SELF(gen[5630]),
			.cell_state(gen[5630])
		); 

/******************* CELL 5631 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5631 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5535]),
			.N(gen[5536]),
			.NE(gen[5537]),

			.O(gen[5630]),
			.E(gen[5632]),

			.SO(gen[5725]),
			.S(gen[5726]),
			.SE(gen[5727]),

			.SELF(gen[5631]),
			.cell_state(gen[5631])
		); 

/******************* CELL 5632 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5632 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5536]),
			.N(gen[5537]),
			.NE(gen[5538]),

			.O(gen[5631]),
			.E(gen[5633]),

			.SO(gen[5726]),
			.S(gen[5727]),
			.SE(gen[5728]),

			.SELF(gen[5632]),
			.cell_state(gen[5632])
		); 

/******************* CELL 5633 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5633 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5537]),
			.N(gen[5538]),
			.NE(gen[5539]),

			.O(gen[5632]),
			.E(gen[5634]),

			.SO(gen[5727]),
			.S(gen[5728]),
			.SE(gen[5729]),

			.SELF(gen[5633]),
			.cell_state(gen[5633])
		); 

/******************* CELL 5634 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5634 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5538]),
			.N(gen[5539]),
			.NE(gen[5540]),

			.O(gen[5633]),
			.E(gen[5635]),

			.SO(gen[5728]),
			.S(gen[5729]),
			.SE(gen[5730]),

			.SELF(gen[5634]),
			.cell_state(gen[5634])
		); 

/******************* CELL 5635 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5635 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5539]),
			.N(gen[5540]),
			.NE(gen[5541]),

			.O(gen[5634]),
			.E(gen[5636]),

			.SO(gen[5729]),
			.S(gen[5730]),
			.SE(gen[5731]),

			.SELF(gen[5635]),
			.cell_state(gen[5635])
		); 

/******************* CELL 5636 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5636 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5540]),
			.N(gen[5541]),
			.NE(gen[5542]),

			.O(gen[5635]),
			.E(gen[5637]),

			.SO(gen[5730]),
			.S(gen[5731]),
			.SE(gen[5732]),

			.SELF(gen[5636]),
			.cell_state(gen[5636])
		); 

/******************* CELL 5637 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5637 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5541]),
			.N(gen[5542]),
			.NE(gen[5543]),

			.O(gen[5636]),
			.E(gen[5638]),

			.SO(gen[5731]),
			.S(gen[5732]),
			.SE(gen[5733]),

			.SELF(gen[5637]),
			.cell_state(gen[5637])
		); 

/******************* CELL 5638 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5638 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5542]),
			.N(gen[5543]),
			.NE(gen[5544]),

			.O(gen[5637]),
			.E(gen[5639]),

			.SO(gen[5732]),
			.S(gen[5733]),
			.SE(gen[5734]),

			.SELF(gen[5638]),
			.cell_state(gen[5638])
		); 

/******************* CELL 5639 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5639 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5543]),
			.N(gen[5544]),
			.NE(gen[5545]),

			.O(gen[5638]),
			.E(gen[5640]),

			.SO(gen[5733]),
			.S(gen[5734]),
			.SE(gen[5735]),

			.SELF(gen[5639]),
			.cell_state(gen[5639])
		); 

/******************* CELL 5640 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5640 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5544]),
			.N(gen[5545]),
			.NE(gen[5546]),

			.O(gen[5639]),
			.E(gen[5641]),

			.SO(gen[5734]),
			.S(gen[5735]),
			.SE(gen[5736]),

			.SELF(gen[5640]),
			.cell_state(gen[5640])
		); 

/******************* CELL 5641 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5641 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5545]),
			.N(gen[5546]),
			.NE(gen[5547]),

			.O(gen[5640]),
			.E(gen[5642]),

			.SO(gen[5735]),
			.S(gen[5736]),
			.SE(gen[5737]),

			.SELF(gen[5641]),
			.cell_state(gen[5641])
		); 

/******************* CELL 5642 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5642 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5546]),
			.N(gen[5547]),
			.NE(gen[5548]),

			.O(gen[5641]),
			.E(gen[5643]),

			.SO(gen[5736]),
			.S(gen[5737]),
			.SE(gen[5738]),

			.SELF(gen[5642]),
			.cell_state(gen[5642])
		); 

/******************* CELL 5643 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5643 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5547]),
			.N(gen[5548]),
			.NE(gen[5549]),

			.O(gen[5642]),
			.E(gen[5644]),

			.SO(gen[5737]),
			.S(gen[5738]),
			.SE(gen[5739]),

			.SELF(gen[5643]),
			.cell_state(gen[5643])
		); 

/******************* CELL 5644 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5644 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5548]),
			.N(gen[5549]),
			.NE(gen[5550]),

			.O(gen[5643]),
			.E(gen[5645]),

			.SO(gen[5738]),
			.S(gen[5739]),
			.SE(gen[5740]),

			.SELF(gen[5644]),
			.cell_state(gen[5644])
		); 

/******************* CELL 5645 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5645 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5549]),
			.N(gen[5550]),
			.NE(gen[5551]),

			.O(gen[5644]),
			.E(gen[5646]),

			.SO(gen[5739]),
			.S(gen[5740]),
			.SE(gen[5741]),

			.SELF(gen[5645]),
			.cell_state(gen[5645])
		); 

/******************* CELL 5646 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5646 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5550]),
			.N(gen[5551]),
			.NE(gen[5552]),

			.O(gen[5645]),
			.E(gen[5647]),

			.SO(gen[5740]),
			.S(gen[5741]),
			.SE(gen[5742]),

			.SELF(gen[5646]),
			.cell_state(gen[5646])
		); 

/******************* CELL 5647 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5647 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5551]),
			.N(gen[5552]),
			.NE(gen[5553]),

			.O(gen[5646]),
			.E(gen[5648]),

			.SO(gen[5741]),
			.S(gen[5742]),
			.SE(gen[5743]),

			.SELF(gen[5647]),
			.cell_state(gen[5647])
		); 

/******************* CELL 5648 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5648 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5552]),
			.N(gen[5553]),
			.NE(gen[5554]),

			.O(gen[5647]),
			.E(gen[5649]),

			.SO(gen[5742]),
			.S(gen[5743]),
			.SE(gen[5744]),

			.SELF(gen[5648]),
			.cell_state(gen[5648])
		); 

/******************* CELL 5649 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5649 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5553]),
			.N(gen[5554]),
			.NE(gen[5555]),

			.O(gen[5648]),
			.E(gen[5650]),

			.SO(gen[5743]),
			.S(gen[5744]),
			.SE(gen[5745]),

			.SELF(gen[5649]),
			.cell_state(gen[5649])
		); 

/******************* CELL 5650 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5650 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5554]),
			.N(gen[5555]),
			.NE(gen[5556]),

			.O(gen[5649]),
			.E(gen[5651]),

			.SO(gen[5744]),
			.S(gen[5745]),
			.SE(gen[5746]),

			.SELF(gen[5650]),
			.cell_state(gen[5650])
		); 

/******************* CELL 5651 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5651 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5555]),
			.N(gen[5556]),
			.NE(gen[5557]),

			.O(gen[5650]),
			.E(gen[5652]),

			.SO(gen[5745]),
			.S(gen[5746]),
			.SE(gen[5747]),

			.SELF(gen[5651]),
			.cell_state(gen[5651])
		); 

/******************* CELL 5652 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5652 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5556]),
			.N(gen[5557]),
			.NE(gen[5558]),

			.O(gen[5651]),
			.E(gen[5653]),

			.SO(gen[5746]),
			.S(gen[5747]),
			.SE(gen[5748]),

			.SELF(gen[5652]),
			.cell_state(gen[5652])
		); 

/******************* CELL 5653 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5653 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5557]),
			.N(gen[5558]),
			.NE(gen[5559]),

			.O(gen[5652]),
			.E(gen[5654]),

			.SO(gen[5747]),
			.S(gen[5748]),
			.SE(gen[5749]),

			.SELF(gen[5653]),
			.cell_state(gen[5653])
		); 

/******************* CELL 5654 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5654 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5558]),
			.N(gen[5559]),
			.NE(gen[5560]),

			.O(gen[5653]),
			.E(gen[5655]),

			.SO(gen[5748]),
			.S(gen[5749]),
			.SE(gen[5750]),

			.SELF(gen[5654]),
			.cell_state(gen[5654])
		); 

/******************* CELL 5655 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5655 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5559]),
			.N(gen[5560]),
			.NE(gen[5561]),

			.O(gen[5654]),
			.E(gen[5656]),

			.SO(gen[5749]),
			.S(gen[5750]),
			.SE(gen[5751]),

			.SELF(gen[5655]),
			.cell_state(gen[5655])
		); 

/******************* CELL 5656 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5656 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5560]),
			.N(gen[5561]),
			.NE(gen[5562]),

			.O(gen[5655]),
			.E(gen[5657]),

			.SO(gen[5750]),
			.S(gen[5751]),
			.SE(gen[5752]),

			.SELF(gen[5656]),
			.cell_state(gen[5656])
		); 

/******************* CELL 5657 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5657 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5561]),
			.N(gen[5562]),
			.NE(gen[5563]),

			.O(gen[5656]),
			.E(gen[5658]),

			.SO(gen[5751]),
			.S(gen[5752]),
			.SE(gen[5753]),

			.SELF(gen[5657]),
			.cell_state(gen[5657])
		); 

/******************* CELL 5658 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5658 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5562]),
			.N(gen[5563]),
			.NE(gen[5564]),

			.O(gen[5657]),
			.E(gen[5659]),

			.SO(gen[5752]),
			.S(gen[5753]),
			.SE(gen[5754]),

			.SELF(gen[5658]),
			.cell_state(gen[5658])
		); 

/******************* CELL 5659 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5659 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5563]),
			.N(gen[5564]),
			.NE(gen[5565]),

			.O(gen[5658]),
			.E(gen[5660]),

			.SO(gen[5753]),
			.S(gen[5754]),
			.SE(gen[5755]),

			.SELF(gen[5659]),
			.cell_state(gen[5659])
		); 

/******************* CELL 5660 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5660 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5564]),
			.N(gen[5565]),
			.NE(gen[5566]),

			.O(gen[5659]),
			.E(gen[5661]),

			.SO(gen[5754]),
			.S(gen[5755]),
			.SE(gen[5756]),

			.SELF(gen[5660]),
			.cell_state(gen[5660])
		); 

/******************* CELL 5661 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5661 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5565]),
			.N(gen[5566]),
			.NE(gen[5567]),

			.O(gen[5660]),
			.E(gen[5662]),

			.SO(gen[5755]),
			.S(gen[5756]),
			.SE(gen[5757]),

			.SELF(gen[5661]),
			.cell_state(gen[5661])
		); 

/******************* CELL 5662 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5662 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5566]),
			.N(gen[5567]),
			.NE(gen[5568]),

			.O(gen[5661]),
			.E(gen[5663]),

			.SO(gen[5756]),
			.S(gen[5757]),
			.SE(gen[5758]),

			.SELF(gen[5662]),
			.cell_state(gen[5662])
		); 

/******************* CELL 5663 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5663 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5567]),
			.N(gen[5568]),
			.NE(gen[5569]),

			.O(gen[5662]),
			.E(gen[5664]),

			.SO(gen[5757]),
			.S(gen[5758]),
			.SE(gen[5759]),

			.SELF(gen[5663]),
			.cell_state(gen[5663])
		); 

/******************* CELL 5664 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5664 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5568]),
			.N(gen[5569]),
			.NE(gen[5570]),

			.O(gen[5663]),
			.E(gen[5665]),

			.SO(gen[5758]),
			.S(gen[5759]),
			.SE(gen[5760]),

			.SELF(gen[5664]),
			.cell_state(gen[5664])
		); 

/******************* CELL 5665 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5665 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5569]),
			.N(gen[5570]),
			.NE(gen[5571]),

			.O(gen[5664]),
			.E(gen[5666]),

			.SO(gen[5759]),
			.S(gen[5760]),
			.SE(gen[5761]),

			.SELF(gen[5665]),
			.cell_state(gen[5665])
		); 

/******************* CELL 5666 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5666 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5570]),
			.N(gen[5571]),
			.NE(gen[5572]),

			.O(gen[5665]),
			.E(gen[5667]),

			.SO(gen[5760]),
			.S(gen[5761]),
			.SE(gen[5762]),

			.SELF(gen[5666]),
			.cell_state(gen[5666])
		); 

/******************* CELL 5667 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5667 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5571]),
			.N(gen[5572]),
			.NE(gen[5573]),

			.O(gen[5666]),
			.E(gen[5668]),

			.SO(gen[5761]),
			.S(gen[5762]),
			.SE(gen[5763]),

			.SELF(gen[5667]),
			.cell_state(gen[5667])
		); 

/******************* CELL 5668 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5668 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5572]),
			.N(gen[5573]),
			.NE(gen[5574]),

			.O(gen[5667]),
			.E(gen[5669]),

			.SO(gen[5762]),
			.S(gen[5763]),
			.SE(gen[5764]),

			.SELF(gen[5668]),
			.cell_state(gen[5668])
		); 

/******************* CELL 5669 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5669 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5573]),
			.N(gen[5574]),
			.NE(gen[5575]),

			.O(gen[5668]),
			.E(gen[5670]),

			.SO(gen[5763]),
			.S(gen[5764]),
			.SE(gen[5765]),

			.SELF(gen[5669]),
			.cell_state(gen[5669])
		); 

/******************* CELL 5670 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5670 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5574]),
			.N(gen[5575]),
			.NE(gen[5576]),

			.O(gen[5669]),
			.E(gen[5671]),

			.SO(gen[5764]),
			.S(gen[5765]),
			.SE(gen[5766]),

			.SELF(gen[5670]),
			.cell_state(gen[5670])
		); 

/******************* CELL 5671 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5671 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5575]),
			.N(gen[5576]),
			.NE(gen[5577]),

			.O(gen[5670]),
			.E(gen[5672]),

			.SO(gen[5765]),
			.S(gen[5766]),
			.SE(gen[5767]),

			.SELF(gen[5671]),
			.cell_state(gen[5671])
		); 

/******************* CELL 5672 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5672 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5576]),
			.N(gen[5577]),
			.NE(gen[5578]),

			.O(gen[5671]),
			.E(gen[5673]),

			.SO(gen[5766]),
			.S(gen[5767]),
			.SE(gen[5768]),

			.SELF(gen[5672]),
			.cell_state(gen[5672])
		); 

/******************* CELL 5673 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5673 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5577]),
			.N(gen[5578]),
			.NE(gen[5579]),

			.O(gen[5672]),
			.E(gen[5674]),

			.SO(gen[5767]),
			.S(gen[5768]),
			.SE(gen[5769]),

			.SELF(gen[5673]),
			.cell_state(gen[5673])
		); 

/******************* CELL 5674 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5674 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5578]),
			.N(gen[5579]),
			.NE(gen[5580]),

			.O(gen[5673]),
			.E(gen[5675]),

			.SO(gen[5768]),
			.S(gen[5769]),
			.SE(gen[5770]),

			.SELF(gen[5674]),
			.cell_state(gen[5674])
		); 

/******************* CELL 5675 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5675 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5579]),
			.N(gen[5580]),
			.NE(gen[5581]),

			.O(gen[5674]),
			.E(gen[5676]),

			.SO(gen[5769]),
			.S(gen[5770]),
			.SE(gen[5771]),

			.SELF(gen[5675]),
			.cell_state(gen[5675])
		); 

/******************* CELL 5676 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5676 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5580]),
			.N(gen[5581]),
			.NE(gen[5582]),

			.O(gen[5675]),
			.E(gen[5677]),

			.SO(gen[5770]),
			.S(gen[5771]),
			.SE(gen[5772]),

			.SELF(gen[5676]),
			.cell_state(gen[5676])
		); 

/******************* CELL 5677 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5677 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5581]),
			.N(gen[5582]),
			.NE(gen[5583]),

			.O(gen[5676]),
			.E(gen[5678]),

			.SO(gen[5771]),
			.S(gen[5772]),
			.SE(gen[5773]),

			.SELF(gen[5677]),
			.cell_state(gen[5677])
		); 

/******************* CELL 5678 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5678 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5582]),
			.N(gen[5583]),
			.NE(gen[5584]),

			.O(gen[5677]),
			.E(gen[5679]),

			.SO(gen[5772]),
			.S(gen[5773]),
			.SE(gen[5774]),

			.SELF(gen[5678]),
			.cell_state(gen[5678])
		); 

/******************* CELL 5679 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5679 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5583]),
			.N(gen[5584]),
			.NE(gen[5585]),

			.O(gen[5678]),
			.E(gen[5680]),

			.SO(gen[5773]),
			.S(gen[5774]),
			.SE(gen[5775]),

			.SELF(gen[5679]),
			.cell_state(gen[5679])
		); 

/******************* CELL 5680 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5680 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5584]),
			.N(gen[5585]),
			.NE(gen[5586]),

			.O(gen[5679]),
			.E(gen[5681]),

			.SO(gen[5774]),
			.S(gen[5775]),
			.SE(gen[5776]),

			.SELF(gen[5680]),
			.cell_state(gen[5680])
		); 

/******************* CELL 5681 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5681 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5585]),
			.N(gen[5586]),
			.NE(gen[5587]),

			.O(gen[5680]),
			.E(gen[5682]),

			.SO(gen[5775]),
			.S(gen[5776]),
			.SE(gen[5777]),

			.SELF(gen[5681]),
			.cell_state(gen[5681])
		); 

/******************* CELL 5682 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5682 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5586]),
			.N(gen[5587]),
			.NE(gen[5588]),

			.O(gen[5681]),
			.E(gen[5683]),

			.SO(gen[5776]),
			.S(gen[5777]),
			.SE(gen[5778]),

			.SELF(gen[5682]),
			.cell_state(gen[5682])
		); 

/******************* CELL 5683 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5683 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5587]),
			.N(gen[5588]),
			.NE(gen[5589]),

			.O(gen[5682]),
			.E(gen[5684]),

			.SO(gen[5777]),
			.S(gen[5778]),
			.SE(gen[5779]),

			.SELF(gen[5683]),
			.cell_state(gen[5683])
		); 

/******************* CELL 5684 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5684 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5588]),
			.N(gen[5589]),
			.NE(gen[5590]),

			.O(gen[5683]),
			.E(gen[5685]),

			.SO(gen[5778]),
			.S(gen[5779]),
			.SE(gen[5780]),

			.SELF(gen[5684]),
			.cell_state(gen[5684])
		); 

/******************* CELL 5685 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5685 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5589]),
			.N(gen[5590]),
			.NE(gen[5591]),

			.O(gen[5684]),
			.E(gen[5686]),

			.SO(gen[5779]),
			.S(gen[5780]),
			.SE(gen[5781]),

			.SELF(gen[5685]),
			.cell_state(gen[5685])
		); 

/******************* CELL 5686 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5686 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5590]),
			.N(gen[5591]),
			.NE(gen[5592]),

			.O(gen[5685]),
			.E(gen[5687]),

			.SO(gen[5780]),
			.S(gen[5781]),
			.SE(gen[5782]),

			.SELF(gen[5686]),
			.cell_state(gen[5686])
		); 

/******************* CELL 5687 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5687 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5591]),
			.N(gen[5592]),
			.NE(gen[5593]),

			.O(gen[5686]),
			.E(gen[5688]),

			.SO(gen[5781]),
			.S(gen[5782]),
			.SE(gen[5783]),

			.SELF(gen[5687]),
			.cell_state(gen[5687])
		); 

/******************* CELL 5688 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5688 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5592]),
			.N(gen[5593]),
			.NE(gen[5594]),

			.O(gen[5687]),
			.E(gen[5689]),

			.SO(gen[5782]),
			.S(gen[5783]),
			.SE(gen[5784]),

			.SELF(gen[5688]),
			.cell_state(gen[5688])
		); 

/******************* CELL 5689 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5689 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5593]),
			.N(gen[5594]),
			.NE(gen[5595]),

			.O(gen[5688]),
			.E(gen[5690]),

			.SO(gen[5783]),
			.S(gen[5784]),
			.SE(gen[5785]),

			.SELF(gen[5689]),
			.cell_state(gen[5689])
		); 

/******************* CELL 5690 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5690 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5594]),
			.N(gen[5595]),
			.NE(gen[5596]),

			.O(gen[5689]),
			.E(gen[5691]),

			.SO(gen[5784]),
			.S(gen[5785]),
			.SE(gen[5786]),

			.SELF(gen[5690]),
			.cell_state(gen[5690])
		); 

/******************* CELL 5691 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5691 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5595]),
			.N(gen[5596]),
			.NE(gen[5597]),

			.O(gen[5690]),
			.E(gen[5692]),

			.SO(gen[5785]),
			.S(gen[5786]),
			.SE(gen[5787]),

			.SELF(gen[5691]),
			.cell_state(gen[5691])
		); 

/******************* CELL 5692 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5692 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5596]),
			.N(gen[5597]),
			.NE(gen[5598]),

			.O(gen[5691]),
			.E(gen[5693]),

			.SO(gen[5786]),
			.S(gen[5787]),
			.SE(gen[5788]),

			.SELF(gen[5692]),
			.cell_state(gen[5692])
		); 

/******************* CELL 5693 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5693 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5597]),
			.N(gen[5598]),
			.NE(gen[5599]),

			.O(gen[5692]),
			.E(gen[5694]),

			.SO(gen[5787]),
			.S(gen[5788]),
			.SE(gen[5789]),

			.SELF(gen[5693]),
			.cell_state(gen[5693])
		); 

/******************* CELL 5694 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5694 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5598]),
			.N(gen[5599]),
			.NE(gen[5600]),

			.O(gen[5693]),
			.E(gen[5695]),

			.SO(gen[5788]),
			.S(gen[5789]),
			.SE(gen[5790]),

			.SELF(gen[5694]),
			.cell_state(gen[5694])
		); 

/******************* CELL 5695 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5695 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5599]),
			.N(gen[5600]),
			.NE(gen[5601]),

			.O(gen[5694]),
			.E(gen[5696]),

			.SO(gen[5789]),
			.S(gen[5790]),
			.SE(gen[5791]),

			.SELF(gen[5695]),
			.cell_state(gen[5695])
		); 

/******************* CELL 5696 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5696 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5600]),
			.N(gen[5601]),
			.NE(gen[5602]),

			.O(gen[5695]),
			.E(gen[5697]),

			.SO(gen[5790]),
			.S(gen[5791]),
			.SE(gen[5792]),

			.SELF(gen[5696]),
			.cell_state(gen[5696])
		); 

/******************* CELL 5697 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5697 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5601]),
			.N(gen[5602]),
			.NE(gen[5603]),

			.O(gen[5696]),
			.E(gen[5698]),

			.SO(gen[5791]),
			.S(gen[5792]),
			.SE(gen[5793]),

			.SELF(gen[5697]),
			.cell_state(gen[5697])
		); 

/******************* CELL 5698 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5698 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5602]),
			.N(gen[5603]),
			.NE(gen[5604]),

			.O(gen[5697]),
			.E(gen[5699]),

			.SO(gen[5792]),
			.S(gen[5793]),
			.SE(gen[5794]),

			.SELF(gen[5698]),
			.cell_state(gen[5698])
		); 

/******************* CELL 5699 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5699 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5603]),
			.N(gen[5604]),
			.NE(gen[5603]),

			.O(gen[5698]),
			.E(gen[5698]),

			.SO(gen[5793]),
			.S(gen[5794]),
			.SE(gen[5793]),

			.SELF(gen[5699]),
			.cell_state(gen[5699])
		); 

/******************* CELL 5700 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5700 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5606]),
			.N(gen[5605]),
			.NE(gen[5606]),

			.O(gen[5701]),
			.E(gen[5701]),

			.SO(gen[5796]),
			.S(gen[5795]),
			.SE(gen[5796]),

			.SELF(gen[5700]),
			.cell_state(gen[5700])
		); 

/******************* CELL 5701 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5701 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5605]),
			.N(gen[5606]),
			.NE(gen[5607]),

			.O(gen[5700]),
			.E(gen[5702]),

			.SO(gen[5795]),
			.S(gen[5796]),
			.SE(gen[5797]),

			.SELF(gen[5701]),
			.cell_state(gen[5701])
		); 

/******************* CELL 5702 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5702 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5606]),
			.N(gen[5607]),
			.NE(gen[5608]),

			.O(gen[5701]),
			.E(gen[5703]),

			.SO(gen[5796]),
			.S(gen[5797]),
			.SE(gen[5798]),

			.SELF(gen[5702]),
			.cell_state(gen[5702])
		); 

/******************* CELL 5703 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5703 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5607]),
			.N(gen[5608]),
			.NE(gen[5609]),

			.O(gen[5702]),
			.E(gen[5704]),

			.SO(gen[5797]),
			.S(gen[5798]),
			.SE(gen[5799]),

			.SELF(gen[5703]),
			.cell_state(gen[5703])
		); 

/******************* CELL 5704 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5704 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5608]),
			.N(gen[5609]),
			.NE(gen[5610]),

			.O(gen[5703]),
			.E(gen[5705]),

			.SO(gen[5798]),
			.S(gen[5799]),
			.SE(gen[5800]),

			.SELF(gen[5704]),
			.cell_state(gen[5704])
		); 

/******************* CELL 5705 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5705 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5609]),
			.N(gen[5610]),
			.NE(gen[5611]),

			.O(gen[5704]),
			.E(gen[5706]),

			.SO(gen[5799]),
			.S(gen[5800]),
			.SE(gen[5801]),

			.SELF(gen[5705]),
			.cell_state(gen[5705])
		); 

/******************* CELL 5706 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5706 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5610]),
			.N(gen[5611]),
			.NE(gen[5612]),

			.O(gen[5705]),
			.E(gen[5707]),

			.SO(gen[5800]),
			.S(gen[5801]),
			.SE(gen[5802]),

			.SELF(gen[5706]),
			.cell_state(gen[5706])
		); 

/******************* CELL 5707 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5707 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5611]),
			.N(gen[5612]),
			.NE(gen[5613]),

			.O(gen[5706]),
			.E(gen[5708]),

			.SO(gen[5801]),
			.S(gen[5802]),
			.SE(gen[5803]),

			.SELF(gen[5707]),
			.cell_state(gen[5707])
		); 

/******************* CELL 5708 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5708 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5612]),
			.N(gen[5613]),
			.NE(gen[5614]),

			.O(gen[5707]),
			.E(gen[5709]),

			.SO(gen[5802]),
			.S(gen[5803]),
			.SE(gen[5804]),

			.SELF(gen[5708]),
			.cell_state(gen[5708])
		); 

/******************* CELL 5709 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5709 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5613]),
			.N(gen[5614]),
			.NE(gen[5615]),

			.O(gen[5708]),
			.E(gen[5710]),

			.SO(gen[5803]),
			.S(gen[5804]),
			.SE(gen[5805]),

			.SELF(gen[5709]),
			.cell_state(gen[5709])
		); 

/******************* CELL 5710 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5710 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5614]),
			.N(gen[5615]),
			.NE(gen[5616]),

			.O(gen[5709]),
			.E(gen[5711]),

			.SO(gen[5804]),
			.S(gen[5805]),
			.SE(gen[5806]),

			.SELF(gen[5710]),
			.cell_state(gen[5710])
		); 

/******************* CELL 5711 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5711 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5615]),
			.N(gen[5616]),
			.NE(gen[5617]),

			.O(gen[5710]),
			.E(gen[5712]),

			.SO(gen[5805]),
			.S(gen[5806]),
			.SE(gen[5807]),

			.SELF(gen[5711]),
			.cell_state(gen[5711])
		); 

/******************* CELL 5712 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5712 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5616]),
			.N(gen[5617]),
			.NE(gen[5618]),

			.O(gen[5711]),
			.E(gen[5713]),

			.SO(gen[5806]),
			.S(gen[5807]),
			.SE(gen[5808]),

			.SELF(gen[5712]),
			.cell_state(gen[5712])
		); 

/******************* CELL 5713 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5713 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5617]),
			.N(gen[5618]),
			.NE(gen[5619]),

			.O(gen[5712]),
			.E(gen[5714]),

			.SO(gen[5807]),
			.S(gen[5808]),
			.SE(gen[5809]),

			.SELF(gen[5713]),
			.cell_state(gen[5713])
		); 

/******************* CELL 5714 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5714 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5618]),
			.N(gen[5619]),
			.NE(gen[5620]),

			.O(gen[5713]),
			.E(gen[5715]),

			.SO(gen[5808]),
			.S(gen[5809]),
			.SE(gen[5810]),

			.SELF(gen[5714]),
			.cell_state(gen[5714])
		); 

/******************* CELL 5715 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5715 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5619]),
			.N(gen[5620]),
			.NE(gen[5621]),

			.O(gen[5714]),
			.E(gen[5716]),

			.SO(gen[5809]),
			.S(gen[5810]),
			.SE(gen[5811]),

			.SELF(gen[5715]),
			.cell_state(gen[5715])
		); 

/******************* CELL 5716 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5716 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5620]),
			.N(gen[5621]),
			.NE(gen[5622]),

			.O(gen[5715]),
			.E(gen[5717]),

			.SO(gen[5810]),
			.S(gen[5811]),
			.SE(gen[5812]),

			.SELF(gen[5716]),
			.cell_state(gen[5716])
		); 

/******************* CELL 5717 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5717 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5621]),
			.N(gen[5622]),
			.NE(gen[5623]),

			.O(gen[5716]),
			.E(gen[5718]),

			.SO(gen[5811]),
			.S(gen[5812]),
			.SE(gen[5813]),

			.SELF(gen[5717]),
			.cell_state(gen[5717])
		); 

/******************* CELL 5718 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5718 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5622]),
			.N(gen[5623]),
			.NE(gen[5624]),

			.O(gen[5717]),
			.E(gen[5719]),

			.SO(gen[5812]),
			.S(gen[5813]),
			.SE(gen[5814]),

			.SELF(gen[5718]),
			.cell_state(gen[5718])
		); 

/******************* CELL 5719 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5719 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5623]),
			.N(gen[5624]),
			.NE(gen[5625]),

			.O(gen[5718]),
			.E(gen[5720]),

			.SO(gen[5813]),
			.S(gen[5814]),
			.SE(gen[5815]),

			.SELF(gen[5719]),
			.cell_state(gen[5719])
		); 

/******************* CELL 5720 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5720 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5624]),
			.N(gen[5625]),
			.NE(gen[5626]),

			.O(gen[5719]),
			.E(gen[5721]),

			.SO(gen[5814]),
			.S(gen[5815]),
			.SE(gen[5816]),

			.SELF(gen[5720]),
			.cell_state(gen[5720])
		); 

/******************* CELL 5721 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5721 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5625]),
			.N(gen[5626]),
			.NE(gen[5627]),

			.O(gen[5720]),
			.E(gen[5722]),

			.SO(gen[5815]),
			.S(gen[5816]),
			.SE(gen[5817]),

			.SELF(gen[5721]),
			.cell_state(gen[5721])
		); 

/******************* CELL 5722 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5722 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5626]),
			.N(gen[5627]),
			.NE(gen[5628]),

			.O(gen[5721]),
			.E(gen[5723]),

			.SO(gen[5816]),
			.S(gen[5817]),
			.SE(gen[5818]),

			.SELF(gen[5722]),
			.cell_state(gen[5722])
		); 

/******************* CELL 5723 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5723 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5627]),
			.N(gen[5628]),
			.NE(gen[5629]),

			.O(gen[5722]),
			.E(gen[5724]),

			.SO(gen[5817]),
			.S(gen[5818]),
			.SE(gen[5819]),

			.SELF(gen[5723]),
			.cell_state(gen[5723])
		); 

/******************* CELL 5724 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5724 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5628]),
			.N(gen[5629]),
			.NE(gen[5630]),

			.O(gen[5723]),
			.E(gen[5725]),

			.SO(gen[5818]),
			.S(gen[5819]),
			.SE(gen[5820]),

			.SELF(gen[5724]),
			.cell_state(gen[5724])
		); 

/******************* CELL 5725 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5725 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5629]),
			.N(gen[5630]),
			.NE(gen[5631]),

			.O(gen[5724]),
			.E(gen[5726]),

			.SO(gen[5819]),
			.S(gen[5820]),
			.SE(gen[5821]),

			.SELF(gen[5725]),
			.cell_state(gen[5725])
		); 

/******************* CELL 5726 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5726 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5630]),
			.N(gen[5631]),
			.NE(gen[5632]),

			.O(gen[5725]),
			.E(gen[5727]),

			.SO(gen[5820]),
			.S(gen[5821]),
			.SE(gen[5822]),

			.SELF(gen[5726]),
			.cell_state(gen[5726])
		); 

/******************* CELL 5727 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5727 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5631]),
			.N(gen[5632]),
			.NE(gen[5633]),

			.O(gen[5726]),
			.E(gen[5728]),

			.SO(gen[5821]),
			.S(gen[5822]),
			.SE(gen[5823]),

			.SELF(gen[5727]),
			.cell_state(gen[5727])
		); 

/******************* CELL 5728 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5728 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5632]),
			.N(gen[5633]),
			.NE(gen[5634]),

			.O(gen[5727]),
			.E(gen[5729]),

			.SO(gen[5822]),
			.S(gen[5823]),
			.SE(gen[5824]),

			.SELF(gen[5728]),
			.cell_state(gen[5728])
		); 

/******************* CELL 5729 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5729 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5633]),
			.N(gen[5634]),
			.NE(gen[5635]),

			.O(gen[5728]),
			.E(gen[5730]),

			.SO(gen[5823]),
			.S(gen[5824]),
			.SE(gen[5825]),

			.SELF(gen[5729]),
			.cell_state(gen[5729])
		); 

/******************* CELL 5730 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5730 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5634]),
			.N(gen[5635]),
			.NE(gen[5636]),

			.O(gen[5729]),
			.E(gen[5731]),

			.SO(gen[5824]),
			.S(gen[5825]),
			.SE(gen[5826]),

			.SELF(gen[5730]),
			.cell_state(gen[5730])
		); 

/******************* CELL 5731 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5731 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5635]),
			.N(gen[5636]),
			.NE(gen[5637]),

			.O(gen[5730]),
			.E(gen[5732]),

			.SO(gen[5825]),
			.S(gen[5826]),
			.SE(gen[5827]),

			.SELF(gen[5731]),
			.cell_state(gen[5731])
		); 

/******************* CELL 5732 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5732 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5636]),
			.N(gen[5637]),
			.NE(gen[5638]),

			.O(gen[5731]),
			.E(gen[5733]),

			.SO(gen[5826]),
			.S(gen[5827]),
			.SE(gen[5828]),

			.SELF(gen[5732]),
			.cell_state(gen[5732])
		); 

/******************* CELL 5733 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5733 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5637]),
			.N(gen[5638]),
			.NE(gen[5639]),

			.O(gen[5732]),
			.E(gen[5734]),

			.SO(gen[5827]),
			.S(gen[5828]),
			.SE(gen[5829]),

			.SELF(gen[5733]),
			.cell_state(gen[5733])
		); 

/******************* CELL 5734 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5734 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5638]),
			.N(gen[5639]),
			.NE(gen[5640]),

			.O(gen[5733]),
			.E(gen[5735]),

			.SO(gen[5828]),
			.S(gen[5829]),
			.SE(gen[5830]),

			.SELF(gen[5734]),
			.cell_state(gen[5734])
		); 

/******************* CELL 5735 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5735 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5639]),
			.N(gen[5640]),
			.NE(gen[5641]),

			.O(gen[5734]),
			.E(gen[5736]),

			.SO(gen[5829]),
			.S(gen[5830]),
			.SE(gen[5831]),

			.SELF(gen[5735]),
			.cell_state(gen[5735])
		); 

/******************* CELL 5736 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5736 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5640]),
			.N(gen[5641]),
			.NE(gen[5642]),

			.O(gen[5735]),
			.E(gen[5737]),

			.SO(gen[5830]),
			.S(gen[5831]),
			.SE(gen[5832]),

			.SELF(gen[5736]),
			.cell_state(gen[5736])
		); 

/******************* CELL 5737 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5737 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5641]),
			.N(gen[5642]),
			.NE(gen[5643]),

			.O(gen[5736]),
			.E(gen[5738]),

			.SO(gen[5831]),
			.S(gen[5832]),
			.SE(gen[5833]),

			.SELF(gen[5737]),
			.cell_state(gen[5737])
		); 

/******************* CELL 5738 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5738 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5642]),
			.N(gen[5643]),
			.NE(gen[5644]),

			.O(gen[5737]),
			.E(gen[5739]),

			.SO(gen[5832]),
			.S(gen[5833]),
			.SE(gen[5834]),

			.SELF(gen[5738]),
			.cell_state(gen[5738])
		); 

/******************* CELL 5739 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5739 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5643]),
			.N(gen[5644]),
			.NE(gen[5645]),

			.O(gen[5738]),
			.E(gen[5740]),

			.SO(gen[5833]),
			.S(gen[5834]),
			.SE(gen[5835]),

			.SELF(gen[5739]),
			.cell_state(gen[5739])
		); 

/******************* CELL 5740 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5740 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5644]),
			.N(gen[5645]),
			.NE(gen[5646]),

			.O(gen[5739]),
			.E(gen[5741]),

			.SO(gen[5834]),
			.S(gen[5835]),
			.SE(gen[5836]),

			.SELF(gen[5740]),
			.cell_state(gen[5740])
		); 

/******************* CELL 5741 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5741 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5645]),
			.N(gen[5646]),
			.NE(gen[5647]),

			.O(gen[5740]),
			.E(gen[5742]),

			.SO(gen[5835]),
			.S(gen[5836]),
			.SE(gen[5837]),

			.SELF(gen[5741]),
			.cell_state(gen[5741])
		); 

/******************* CELL 5742 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5742 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5646]),
			.N(gen[5647]),
			.NE(gen[5648]),

			.O(gen[5741]),
			.E(gen[5743]),

			.SO(gen[5836]),
			.S(gen[5837]),
			.SE(gen[5838]),

			.SELF(gen[5742]),
			.cell_state(gen[5742])
		); 

/******************* CELL 5743 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5743 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5647]),
			.N(gen[5648]),
			.NE(gen[5649]),

			.O(gen[5742]),
			.E(gen[5744]),

			.SO(gen[5837]),
			.S(gen[5838]),
			.SE(gen[5839]),

			.SELF(gen[5743]),
			.cell_state(gen[5743])
		); 

/******************* CELL 5744 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5744 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5648]),
			.N(gen[5649]),
			.NE(gen[5650]),

			.O(gen[5743]),
			.E(gen[5745]),

			.SO(gen[5838]),
			.S(gen[5839]),
			.SE(gen[5840]),

			.SELF(gen[5744]),
			.cell_state(gen[5744])
		); 

/******************* CELL 5745 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5745 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5649]),
			.N(gen[5650]),
			.NE(gen[5651]),

			.O(gen[5744]),
			.E(gen[5746]),

			.SO(gen[5839]),
			.S(gen[5840]),
			.SE(gen[5841]),

			.SELF(gen[5745]),
			.cell_state(gen[5745])
		); 

/******************* CELL 5746 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5746 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5650]),
			.N(gen[5651]),
			.NE(gen[5652]),

			.O(gen[5745]),
			.E(gen[5747]),

			.SO(gen[5840]),
			.S(gen[5841]),
			.SE(gen[5842]),

			.SELF(gen[5746]),
			.cell_state(gen[5746])
		); 

/******************* CELL 5747 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5747 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5651]),
			.N(gen[5652]),
			.NE(gen[5653]),

			.O(gen[5746]),
			.E(gen[5748]),

			.SO(gen[5841]),
			.S(gen[5842]),
			.SE(gen[5843]),

			.SELF(gen[5747]),
			.cell_state(gen[5747])
		); 

/******************* CELL 5748 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5748 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5652]),
			.N(gen[5653]),
			.NE(gen[5654]),

			.O(gen[5747]),
			.E(gen[5749]),

			.SO(gen[5842]),
			.S(gen[5843]),
			.SE(gen[5844]),

			.SELF(gen[5748]),
			.cell_state(gen[5748])
		); 

/******************* CELL 5749 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5749 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5653]),
			.N(gen[5654]),
			.NE(gen[5655]),

			.O(gen[5748]),
			.E(gen[5750]),

			.SO(gen[5843]),
			.S(gen[5844]),
			.SE(gen[5845]),

			.SELF(gen[5749]),
			.cell_state(gen[5749])
		); 

/******************* CELL 5750 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5750 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5654]),
			.N(gen[5655]),
			.NE(gen[5656]),

			.O(gen[5749]),
			.E(gen[5751]),

			.SO(gen[5844]),
			.S(gen[5845]),
			.SE(gen[5846]),

			.SELF(gen[5750]),
			.cell_state(gen[5750])
		); 

/******************* CELL 5751 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5751 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5655]),
			.N(gen[5656]),
			.NE(gen[5657]),

			.O(gen[5750]),
			.E(gen[5752]),

			.SO(gen[5845]),
			.S(gen[5846]),
			.SE(gen[5847]),

			.SELF(gen[5751]),
			.cell_state(gen[5751])
		); 

/******************* CELL 5752 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5752 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5656]),
			.N(gen[5657]),
			.NE(gen[5658]),

			.O(gen[5751]),
			.E(gen[5753]),

			.SO(gen[5846]),
			.S(gen[5847]),
			.SE(gen[5848]),

			.SELF(gen[5752]),
			.cell_state(gen[5752])
		); 

/******************* CELL 5753 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5753 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5657]),
			.N(gen[5658]),
			.NE(gen[5659]),

			.O(gen[5752]),
			.E(gen[5754]),

			.SO(gen[5847]),
			.S(gen[5848]),
			.SE(gen[5849]),

			.SELF(gen[5753]),
			.cell_state(gen[5753])
		); 

/******************* CELL 5754 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5754 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5658]),
			.N(gen[5659]),
			.NE(gen[5660]),

			.O(gen[5753]),
			.E(gen[5755]),

			.SO(gen[5848]),
			.S(gen[5849]),
			.SE(gen[5850]),

			.SELF(gen[5754]),
			.cell_state(gen[5754])
		); 

/******************* CELL 5755 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5755 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5659]),
			.N(gen[5660]),
			.NE(gen[5661]),

			.O(gen[5754]),
			.E(gen[5756]),

			.SO(gen[5849]),
			.S(gen[5850]),
			.SE(gen[5851]),

			.SELF(gen[5755]),
			.cell_state(gen[5755])
		); 

/******************* CELL 5756 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5756 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5660]),
			.N(gen[5661]),
			.NE(gen[5662]),

			.O(gen[5755]),
			.E(gen[5757]),

			.SO(gen[5850]),
			.S(gen[5851]),
			.SE(gen[5852]),

			.SELF(gen[5756]),
			.cell_state(gen[5756])
		); 

/******************* CELL 5757 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5757 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5661]),
			.N(gen[5662]),
			.NE(gen[5663]),

			.O(gen[5756]),
			.E(gen[5758]),

			.SO(gen[5851]),
			.S(gen[5852]),
			.SE(gen[5853]),

			.SELF(gen[5757]),
			.cell_state(gen[5757])
		); 

/******************* CELL 5758 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5758 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5662]),
			.N(gen[5663]),
			.NE(gen[5664]),

			.O(gen[5757]),
			.E(gen[5759]),

			.SO(gen[5852]),
			.S(gen[5853]),
			.SE(gen[5854]),

			.SELF(gen[5758]),
			.cell_state(gen[5758])
		); 

/******************* CELL 5759 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5759 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5663]),
			.N(gen[5664]),
			.NE(gen[5665]),

			.O(gen[5758]),
			.E(gen[5760]),

			.SO(gen[5853]),
			.S(gen[5854]),
			.SE(gen[5855]),

			.SELF(gen[5759]),
			.cell_state(gen[5759])
		); 

/******************* CELL 5760 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5760 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5664]),
			.N(gen[5665]),
			.NE(gen[5666]),

			.O(gen[5759]),
			.E(gen[5761]),

			.SO(gen[5854]),
			.S(gen[5855]),
			.SE(gen[5856]),

			.SELF(gen[5760]),
			.cell_state(gen[5760])
		); 

/******************* CELL 5761 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5761 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5665]),
			.N(gen[5666]),
			.NE(gen[5667]),

			.O(gen[5760]),
			.E(gen[5762]),

			.SO(gen[5855]),
			.S(gen[5856]),
			.SE(gen[5857]),

			.SELF(gen[5761]),
			.cell_state(gen[5761])
		); 

/******************* CELL 5762 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5762 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5666]),
			.N(gen[5667]),
			.NE(gen[5668]),

			.O(gen[5761]),
			.E(gen[5763]),

			.SO(gen[5856]),
			.S(gen[5857]),
			.SE(gen[5858]),

			.SELF(gen[5762]),
			.cell_state(gen[5762])
		); 

/******************* CELL 5763 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5763 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5667]),
			.N(gen[5668]),
			.NE(gen[5669]),

			.O(gen[5762]),
			.E(gen[5764]),

			.SO(gen[5857]),
			.S(gen[5858]),
			.SE(gen[5859]),

			.SELF(gen[5763]),
			.cell_state(gen[5763])
		); 

/******************* CELL 5764 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5764 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5668]),
			.N(gen[5669]),
			.NE(gen[5670]),

			.O(gen[5763]),
			.E(gen[5765]),

			.SO(gen[5858]),
			.S(gen[5859]),
			.SE(gen[5860]),

			.SELF(gen[5764]),
			.cell_state(gen[5764])
		); 

/******************* CELL 5765 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5765 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5669]),
			.N(gen[5670]),
			.NE(gen[5671]),

			.O(gen[5764]),
			.E(gen[5766]),

			.SO(gen[5859]),
			.S(gen[5860]),
			.SE(gen[5861]),

			.SELF(gen[5765]),
			.cell_state(gen[5765])
		); 

/******************* CELL 5766 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5766 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5670]),
			.N(gen[5671]),
			.NE(gen[5672]),

			.O(gen[5765]),
			.E(gen[5767]),

			.SO(gen[5860]),
			.S(gen[5861]),
			.SE(gen[5862]),

			.SELF(gen[5766]),
			.cell_state(gen[5766])
		); 

/******************* CELL 5767 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5767 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5671]),
			.N(gen[5672]),
			.NE(gen[5673]),

			.O(gen[5766]),
			.E(gen[5768]),

			.SO(gen[5861]),
			.S(gen[5862]),
			.SE(gen[5863]),

			.SELF(gen[5767]),
			.cell_state(gen[5767])
		); 

/******************* CELL 5768 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5768 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5672]),
			.N(gen[5673]),
			.NE(gen[5674]),

			.O(gen[5767]),
			.E(gen[5769]),

			.SO(gen[5862]),
			.S(gen[5863]),
			.SE(gen[5864]),

			.SELF(gen[5768]),
			.cell_state(gen[5768])
		); 

/******************* CELL 5769 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5769 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5673]),
			.N(gen[5674]),
			.NE(gen[5675]),

			.O(gen[5768]),
			.E(gen[5770]),

			.SO(gen[5863]),
			.S(gen[5864]),
			.SE(gen[5865]),

			.SELF(gen[5769]),
			.cell_state(gen[5769])
		); 

/******************* CELL 5770 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5770 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5674]),
			.N(gen[5675]),
			.NE(gen[5676]),

			.O(gen[5769]),
			.E(gen[5771]),

			.SO(gen[5864]),
			.S(gen[5865]),
			.SE(gen[5866]),

			.SELF(gen[5770]),
			.cell_state(gen[5770])
		); 

/******************* CELL 5771 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5771 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5675]),
			.N(gen[5676]),
			.NE(gen[5677]),

			.O(gen[5770]),
			.E(gen[5772]),

			.SO(gen[5865]),
			.S(gen[5866]),
			.SE(gen[5867]),

			.SELF(gen[5771]),
			.cell_state(gen[5771])
		); 

/******************* CELL 5772 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5772 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5676]),
			.N(gen[5677]),
			.NE(gen[5678]),

			.O(gen[5771]),
			.E(gen[5773]),

			.SO(gen[5866]),
			.S(gen[5867]),
			.SE(gen[5868]),

			.SELF(gen[5772]),
			.cell_state(gen[5772])
		); 

/******************* CELL 5773 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5773 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5677]),
			.N(gen[5678]),
			.NE(gen[5679]),

			.O(gen[5772]),
			.E(gen[5774]),

			.SO(gen[5867]),
			.S(gen[5868]),
			.SE(gen[5869]),

			.SELF(gen[5773]),
			.cell_state(gen[5773])
		); 

/******************* CELL 5774 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5774 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5678]),
			.N(gen[5679]),
			.NE(gen[5680]),

			.O(gen[5773]),
			.E(gen[5775]),

			.SO(gen[5868]),
			.S(gen[5869]),
			.SE(gen[5870]),

			.SELF(gen[5774]),
			.cell_state(gen[5774])
		); 

/******************* CELL 5775 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5775 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5679]),
			.N(gen[5680]),
			.NE(gen[5681]),

			.O(gen[5774]),
			.E(gen[5776]),

			.SO(gen[5869]),
			.S(gen[5870]),
			.SE(gen[5871]),

			.SELF(gen[5775]),
			.cell_state(gen[5775])
		); 

/******************* CELL 5776 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5776 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5680]),
			.N(gen[5681]),
			.NE(gen[5682]),

			.O(gen[5775]),
			.E(gen[5777]),

			.SO(gen[5870]),
			.S(gen[5871]),
			.SE(gen[5872]),

			.SELF(gen[5776]),
			.cell_state(gen[5776])
		); 

/******************* CELL 5777 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5777 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5681]),
			.N(gen[5682]),
			.NE(gen[5683]),

			.O(gen[5776]),
			.E(gen[5778]),

			.SO(gen[5871]),
			.S(gen[5872]),
			.SE(gen[5873]),

			.SELF(gen[5777]),
			.cell_state(gen[5777])
		); 

/******************* CELL 5778 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5778 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5682]),
			.N(gen[5683]),
			.NE(gen[5684]),

			.O(gen[5777]),
			.E(gen[5779]),

			.SO(gen[5872]),
			.S(gen[5873]),
			.SE(gen[5874]),

			.SELF(gen[5778]),
			.cell_state(gen[5778])
		); 

/******************* CELL 5779 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5779 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5683]),
			.N(gen[5684]),
			.NE(gen[5685]),

			.O(gen[5778]),
			.E(gen[5780]),

			.SO(gen[5873]),
			.S(gen[5874]),
			.SE(gen[5875]),

			.SELF(gen[5779]),
			.cell_state(gen[5779])
		); 

/******************* CELL 5780 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5780 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5684]),
			.N(gen[5685]),
			.NE(gen[5686]),

			.O(gen[5779]),
			.E(gen[5781]),

			.SO(gen[5874]),
			.S(gen[5875]),
			.SE(gen[5876]),

			.SELF(gen[5780]),
			.cell_state(gen[5780])
		); 

/******************* CELL 5781 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5781 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5685]),
			.N(gen[5686]),
			.NE(gen[5687]),

			.O(gen[5780]),
			.E(gen[5782]),

			.SO(gen[5875]),
			.S(gen[5876]),
			.SE(gen[5877]),

			.SELF(gen[5781]),
			.cell_state(gen[5781])
		); 

/******************* CELL 5782 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5782 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5686]),
			.N(gen[5687]),
			.NE(gen[5688]),

			.O(gen[5781]),
			.E(gen[5783]),

			.SO(gen[5876]),
			.S(gen[5877]),
			.SE(gen[5878]),

			.SELF(gen[5782]),
			.cell_state(gen[5782])
		); 

/******************* CELL 5783 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5783 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5687]),
			.N(gen[5688]),
			.NE(gen[5689]),

			.O(gen[5782]),
			.E(gen[5784]),

			.SO(gen[5877]),
			.S(gen[5878]),
			.SE(gen[5879]),

			.SELF(gen[5783]),
			.cell_state(gen[5783])
		); 

/******************* CELL 5784 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5784 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5688]),
			.N(gen[5689]),
			.NE(gen[5690]),

			.O(gen[5783]),
			.E(gen[5785]),

			.SO(gen[5878]),
			.S(gen[5879]),
			.SE(gen[5880]),

			.SELF(gen[5784]),
			.cell_state(gen[5784])
		); 

/******************* CELL 5785 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5785 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5689]),
			.N(gen[5690]),
			.NE(gen[5691]),

			.O(gen[5784]),
			.E(gen[5786]),

			.SO(gen[5879]),
			.S(gen[5880]),
			.SE(gen[5881]),

			.SELF(gen[5785]),
			.cell_state(gen[5785])
		); 

/******************* CELL 5786 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5786 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5690]),
			.N(gen[5691]),
			.NE(gen[5692]),

			.O(gen[5785]),
			.E(gen[5787]),

			.SO(gen[5880]),
			.S(gen[5881]),
			.SE(gen[5882]),

			.SELF(gen[5786]),
			.cell_state(gen[5786])
		); 

/******************* CELL 5787 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5787 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5691]),
			.N(gen[5692]),
			.NE(gen[5693]),

			.O(gen[5786]),
			.E(gen[5788]),

			.SO(gen[5881]),
			.S(gen[5882]),
			.SE(gen[5883]),

			.SELF(gen[5787]),
			.cell_state(gen[5787])
		); 

/******************* CELL 5788 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5788 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5692]),
			.N(gen[5693]),
			.NE(gen[5694]),

			.O(gen[5787]),
			.E(gen[5789]),

			.SO(gen[5882]),
			.S(gen[5883]),
			.SE(gen[5884]),

			.SELF(gen[5788]),
			.cell_state(gen[5788])
		); 

/******************* CELL 5789 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5789 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5693]),
			.N(gen[5694]),
			.NE(gen[5695]),

			.O(gen[5788]),
			.E(gen[5790]),

			.SO(gen[5883]),
			.S(gen[5884]),
			.SE(gen[5885]),

			.SELF(gen[5789]),
			.cell_state(gen[5789])
		); 

/******************* CELL 5790 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5790 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5694]),
			.N(gen[5695]),
			.NE(gen[5696]),

			.O(gen[5789]),
			.E(gen[5791]),

			.SO(gen[5884]),
			.S(gen[5885]),
			.SE(gen[5886]),

			.SELF(gen[5790]),
			.cell_state(gen[5790])
		); 

/******************* CELL 5791 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5791 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5695]),
			.N(gen[5696]),
			.NE(gen[5697]),

			.O(gen[5790]),
			.E(gen[5792]),

			.SO(gen[5885]),
			.S(gen[5886]),
			.SE(gen[5887]),

			.SELF(gen[5791]),
			.cell_state(gen[5791])
		); 

/******************* CELL 5792 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5792 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5696]),
			.N(gen[5697]),
			.NE(gen[5698]),

			.O(gen[5791]),
			.E(gen[5793]),

			.SO(gen[5886]),
			.S(gen[5887]),
			.SE(gen[5888]),

			.SELF(gen[5792]),
			.cell_state(gen[5792])
		); 

/******************* CELL 5793 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5793 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5697]),
			.N(gen[5698]),
			.NE(gen[5699]),

			.O(gen[5792]),
			.E(gen[5794]),

			.SO(gen[5887]),
			.S(gen[5888]),
			.SE(gen[5889]),

			.SELF(gen[5793]),
			.cell_state(gen[5793])
		); 

/******************* CELL 5794 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5794 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5698]),
			.N(gen[5699]),
			.NE(gen[5698]),

			.O(gen[5793]),
			.E(gen[5793]),

			.SO(gen[5888]),
			.S(gen[5889]),
			.SE(gen[5888]),

			.SELF(gen[5794]),
			.cell_state(gen[5794])
		); 

/******************* CELL 5795 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5795 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5701]),
			.N(gen[5700]),
			.NE(gen[5701]),

			.O(gen[5796]),
			.E(gen[5796]),

			.SO(gen[5891]),
			.S(gen[5890]),
			.SE(gen[5891]),

			.SELF(gen[5795]),
			.cell_state(gen[5795])
		); 

/******************* CELL 5796 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5796 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5700]),
			.N(gen[5701]),
			.NE(gen[5702]),

			.O(gen[5795]),
			.E(gen[5797]),

			.SO(gen[5890]),
			.S(gen[5891]),
			.SE(gen[5892]),

			.SELF(gen[5796]),
			.cell_state(gen[5796])
		); 

/******************* CELL 5797 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5797 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5701]),
			.N(gen[5702]),
			.NE(gen[5703]),

			.O(gen[5796]),
			.E(gen[5798]),

			.SO(gen[5891]),
			.S(gen[5892]),
			.SE(gen[5893]),

			.SELF(gen[5797]),
			.cell_state(gen[5797])
		); 

/******************* CELL 5798 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5798 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5702]),
			.N(gen[5703]),
			.NE(gen[5704]),

			.O(gen[5797]),
			.E(gen[5799]),

			.SO(gen[5892]),
			.S(gen[5893]),
			.SE(gen[5894]),

			.SELF(gen[5798]),
			.cell_state(gen[5798])
		); 

/******************* CELL 5799 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5799 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5703]),
			.N(gen[5704]),
			.NE(gen[5705]),

			.O(gen[5798]),
			.E(gen[5800]),

			.SO(gen[5893]),
			.S(gen[5894]),
			.SE(gen[5895]),

			.SELF(gen[5799]),
			.cell_state(gen[5799])
		); 

/******************* CELL 5800 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5800 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5704]),
			.N(gen[5705]),
			.NE(gen[5706]),

			.O(gen[5799]),
			.E(gen[5801]),

			.SO(gen[5894]),
			.S(gen[5895]),
			.SE(gen[5896]),

			.SELF(gen[5800]),
			.cell_state(gen[5800])
		); 

/******************* CELL 5801 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5801 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5705]),
			.N(gen[5706]),
			.NE(gen[5707]),

			.O(gen[5800]),
			.E(gen[5802]),

			.SO(gen[5895]),
			.S(gen[5896]),
			.SE(gen[5897]),

			.SELF(gen[5801]),
			.cell_state(gen[5801])
		); 

/******************* CELL 5802 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5802 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5706]),
			.N(gen[5707]),
			.NE(gen[5708]),

			.O(gen[5801]),
			.E(gen[5803]),

			.SO(gen[5896]),
			.S(gen[5897]),
			.SE(gen[5898]),

			.SELF(gen[5802]),
			.cell_state(gen[5802])
		); 

/******************* CELL 5803 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5803 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5707]),
			.N(gen[5708]),
			.NE(gen[5709]),

			.O(gen[5802]),
			.E(gen[5804]),

			.SO(gen[5897]),
			.S(gen[5898]),
			.SE(gen[5899]),

			.SELF(gen[5803]),
			.cell_state(gen[5803])
		); 

/******************* CELL 5804 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5804 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5708]),
			.N(gen[5709]),
			.NE(gen[5710]),

			.O(gen[5803]),
			.E(gen[5805]),

			.SO(gen[5898]),
			.S(gen[5899]),
			.SE(gen[5900]),

			.SELF(gen[5804]),
			.cell_state(gen[5804])
		); 

/******************* CELL 5805 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5805 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5709]),
			.N(gen[5710]),
			.NE(gen[5711]),

			.O(gen[5804]),
			.E(gen[5806]),

			.SO(gen[5899]),
			.S(gen[5900]),
			.SE(gen[5901]),

			.SELF(gen[5805]),
			.cell_state(gen[5805])
		); 

/******************* CELL 5806 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5806 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5710]),
			.N(gen[5711]),
			.NE(gen[5712]),

			.O(gen[5805]),
			.E(gen[5807]),

			.SO(gen[5900]),
			.S(gen[5901]),
			.SE(gen[5902]),

			.SELF(gen[5806]),
			.cell_state(gen[5806])
		); 

/******************* CELL 5807 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5807 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5711]),
			.N(gen[5712]),
			.NE(gen[5713]),

			.O(gen[5806]),
			.E(gen[5808]),

			.SO(gen[5901]),
			.S(gen[5902]),
			.SE(gen[5903]),

			.SELF(gen[5807]),
			.cell_state(gen[5807])
		); 

/******************* CELL 5808 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5808 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5712]),
			.N(gen[5713]),
			.NE(gen[5714]),

			.O(gen[5807]),
			.E(gen[5809]),

			.SO(gen[5902]),
			.S(gen[5903]),
			.SE(gen[5904]),

			.SELF(gen[5808]),
			.cell_state(gen[5808])
		); 

/******************* CELL 5809 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5809 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5713]),
			.N(gen[5714]),
			.NE(gen[5715]),

			.O(gen[5808]),
			.E(gen[5810]),

			.SO(gen[5903]),
			.S(gen[5904]),
			.SE(gen[5905]),

			.SELF(gen[5809]),
			.cell_state(gen[5809])
		); 

/******************* CELL 5810 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5810 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5714]),
			.N(gen[5715]),
			.NE(gen[5716]),

			.O(gen[5809]),
			.E(gen[5811]),

			.SO(gen[5904]),
			.S(gen[5905]),
			.SE(gen[5906]),

			.SELF(gen[5810]),
			.cell_state(gen[5810])
		); 

/******************* CELL 5811 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5811 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5715]),
			.N(gen[5716]),
			.NE(gen[5717]),

			.O(gen[5810]),
			.E(gen[5812]),

			.SO(gen[5905]),
			.S(gen[5906]),
			.SE(gen[5907]),

			.SELF(gen[5811]),
			.cell_state(gen[5811])
		); 

/******************* CELL 5812 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5812 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5716]),
			.N(gen[5717]),
			.NE(gen[5718]),

			.O(gen[5811]),
			.E(gen[5813]),

			.SO(gen[5906]),
			.S(gen[5907]),
			.SE(gen[5908]),

			.SELF(gen[5812]),
			.cell_state(gen[5812])
		); 

/******************* CELL 5813 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5813 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5717]),
			.N(gen[5718]),
			.NE(gen[5719]),

			.O(gen[5812]),
			.E(gen[5814]),

			.SO(gen[5907]),
			.S(gen[5908]),
			.SE(gen[5909]),

			.SELF(gen[5813]),
			.cell_state(gen[5813])
		); 

/******************* CELL 5814 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5814 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5718]),
			.N(gen[5719]),
			.NE(gen[5720]),

			.O(gen[5813]),
			.E(gen[5815]),

			.SO(gen[5908]),
			.S(gen[5909]),
			.SE(gen[5910]),

			.SELF(gen[5814]),
			.cell_state(gen[5814])
		); 

/******************* CELL 5815 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5815 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5719]),
			.N(gen[5720]),
			.NE(gen[5721]),

			.O(gen[5814]),
			.E(gen[5816]),

			.SO(gen[5909]),
			.S(gen[5910]),
			.SE(gen[5911]),

			.SELF(gen[5815]),
			.cell_state(gen[5815])
		); 

/******************* CELL 5816 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5816 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5720]),
			.N(gen[5721]),
			.NE(gen[5722]),

			.O(gen[5815]),
			.E(gen[5817]),

			.SO(gen[5910]),
			.S(gen[5911]),
			.SE(gen[5912]),

			.SELF(gen[5816]),
			.cell_state(gen[5816])
		); 

/******************* CELL 5817 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5817 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5721]),
			.N(gen[5722]),
			.NE(gen[5723]),

			.O(gen[5816]),
			.E(gen[5818]),

			.SO(gen[5911]),
			.S(gen[5912]),
			.SE(gen[5913]),

			.SELF(gen[5817]),
			.cell_state(gen[5817])
		); 

/******************* CELL 5818 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5818 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5722]),
			.N(gen[5723]),
			.NE(gen[5724]),

			.O(gen[5817]),
			.E(gen[5819]),

			.SO(gen[5912]),
			.S(gen[5913]),
			.SE(gen[5914]),

			.SELF(gen[5818]),
			.cell_state(gen[5818])
		); 

/******************* CELL 5819 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5819 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5723]),
			.N(gen[5724]),
			.NE(gen[5725]),

			.O(gen[5818]),
			.E(gen[5820]),

			.SO(gen[5913]),
			.S(gen[5914]),
			.SE(gen[5915]),

			.SELF(gen[5819]),
			.cell_state(gen[5819])
		); 

/******************* CELL 5820 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5820 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5724]),
			.N(gen[5725]),
			.NE(gen[5726]),

			.O(gen[5819]),
			.E(gen[5821]),

			.SO(gen[5914]),
			.S(gen[5915]),
			.SE(gen[5916]),

			.SELF(gen[5820]),
			.cell_state(gen[5820])
		); 

/******************* CELL 5821 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5821 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5725]),
			.N(gen[5726]),
			.NE(gen[5727]),

			.O(gen[5820]),
			.E(gen[5822]),

			.SO(gen[5915]),
			.S(gen[5916]),
			.SE(gen[5917]),

			.SELF(gen[5821]),
			.cell_state(gen[5821])
		); 

/******************* CELL 5822 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5822 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5726]),
			.N(gen[5727]),
			.NE(gen[5728]),

			.O(gen[5821]),
			.E(gen[5823]),

			.SO(gen[5916]),
			.S(gen[5917]),
			.SE(gen[5918]),

			.SELF(gen[5822]),
			.cell_state(gen[5822])
		); 

/******************* CELL 5823 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5823 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5727]),
			.N(gen[5728]),
			.NE(gen[5729]),

			.O(gen[5822]),
			.E(gen[5824]),

			.SO(gen[5917]),
			.S(gen[5918]),
			.SE(gen[5919]),

			.SELF(gen[5823]),
			.cell_state(gen[5823])
		); 

/******************* CELL 5824 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5824 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5728]),
			.N(gen[5729]),
			.NE(gen[5730]),

			.O(gen[5823]),
			.E(gen[5825]),

			.SO(gen[5918]),
			.S(gen[5919]),
			.SE(gen[5920]),

			.SELF(gen[5824]),
			.cell_state(gen[5824])
		); 

/******************* CELL 5825 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5825 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5729]),
			.N(gen[5730]),
			.NE(gen[5731]),

			.O(gen[5824]),
			.E(gen[5826]),

			.SO(gen[5919]),
			.S(gen[5920]),
			.SE(gen[5921]),

			.SELF(gen[5825]),
			.cell_state(gen[5825])
		); 

/******************* CELL 5826 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5826 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5730]),
			.N(gen[5731]),
			.NE(gen[5732]),

			.O(gen[5825]),
			.E(gen[5827]),

			.SO(gen[5920]),
			.S(gen[5921]),
			.SE(gen[5922]),

			.SELF(gen[5826]),
			.cell_state(gen[5826])
		); 

/******************* CELL 5827 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5827 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5731]),
			.N(gen[5732]),
			.NE(gen[5733]),

			.O(gen[5826]),
			.E(gen[5828]),

			.SO(gen[5921]),
			.S(gen[5922]),
			.SE(gen[5923]),

			.SELF(gen[5827]),
			.cell_state(gen[5827])
		); 

/******************* CELL 5828 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5828 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5732]),
			.N(gen[5733]),
			.NE(gen[5734]),

			.O(gen[5827]),
			.E(gen[5829]),

			.SO(gen[5922]),
			.S(gen[5923]),
			.SE(gen[5924]),

			.SELF(gen[5828]),
			.cell_state(gen[5828])
		); 

/******************* CELL 5829 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5829 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5733]),
			.N(gen[5734]),
			.NE(gen[5735]),

			.O(gen[5828]),
			.E(gen[5830]),

			.SO(gen[5923]),
			.S(gen[5924]),
			.SE(gen[5925]),

			.SELF(gen[5829]),
			.cell_state(gen[5829])
		); 

/******************* CELL 5830 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5830 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5734]),
			.N(gen[5735]),
			.NE(gen[5736]),

			.O(gen[5829]),
			.E(gen[5831]),

			.SO(gen[5924]),
			.S(gen[5925]),
			.SE(gen[5926]),

			.SELF(gen[5830]),
			.cell_state(gen[5830])
		); 

/******************* CELL 5831 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5831 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5735]),
			.N(gen[5736]),
			.NE(gen[5737]),

			.O(gen[5830]),
			.E(gen[5832]),

			.SO(gen[5925]),
			.S(gen[5926]),
			.SE(gen[5927]),

			.SELF(gen[5831]),
			.cell_state(gen[5831])
		); 

/******************* CELL 5832 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5832 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5736]),
			.N(gen[5737]),
			.NE(gen[5738]),

			.O(gen[5831]),
			.E(gen[5833]),

			.SO(gen[5926]),
			.S(gen[5927]),
			.SE(gen[5928]),

			.SELF(gen[5832]),
			.cell_state(gen[5832])
		); 

/******************* CELL 5833 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5833 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5737]),
			.N(gen[5738]),
			.NE(gen[5739]),

			.O(gen[5832]),
			.E(gen[5834]),

			.SO(gen[5927]),
			.S(gen[5928]),
			.SE(gen[5929]),

			.SELF(gen[5833]),
			.cell_state(gen[5833])
		); 

/******************* CELL 5834 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5834 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5738]),
			.N(gen[5739]),
			.NE(gen[5740]),

			.O(gen[5833]),
			.E(gen[5835]),

			.SO(gen[5928]),
			.S(gen[5929]),
			.SE(gen[5930]),

			.SELF(gen[5834]),
			.cell_state(gen[5834])
		); 

/******************* CELL 5835 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5835 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5739]),
			.N(gen[5740]),
			.NE(gen[5741]),

			.O(gen[5834]),
			.E(gen[5836]),

			.SO(gen[5929]),
			.S(gen[5930]),
			.SE(gen[5931]),

			.SELF(gen[5835]),
			.cell_state(gen[5835])
		); 

/******************* CELL 5836 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5836 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5740]),
			.N(gen[5741]),
			.NE(gen[5742]),

			.O(gen[5835]),
			.E(gen[5837]),

			.SO(gen[5930]),
			.S(gen[5931]),
			.SE(gen[5932]),

			.SELF(gen[5836]),
			.cell_state(gen[5836])
		); 

/******************* CELL 5837 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5837 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5741]),
			.N(gen[5742]),
			.NE(gen[5743]),

			.O(gen[5836]),
			.E(gen[5838]),

			.SO(gen[5931]),
			.S(gen[5932]),
			.SE(gen[5933]),

			.SELF(gen[5837]),
			.cell_state(gen[5837])
		); 

/******************* CELL 5838 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5838 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5742]),
			.N(gen[5743]),
			.NE(gen[5744]),

			.O(gen[5837]),
			.E(gen[5839]),

			.SO(gen[5932]),
			.S(gen[5933]),
			.SE(gen[5934]),

			.SELF(gen[5838]),
			.cell_state(gen[5838])
		); 

/******************* CELL 5839 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5839 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5743]),
			.N(gen[5744]),
			.NE(gen[5745]),

			.O(gen[5838]),
			.E(gen[5840]),

			.SO(gen[5933]),
			.S(gen[5934]),
			.SE(gen[5935]),

			.SELF(gen[5839]),
			.cell_state(gen[5839])
		); 

/******************* CELL 5840 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5840 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5744]),
			.N(gen[5745]),
			.NE(gen[5746]),

			.O(gen[5839]),
			.E(gen[5841]),

			.SO(gen[5934]),
			.S(gen[5935]),
			.SE(gen[5936]),

			.SELF(gen[5840]),
			.cell_state(gen[5840])
		); 

/******************* CELL 5841 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5841 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5745]),
			.N(gen[5746]),
			.NE(gen[5747]),

			.O(gen[5840]),
			.E(gen[5842]),

			.SO(gen[5935]),
			.S(gen[5936]),
			.SE(gen[5937]),

			.SELF(gen[5841]),
			.cell_state(gen[5841])
		); 

/******************* CELL 5842 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5842 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5746]),
			.N(gen[5747]),
			.NE(gen[5748]),

			.O(gen[5841]),
			.E(gen[5843]),

			.SO(gen[5936]),
			.S(gen[5937]),
			.SE(gen[5938]),

			.SELF(gen[5842]),
			.cell_state(gen[5842])
		); 

/******************* CELL 5843 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5843 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5747]),
			.N(gen[5748]),
			.NE(gen[5749]),

			.O(gen[5842]),
			.E(gen[5844]),

			.SO(gen[5937]),
			.S(gen[5938]),
			.SE(gen[5939]),

			.SELF(gen[5843]),
			.cell_state(gen[5843])
		); 

/******************* CELL 5844 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5844 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5748]),
			.N(gen[5749]),
			.NE(gen[5750]),

			.O(gen[5843]),
			.E(gen[5845]),

			.SO(gen[5938]),
			.S(gen[5939]),
			.SE(gen[5940]),

			.SELF(gen[5844]),
			.cell_state(gen[5844])
		); 

/******************* CELL 5845 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5845 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5749]),
			.N(gen[5750]),
			.NE(gen[5751]),

			.O(gen[5844]),
			.E(gen[5846]),

			.SO(gen[5939]),
			.S(gen[5940]),
			.SE(gen[5941]),

			.SELF(gen[5845]),
			.cell_state(gen[5845])
		); 

/******************* CELL 5846 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5846 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5750]),
			.N(gen[5751]),
			.NE(gen[5752]),

			.O(gen[5845]),
			.E(gen[5847]),

			.SO(gen[5940]),
			.S(gen[5941]),
			.SE(gen[5942]),

			.SELF(gen[5846]),
			.cell_state(gen[5846])
		); 

/******************* CELL 5847 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5847 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5751]),
			.N(gen[5752]),
			.NE(gen[5753]),

			.O(gen[5846]),
			.E(gen[5848]),

			.SO(gen[5941]),
			.S(gen[5942]),
			.SE(gen[5943]),

			.SELF(gen[5847]),
			.cell_state(gen[5847])
		); 

/******************* CELL 5848 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5848 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5752]),
			.N(gen[5753]),
			.NE(gen[5754]),

			.O(gen[5847]),
			.E(gen[5849]),

			.SO(gen[5942]),
			.S(gen[5943]),
			.SE(gen[5944]),

			.SELF(gen[5848]),
			.cell_state(gen[5848])
		); 

/******************* CELL 5849 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5849 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5753]),
			.N(gen[5754]),
			.NE(gen[5755]),

			.O(gen[5848]),
			.E(gen[5850]),

			.SO(gen[5943]),
			.S(gen[5944]),
			.SE(gen[5945]),

			.SELF(gen[5849]),
			.cell_state(gen[5849])
		); 

/******************* CELL 5850 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5850 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5754]),
			.N(gen[5755]),
			.NE(gen[5756]),

			.O(gen[5849]),
			.E(gen[5851]),

			.SO(gen[5944]),
			.S(gen[5945]),
			.SE(gen[5946]),

			.SELF(gen[5850]),
			.cell_state(gen[5850])
		); 

/******************* CELL 5851 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5851 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5755]),
			.N(gen[5756]),
			.NE(gen[5757]),

			.O(gen[5850]),
			.E(gen[5852]),

			.SO(gen[5945]),
			.S(gen[5946]),
			.SE(gen[5947]),

			.SELF(gen[5851]),
			.cell_state(gen[5851])
		); 

/******************* CELL 5852 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5852 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5756]),
			.N(gen[5757]),
			.NE(gen[5758]),

			.O(gen[5851]),
			.E(gen[5853]),

			.SO(gen[5946]),
			.S(gen[5947]),
			.SE(gen[5948]),

			.SELF(gen[5852]),
			.cell_state(gen[5852])
		); 

/******************* CELL 5853 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5853 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5757]),
			.N(gen[5758]),
			.NE(gen[5759]),

			.O(gen[5852]),
			.E(gen[5854]),

			.SO(gen[5947]),
			.S(gen[5948]),
			.SE(gen[5949]),

			.SELF(gen[5853]),
			.cell_state(gen[5853])
		); 

/******************* CELL 5854 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5854 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5758]),
			.N(gen[5759]),
			.NE(gen[5760]),

			.O(gen[5853]),
			.E(gen[5855]),

			.SO(gen[5948]),
			.S(gen[5949]),
			.SE(gen[5950]),

			.SELF(gen[5854]),
			.cell_state(gen[5854])
		); 

/******************* CELL 5855 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5855 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5759]),
			.N(gen[5760]),
			.NE(gen[5761]),

			.O(gen[5854]),
			.E(gen[5856]),

			.SO(gen[5949]),
			.S(gen[5950]),
			.SE(gen[5951]),

			.SELF(gen[5855]),
			.cell_state(gen[5855])
		); 

/******************* CELL 5856 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5856 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5760]),
			.N(gen[5761]),
			.NE(gen[5762]),

			.O(gen[5855]),
			.E(gen[5857]),

			.SO(gen[5950]),
			.S(gen[5951]),
			.SE(gen[5952]),

			.SELF(gen[5856]),
			.cell_state(gen[5856])
		); 

/******************* CELL 5857 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5857 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5761]),
			.N(gen[5762]),
			.NE(gen[5763]),

			.O(gen[5856]),
			.E(gen[5858]),

			.SO(gen[5951]),
			.S(gen[5952]),
			.SE(gen[5953]),

			.SELF(gen[5857]),
			.cell_state(gen[5857])
		); 

/******************* CELL 5858 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5858 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5762]),
			.N(gen[5763]),
			.NE(gen[5764]),

			.O(gen[5857]),
			.E(gen[5859]),

			.SO(gen[5952]),
			.S(gen[5953]),
			.SE(gen[5954]),

			.SELF(gen[5858]),
			.cell_state(gen[5858])
		); 

/******************* CELL 5859 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5859 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5763]),
			.N(gen[5764]),
			.NE(gen[5765]),

			.O(gen[5858]),
			.E(gen[5860]),

			.SO(gen[5953]),
			.S(gen[5954]),
			.SE(gen[5955]),

			.SELF(gen[5859]),
			.cell_state(gen[5859])
		); 

/******************* CELL 5860 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5860 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5764]),
			.N(gen[5765]),
			.NE(gen[5766]),

			.O(gen[5859]),
			.E(gen[5861]),

			.SO(gen[5954]),
			.S(gen[5955]),
			.SE(gen[5956]),

			.SELF(gen[5860]),
			.cell_state(gen[5860])
		); 

/******************* CELL 5861 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5861 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5765]),
			.N(gen[5766]),
			.NE(gen[5767]),

			.O(gen[5860]),
			.E(gen[5862]),

			.SO(gen[5955]),
			.S(gen[5956]),
			.SE(gen[5957]),

			.SELF(gen[5861]),
			.cell_state(gen[5861])
		); 

/******************* CELL 5862 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5862 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5766]),
			.N(gen[5767]),
			.NE(gen[5768]),

			.O(gen[5861]),
			.E(gen[5863]),

			.SO(gen[5956]),
			.S(gen[5957]),
			.SE(gen[5958]),

			.SELF(gen[5862]),
			.cell_state(gen[5862])
		); 

/******************* CELL 5863 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5863 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5767]),
			.N(gen[5768]),
			.NE(gen[5769]),

			.O(gen[5862]),
			.E(gen[5864]),

			.SO(gen[5957]),
			.S(gen[5958]),
			.SE(gen[5959]),

			.SELF(gen[5863]),
			.cell_state(gen[5863])
		); 

/******************* CELL 5864 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5864 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5768]),
			.N(gen[5769]),
			.NE(gen[5770]),

			.O(gen[5863]),
			.E(gen[5865]),

			.SO(gen[5958]),
			.S(gen[5959]),
			.SE(gen[5960]),

			.SELF(gen[5864]),
			.cell_state(gen[5864])
		); 

/******************* CELL 5865 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5865 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5769]),
			.N(gen[5770]),
			.NE(gen[5771]),

			.O(gen[5864]),
			.E(gen[5866]),

			.SO(gen[5959]),
			.S(gen[5960]),
			.SE(gen[5961]),

			.SELF(gen[5865]),
			.cell_state(gen[5865])
		); 

/******************* CELL 5866 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5866 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5770]),
			.N(gen[5771]),
			.NE(gen[5772]),

			.O(gen[5865]),
			.E(gen[5867]),

			.SO(gen[5960]),
			.S(gen[5961]),
			.SE(gen[5962]),

			.SELF(gen[5866]),
			.cell_state(gen[5866])
		); 

/******************* CELL 5867 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5867 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5771]),
			.N(gen[5772]),
			.NE(gen[5773]),

			.O(gen[5866]),
			.E(gen[5868]),

			.SO(gen[5961]),
			.S(gen[5962]),
			.SE(gen[5963]),

			.SELF(gen[5867]),
			.cell_state(gen[5867])
		); 

/******************* CELL 5868 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5868 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5772]),
			.N(gen[5773]),
			.NE(gen[5774]),

			.O(gen[5867]),
			.E(gen[5869]),

			.SO(gen[5962]),
			.S(gen[5963]),
			.SE(gen[5964]),

			.SELF(gen[5868]),
			.cell_state(gen[5868])
		); 

/******************* CELL 5869 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5869 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5773]),
			.N(gen[5774]),
			.NE(gen[5775]),

			.O(gen[5868]),
			.E(gen[5870]),

			.SO(gen[5963]),
			.S(gen[5964]),
			.SE(gen[5965]),

			.SELF(gen[5869]),
			.cell_state(gen[5869])
		); 

/******************* CELL 5870 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5870 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5774]),
			.N(gen[5775]),
			.NE(gen[5776]),

			.O(gen[5869]),
			.E(gen[5871]),

			.SO(gen[5964]),
			.S(gen[5965]),
			.SE(gen[5966]),

			.SELF(gen[5870]),
			.cell_state(gen[5870])
		); 

/******************* CELL 5871 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5871 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5775]),
			.N(gen[5776]),
			.NE(gen[5777]),

			.O(gen[5870]),
			.E(gen[5872]),

			.SO(gen[5965]),
			.S(gen[5966]),
			.SE(gen[5967]),

			.SELF(gen[5871]),
			.cell_state(gen[5871])
		); 

/******************* CELL 5872 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5872 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5776]),
			.N(gen[5777]),
			.NE(gen[5778]),

			.O(gen[5871]),
			.E(gen[5873]),

			.SO(gen[5966]),
			.S(gen[5967]),
			.SE(gen[5968]),

			.SELF(gen[5872]),
			.cell_state(gen[5872])
		); 

/******************* CELL 5873 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5873 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5777]),
			.N(gen[5778]),
			.NE(gen[5779]),

			.O(gen[5872]),
			.E(gen[5874]),

			.SO(gen[5967]),
			.S(gen[5968]),
			.SE(gen[5969]),

			.SELF(gen[5873]),
			.cell_state(gen[5873])
		); 

/******************* CELL 5874 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5874 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5778]),
			.N(gen[5779]),
			.NE(gen[5780]),

			.O(gen[5873]),
			.E(gen[5875]),

			.SO(gen[5968]),
			.S(gen[5969]),
			.SE(gen[5970]),

			.SELF(gen[5874]),
			.cell_state(gen[5874])
		); 

/******************* CELL 5875 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5875 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5779]),
			.N(gen[5780]),
			.NE(gen[5781]),

			.O(gen[5874]),
			.E(gen[5876]),

			.SO(gen[5969]),
			.S(gen[5970]),
			.SE(gen[5971]),

			.SELF(gen[5875]),
			.cell_state(gen[5875])
		); 

/******************* CELL 5876 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5876 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5780]),
			.N(gen[5781]),
			.NE(gen[5782]),

			.O(gen[5875]),
			.E(gen[5877]),

			.SO(gen[5970]),
			.S(gen[5971]),
			.SE(gen[5972]),

			.SELF(gen[5876]),
			.cell_state(gen[5876])
		); 

/******************* CELL 5877 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5877 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5781]),
			.N(gen[5782]),
			.NE(gen[5783]),

			.O(gen[5876]),
			.E(gen[5878]),

			.SO(gen[5971]),
			.S(gen[5972]),
			.SE(gen[5973]),

			.SELF(gen[5877]),
			.cell_state(gen[5877])
		); 

/******************* CELL 5878 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5878 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5782]),
			.N(gen[5783]),
			.NE(gen[5784]),

			.O(gen[5877]),
			.E(gen[5879]),

			.SO(gen[5972]),
			.S(gen[5973]),
			.SE(gen[5974]),

			.SELF(gen[5878]),
			.cell_state(gen[5878])
		); 

/******************* CELL 5879 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5879 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5783]),
			.N(gen[5784]),
			.NE(gen[5785]),

			.O(gen[5878]),
			.E(gen[5880]),

			.SO(gen[5973]),
			.S(gen[5974]),
			.SE(gen[5975]),

			.SELF(gen[5879]),
			.cell_state(gen[5879])
		); 

/******************* CELL 5880 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5880 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5784]),
			.N(gen[5785]),
			.NE(gen[5786]),

			.O(gen[5879]),
			.E(gen[5881]),

			.SO(gen[5974]),
			.S(gen[5975]),
			.SE(gen[5976]),

			.SELF(gen[5880]),
			.cell_state(gen[5880])
		); 

/******************* CELL 5881 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5881 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5785]),
			.N(gen[5786]),
			.NE(gen[5787]),

			.O(gen[5880]),
			.E(gen[5882]),

			.SO(gen[5975]),
			.S(gen[5976]),
			.SE(gen[5977]),

			.SELF(gen[5881]),
			.cell_state(gen[5881])
		); 

/******************* CELL 5882 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5882 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5786]),
			.N(gen[5787]),
			.NE(gen[5788]),

			.O(gen[5881]),
			.E(gen[5883]),

			.SO(gen[5976]),
			.S(gen[5977]),
			.SE(gen[5978]),

			.SELF(gen[5882]),
			.cell_state(gen[5882])
		); 

/******************* CELL 5883 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5883 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5787]),
			.N(gen[5788]),
			.NE(gen[5789]),

			.O(gen[5882]),
			.E(gen[5884]),

			.SO(gen[5977]),
			.S(gen[5978]),
			.SE(gen[5979]),

			.SELF(gen[5883]),
			.cell_state(gen[5883])
		); 

/******************* CELL 5884 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5884 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5788]),
			.N(gen[5789]),
			.NE(gen[5790]),

			.O(gen[5883]),
			.E(gen[5885]),

			.SO(gen[5978]),
			.S(gen[5979]),
			.SE(gen[5980]),

			.SELF(gen[5884]),
			.cell_state(gen[5884])
		); 

/******************* CELL 5885 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5885 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5789]),
			.N(gen[5790]),
			.NE(gen[5791]),

			.O(gen[5884]),
			.E(gen[5886]),

			.SO(gen[5979]),
			.S(gen[5980]),
			.SE(gen[5981]),

			.SELF(gen[5885]),
			.cell_state(gen[5885])
		); 

/******************* CELL 5886 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5886 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5790]),
			.N(gen[5791]),
			.NE(gen[5792]),

			.O(gen[5885]),
			.E(gen[5887]),

			.SO(gen[5980]),
			.S(gen[5981]),
			.SE(gen[5982]),

			.SELF(gen[5886]),
			.cell_state(gen[5886])
		); 

/******************* CELL 5887 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5887 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5791]),
			.N(gen[5792]),
			.NE(gen[5793]),

			.O(gen[5886]),
			.E(gen[5888]),

			.SO(gen[5981]),
			.S(gen[5982]),
			.SE(gen[5983]),

			.SELF(gen[5887]),
			.cell_state(gen[5887])
		); 

/******************* CELL 5888 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5888 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5792]),
			.N(gen[5793]),
			.NE(gen[5794]),

			.O(gen[5887]),
			.E(gen[5889]),

			.SO(gen[5982]),
			.S(gen[5983]),
			.SE(gen[5984]),

			.SELF(gen[5888]),
			.cell_state(gen[5888])
		); 

/******************* CELL 5889 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5889 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5793]),
			.N(gen[5794]),
			.NE(gen[5793]),

			.O(gen[5888]),
			.E(gen[5888]),

			.SO(gen[5983]),
			.S(gen[5984]),
			.SE(gen[5983]),

			.SELF(gen[5889]),
			.cell_state(gen[5889])
		); 

/******************* CELL 5890 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5890 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5796]),
			.N(gen[5795]),
			.NE(gen[5796]),

			.O(gen[5891]),
			.E(gen[5891]),

			.SO(gen[5986]),
			.S(gen[5985]),
			.SE(gen[5986]),

			.SELF(gen[5890]),
			.cell_state(gen[5890])
		); 

/******************* CELL 5891 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5891 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5795]),
			.N(gen[5796]),
			.NE(gen[5797]),

			.O(gen[5890]),
			.E(gen[5892]),

			.SO(gen[5985]),
			.S(gen[5986]),
			.SE(gen[5987]),

			.SELF(gen[5891]),
			.cell_state(gen[5891])
		); 

/******************* CELL 5892 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5892 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5796]),
			.N(gen[5797]),
			.NE(gen[5798]),

			.O(gen[5891]),
			.E(gen[5893]),

			.SO(gen[5986]),
			.S(gen[5987]),
			.SE(gen[5988]),

			.SELF(gen[5892]),
			.cell_state(gen[5892])
		); 

/******************* CELL 5893 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5893 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5797]),
			.N(gen[5798]),
			.NE(gen[5799]),

			.O(gen[5892]),
			.E(gen[5894]),

			.SO(gen[5987]),
			.S(gen[5988]),
			.SE(gen[5989]),

			.SELF(gen[5893]),
			.cell_state(gen[5893])
		); 

/******************* CELL 5894 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5894 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5798]),
			.N(gen[5799]),
			.NE(gen[5800]),

			.O(gen[5893]),
			.E(gen[5895]),

			.SO(gen[5988]),
			.S(gen[5989]),
			.SE(gen[5990]),

			.SELF(gen[5894]),
			.cell_state(gen[5894])
		); 

/******************* CELL 5895 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5895 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5799]),
			.N(gen[5800]),
			.NE(gen[5801]),

			.O(gen[5894]),
			.E(gen[5896]),

			.SO(gen[5989]),
			.S(gen[5990]),
			.SE(gen[5991]),

			.SELF(gen[5895]),
			.cell_state(gen[5895])
		); 

/******************* CELL 5896 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5896 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5800]),
			.N(gen[5801]),
			.NE(gen[5802]),

			.O(gen[5895]),
			.E(gen[5897]),

			.SO(gen[5990]),
			.S(gen[5991]),
			.SE(gen[5992]),

			.SELF(gen[5896]),
			.cell_state(gen[5896])
		); 

/******************* CELL 5897 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5897 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5801]),
			.N(gen[5802]),
			.NE(gen[5803]),

			.O(gen[5896]),
			.E(gen[5898]),

			.SO(gen[5991]),
			.S(gen[5992]),
			.SE(gen[5993]),

			.SELF(gen[5897]),
			.cell_state(gen[5897])
		); 

/******************* CELL 5898 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5898 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5802]),
			.N(gen[5803]),
			.NE(gen[5804]),

			.O(gen[5897]),
			.E(gen[5899]),

			.SO(gen[5992]),
			.S(gen[5993]),
			.SE(gen[5994]),

			.SELF(gen[5898]),
			.cell_state(gen[5898])
		); 

/******************* CELL 5899 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5899 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5803]),
			.N(gen[5804]),
			.NE(gen[5805]),

			.O(gen[5898]),
			.E(gen[5900]),

			.SO(gen[5993]),
			.S(gen[5994]),
			.SE(gen[5995]),

			.SELF(gen[5899]),
			.cell_state(gen[5899])
		); 

/******************* CELL 5900 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5900 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5804]),
			.N(gen[5805]),
			.NE(gen[5806]),

			.O(gen[5899]),
			.E(gen[5901]),

			.SO(gen[5994]),
			.S(gen[5995]),
			.SE(gen[5996]),

			.SELF(gen[5900]),
			.cell_state(gen[5900])
		); 

/******************* CELL 5901 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5901 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5805]),
			.N(gen[5806]),
			.NE(gen[5807]),

			.O(gen[5900]),
			.E(gen[5902]),

			.SO(gen[5995]),
			.S(gen[5996]),
			.SE(gen[5997]),

			.SELF(gen[5901]),
			.cell_state(gen[5901])
		); 

/******************* CELL 5902 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5902 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5806]),
			.N(gen[5807]),
			.NE(gen[5808]),

			.O(gen[5901]),
			.E(gen[5903]),

			.SO(gen[5996]),
			.S(gen[5997]),
			.SE(gen[5998]),

			.SELF(gen[5902]),
			.cell_state(gen[5902])
		); 

/******************* CELL 5903 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5903 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5807]),
			.N(gen[5808]),
			.NE(gen[5809]),

			.O(gen[5902]),
			.E(gen[5904]),

			.SO(gen[5997]),
			.S(gen[5998]),
			.SE(gen[5999]),

			.SELF(gen[5903]),
			.cell_state(gen[5903])
		); 

/******************* CELL 5904 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5904 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5808]),
			.N(gen[5809]),
			.NE(gen[5810]),

			.O(gen[5903]),
			.E(gen[5905]),

			.SO(gen[5998]),
			.S(gen[5999]),
			.SE(gen[6000]),

			.SELF(gen[5904]),
			.cell_state(gen[5904])
		); 

/******************* CELL 5905 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5905 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5809]),
			.N(gen[5810]),
			.NE(gen[5811]),

			.O(gen[5904]),
			.E(gen[5906]),

			.SO(gen[5999]),
			.S(gen[6000]),
			.SE(gen[6001]),

			.SELF(gen[5905]),
			.cell_state(gen[5905])
		); 

/******************* CELL 5906 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5906 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5810]),
			.N(gen[5811]),
			.NE(gen[5812]),

			.O(gen[5905]),
			.E(gen[5907]),

			.SO(gen[6000]),
			.S(gen[6001]),
			.SE(gen[6002]),

			.SELF(gen[5906]),
			.cell_state(gen[5906])
		); 

/******************* CELL 5907 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5907 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5811]),
			.N(gen[5812]),
			.NE(gen[5813]),

			.O(gen[5906]),
			.E(gen[5908]),

			.SO(gen[6001]),
			.S(gen[6002]),
			.SE(gen[6003]),

			.SELF(gen[5907]),
			.cell_state(gen[5907])
		); 

/******************* CELL 5908 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5908 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5812]),
			.N(gen[5813]),
			.NE(gen[5814]),

			.O(gen[5907]),
			.E(gen[5909]),

			.SO(gen[6002]),
			.S(gen[6003]),
			.SE(gen[6004]),

			.SELF(gen[5908]),
			.cell_state(gen[5908])
		); 

/******************* CELL 5909 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5909 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5813]),
			.N(gen[5814]),
			.NE(gen[5815]),

			.O(gen[5908]),
			.E(gen[5910]),

			.SO(gen[6003]),
			.S(gen[6004]),
			.SE(gen[6005]),

			.SELF(gen[5909]),
			.cell_state(gen[5909])
		); 

/******************* CELL 5910 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5910 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5814]),
			.N(gen[5815]),
			.NE(gen[5816]),

			.O(gen[5909]),
			.E(gen[5911]),

			.SO(gen[6004]),
			.S(gen[6005]),
			.SE(gen[6006]),

			.SELF(gen[5910]),
			.cell_state(gen[5910])
		); 

/******************* CELL 5911 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5911 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5815]),
			.N(gen[5816]),
			.NE(gen[5817]),

			.O(gen[5910]),
			.E(gen[5912]),

			.SO(gen[6005]),
			.S(gen[6006]),
			.SE(gen[6007]),

			.SELF(gen[5911]),
			.cell_state(gen[5911])
		); 

/******************* CELL 5912 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5912 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5816]),
			.N(gen[5817]),
			.NE(gen[5818]),

			.O(gen[5911]),
			.E(gen[5913]),

			.SO(gen[6006]),
			.S(gen[6007]),
			.SE(gen[6008]),

			.SELF(gen[5912]),
			.cell_state(gen[5912])
		); 

/******************* CELL 5913 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5913 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5817]),
			.N(gen[5818]),
			.NE(gen[5819]),

			.O(gen[5912]),
			.E(gen[5914]),

			.SO(gen[6007]),
			.S(gen[6008]),
			.SE(gen[6009]),

			.SELF(gen[5913]),
			.cell_state(gen[5913])
		); 

/******************* CELL 5914 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5914 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5818]),
			.N(gen[5819]),
			.NE(gen[5820]),

			.O(gen[5913]),
			.E(gen[5915]),

			.SO(gen[6008]),
			.S(gen[6009]),
			.SE(gen[6010]),

			.SELF(gen[5914]),
			.cell_state(gen[5914])
		); 

/******************* CELL 5915 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5915 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5819]),
			.N(gen[5820]),
			.NE(gen[5821]),

			.O(gen[5914]),
			.E(gen[5916]),

			.SO(gen[6009]),
			.S(gen[6010]),
			.SE(gen[6011]),

			.SELF(gen[5915]),
			.cell_state(gen[5915])
		); 

/******************* CELL 5916 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5916 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5820]),
			.N(gen[5821]),
			.NE(gen[5822]),

			.O(gen[5915]),
			.E(gen[5917]),

			.SO(gen[6010]),
			.S(gen[6011]),
			.SE(gen[6012]),

			.SELF(gen[5916]),
			.cell_state(gen[5916])
		); 

/******************* CELL 5917 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5917 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5821]),
			.N(gen[5822]),
			.NE(gen[5823]),

			.O(gen[5916]),
			.E(gen[5918]),

			.SO(gen[6011]),
			.S(gen[6012]),
			.SE(gen[6013]),

			.SELF(gen[5917]),
			.cell_state(gen[5917])
		); 

/******************* CELL 5918 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5918 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5822]),
			.N(gen[5823]),
			.NE(gen[5824]),

			.O(gen[5917]),
			.E(gen[5919]),

			.SO(gen[6012]),
			.S(gen[6013]),
			.SE(gen[6014]),

			.SELF(gen[5918]),
			.cell_state(gen[5918])
		); 

/******************* CELL 5919 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5919 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5823]),
			.N(gen[5824]),
			.NE(gen[5825]),

			.O(gen[5918]),
			.E(gen[5920]),

			.SO(gen[6013]),
			.S(gen[6014]),
			.SE(gen[6015]),

			.SELF(gen[5919]),
			.cell_state(gen[5919])
		); 

/******************* CELL 5920 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5920 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5824]),
			.N(gen[5825]),
			.NE(gen[5826]),

			.O(gen[5919]),
			.E(gen[5921]),

			.SO(gen[6014]),
			.S(gen[6015]),
			.SE(gen[6016]),

			.SELF(gen[5920]),
			.cell_state(gen[5920])
		); 

/******************* CELL 5921 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5921 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5825]),
			.N(gen[5826]),
			.NE(gen[5827]),

			.O(gen[5920]),
			.E(gen[5922]),

			.SO(gen[6015]),
			.S(gen[6016]),
			.SE(gen[6017]),

			.SELF(gen[5921]),
			.cell_state(gen[5921])
		); 

/******************* CELL 5922 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5922 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5826]),
			.N(gen[5827]),
			.NE(gen[5828]),

			.O(gen[5921]),
			.E(gen[5923]),

			.SO(gen[6016]),
			.S(gen[6017]),
			.SE(gen[6018]),

			.SELF(gen[5922]),
			.cell_state(gen[5922])
		); 

/******************* CELL 5923 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5923 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5827]),
			.N(gen[5828]),
			.NE(gen[5829]),

			.O(gen[5922]),
			.E(gen[5924]),

			.SO(gen[6017]),
			.S(gen[6018]),
			.SE(gen[6019]),

			.SELF(gen[5923]),
			.cell_state(gen[5923])
		); 

/******************* CELL 5924 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5924 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5828]),
			.N(gen[5829]),
			.NE(gen[5830]),

			.O(gen[5923]),
			.E(gen[5925]),

			.SO(gen[6018]),
			.S(gen[6019]),
			.SE(gen[6020]),

			.SELF(gen[5924]),
			.cell_state(gen[5924])
		); 

/******************* CELL 5925 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5925 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5829]),
			.N(gen[5830]),
			.NE(gen[5831]),

			.O(gen[5924]),
			.E(gen[5926]),

			.SO(gen[6019]),
			.S(gen[6020]),
			.SE(gen[6021]),

			.SELF(gen[5925]),
			.cell_state(gen[5925])
		); 

/******************* CELL 5926 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5926 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5830]),
			.N(gen[5831]),
			.NE(gen[5832]),

			.O(gen[5925]),
			.E(gen[5927]),

			.SO(gen[6020]),
			.S(gen[6021]),
			.SE(gen[6022]),

			.SELF(gen[5926]),
			.cell_state(gen[5926])
		); 

/******************* CELL 5927 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5927 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5831]),
			.N(gen[5832]),
			.NE(gen[5833]),

			.O(gen[5926]),
			.E(gen[5928]),

			.SO(gen[6021]),
			.S(gen[6022]),
			.SE(gen[6023]),

			.SELF(gen[5927]),
			.cell_state(gen[5927])
		); 

/******************* CELL 5928 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5928 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5832]),
			.N(gen[5833]),
			.NE(gen[5834]),

			.O(gen[5927]),
			.E(gen[5929]),

			.SO(gen[6022]),
			.S(gen[6023]),
			.SE(gen[6024]),

			.SELF(gen[5928]),
			.cell_state(gen[5928])
		); 

/******************* CELL 5929 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5929 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5833]),
			.N(gen[5834]),
			.NE(gen[5835]),

			.O(gen[5928]),
			.E(gen[5930]),

			.SO(gen[6023]),
			.S(gen[6024]),
			.SE(gen[6025]),

			.SELF(gen[5929]),
			.cell_state(gen[5929])
		); 

/******************* CELL 5930 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5930 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5834]),
			.N(gen[5835]),
			.NE(gen[5836]),

			.O(gen[5929]),
			.E(gen[5931]),

			.SO(gen[6024]),
			.S(gen[6025]),
			.SE(gen[6026]),

			.SELF(gen[5930]),
			.cell_state(gen[5930])
		); 

/******************* CELL 5931 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5931 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5835]),
			.N(gen[5836]),
			.NE(gen[5837]),

			.O(gen[5930]),
			.E(gen[5932]),

			.SO(gen[6025]),
			.S(gen[6026]),
			.SE(gen[6027]),

			.SELF(gen[5931]),
			.cell_state(gen[5931])
		); 

/******************* CELL 5932 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5932 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5836]),
			.N(gen[5837]),
			.NE(gen[5838]),

			.O(gen[5931]),
			.E(gen[5933]),

			.SO(gen[6026]),
			.S(gen[6027]),
			.SE(gen[6028]),

			.SELF(gen[5932]),
			.cell_state(gen[5932])
		); 

/******************* CELL 5933 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5933 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5837]),
			.N(gen[5838]),
			.NE(gen[5839]),

			.O(gen[5932]),
			.E(gen[5934]),

			.SO(gen[6027]),
			.S(gen[6028]),
			.SE(gen[6029]),

			.SELF(gen[5933]),
			.cell_state(gen[5933])
		); 

/******************* CELL 5934 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5934 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5838]),
			.N(gen[5839]),
			.NE(gen[5840]),

			.O(gen[5933]),
			.E(gen[5935]),

			.SO(gen[6028]),
			.S(gen[6029]),
			.SE(gen[6030]),

			.SELF(gen[5934]),
			.cell_state(gen[5934])
		); 

/******************* CELL 5935 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5935 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5839]),
			.N(gen[5840]),
			.NE(gen[5841]),

			.O(gen[5934]),
			.E(gen[5936]),

			.SO(gen[6029]),
			.S(gen[6030]),
			.SE(gen[6031]),

			.SELF(gen[5935]),
			.cell_state(gen[5935])
		); 

/******************* CELL 5936 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5936 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5840]),
			.N(gen[5841]),
			.NE(gen[5842]),

			.O(gen[5935]),
			.E(gen[5937]),

			.SO(gen[6030]),
			.S(gen[6031]),
			.SE(gen[6032]),

			.SELF(gen[5936]),
			.cell_state(gen[5936])
		); 

/******************* CELL 5937 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5937 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5841]),
			.N(gen[5842]),
			.NE(gen[5843]),

			.O(gen[5936]),
			.E(gen[5938]),

			.SO(gen[6031]),
			.S(gen[6032]),
			.SE(gen[6033]),

			.SELF(gen[5937]),
			.cell_state(gen[5937])
		); 

/******************* CELL 5938 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5938 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5842]),
			.N(gen[5843]),
			.NE(gen[5844]),

			.O(gen[5937]),
			.E(gen[5939]),

			.SO(gen[6032]),
			.S(gen[6033]),
			.SE(gen[6034]),

			.SELF(gen[5938]),
			.cell_state(gen[5938])
		); 

/******************* CELL 5939 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5939 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5843]),
			.N(gen[5844]),
			.NE(gen[5845]),

			.O(gen[5938]),
			.E(gen[5940]),

			.SO(gen[6033]),
			.S(gen[6034]),
			.SE(gen[6035]),

			.SELF(gen[5939]),
			.cell_state(gen[5939])
		); 

/******************* CELL 5940 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5940 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5844]),
			.N(gen[5845]),
			.NE(gen[5846]),

			.O(gen[5939]),
			.E(gen[5941]),

			.SO(gen[6034]),
			.S(gen[6035]),
			.SE(gen[6036]),

			.SELF(gen[5940]),
			.cell_state(gen[5940])
		); 

/******************* CELL 5941 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5941 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5845]),
			.N(gen[5846]),
			.NE(gen[5847]),

			.O(gen[5940]),
			.E(gen[5942]),

			.SO(gen[6035]),
			.S(gen[6036]),
			.SE(gen[6037]),

			.SELF(gen[5941]),
			.cell_state(gen[5941])
		); 

/******************* CELL 5942 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5942 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5846]),
			.N(gen[5847]),
			.NE(gen[5848]),

			.O(gen[5941]),
			.E(gen[5943]),

			.SO(gen[6036]),
			.S(gen[6037]),
			.SE(gen[6038]),

			.SELF(gen[5942]),
			.cell_state(gen[5942])
		); 

/******************* CELL 5943 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5943 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5847]),
			.N(gen[5848]),
			.NE(gen[5849]),

			.O(gen[5942]),
			.E(gen[5944]),

			.SO(gen[6037]),
			.S(gen[6038]),
			.SE(gen[6039]),

			.SELF(gen[5943]),
			.cell_state(gen[5943])
		); 

/******************* CELL 5944 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5944 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5848]),
			.N(gen[5849]),
			.NE(gen[5850]),

			.O(gen[5943]),
			.E(gen[5945]),

			.SO(gen[6038]),
			.S(gen[6039]),
			.SE(gen[6040]),

			.SELF(gen[5944]),
			.cell_state(gen[5944])
		); 

/******************* CELL 5945 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5945 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5849]),
			.N(gen[5850]),
			.NE(gen[5851]),

			.O(gen[5944]),
			.E(gen[5946]),

			.SO(gen[6039]),
			.S(gen[6040]),
			.SE(gen[6041]),

			.SELF(gen[5945]),
			.cell_state(gen[5945])
		); 

/******************* CELL 5946 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5946 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5850]),
			.N(gen[5851]),
			.NE(gen[5852]),

			.O(gen[5945]),
			.E(gen[5947]),

			.SO(gen[6040]),
			.S(gen[6041]),
			.SE(gen[6042]),

			.SELF(gen[5946]),
			.cell_state(gen[5946])
		); 

/******************* CELL 5947 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5947 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5851]),
			.N(gen[5852]),
			.NE(gen[5853]),

			.O(gen[5946]),
			.E(gen[5948]),

			.SO(gen[6041]),
			.S(gen[6042]),
			.SE(gen[6043]),

			.SELF(gen[5947]),
			.cell_state(gen[5947])
		); 

/******************* CELL 5948 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5948 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5852]),
			.N(gen[5853]),
			.NE(gen[5854]),

			.O(gen[5947]),
			.E(gen[5949]),

			.SO(gen[6042]),
			.S(gen[6043]),
			.SE(gen[6044]),

			.SELF(gen[5948]),
			.cell_state(gen[5948])
		); 

/******************* CELL 5949 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5949 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5853]),
			.N(gen[5854]),
			.NE(gen[5855]),

			.O(gen[5948]),
			.E(gen[5950]),

			.SO(gen[6043]),
			.S(gen[6044]),
			.SE(gen[6045]),

			.SELF(gen[5949]),
			.cell_state(gen[5949])
		); 

/******************* CELL 5950 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5950 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5854]),
			.N(gen[5855]),
			.NE(gen[5856]),

			.O(gen[5949]),
			.E(gen[5951]),

			.SO(gen[6044]),
			.S(gen[6045]),
			.SE(gen[6046]),

			.SELF(gen[5950]),
			.cell_state(gen[5950])
		); 

/******************* CELL 5951 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5951 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5855]),
			.N(gen[5856]),
			.NE(gen[5857]),

			.O(gen[5950]),
			.E(gen[5952]),

			.SO(gen[6045]),
			.S(gen[6046]),
			.SE(gen[6047]),

			.SELF(gen[5951]),
			.cell_state(gen[5951])
		); 

/******************* CELL 5952 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5952 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5856]),
			.N(gen[5857]),
			.NE(gen[5858]),

			.O(gen[5951]),
			.E(gen[5953]),

			.SO(gen[6046]),
			.S(gen[6047]),
			.SE(gen[6048]),

			.SELF(gen[5952]),
			.cell_state(gen[5952])
		); 

/******************* CELL 5953 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5953 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5857]),
			.N(gen[5858]),
			.NE(gen[5859]),

			.O(gen[5952]),
			.E(gen[5954]),

			.SO(gen[6047]),
			.S(gen[6048]),
			.SE(gen[6049]),

			.SELF(gen[5953]),
			.cell_state(gen[5953])
		); 

/******************* CELL 5954 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5954 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5858]),
			.N(gen[5859]),
			.NE(gen[5860]),

			.O(gen[5953]),
			.E(gen[5955]),

			.SO(gen[6048]),
			.S(gen[6049]),
			.SE(gen[6050]),

			.SELF(gen[5954]),
			.cell_state(gen[5954])
		); 

/******************* CELL 5955 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5955 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5859]),
			.N(gen[5860]),
			.NE(gen[5861]),

			.O(gen[5954]),
			.E(gen[5956]),

			.SO(gen[6049]),
			.S(gen[6050]),
			.SE(gen[6051]),

			.SELF(gen[5955]),
			.cell_state(gen[5955])
		); 

/******************* CELL 5956 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5956 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5860]),
			.N(gen[5861]),
			.NE(gen[5862]),

			.O(gen[5955]),
			.E(gen[5957]),

			.SO(gen[6050]),
			.S(gen[6051]),
			.SE(gen[6052]),

			.SELF(gen[5956]),
			.cell_state(gen[5956])
		); 

/******************* CELL 5957 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5957 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5861]),
			.N(gen[5862]),
			.NE(gen[5863]),

			.O(gen[5956]),
			.E(gen[5958]),

			.SO(gen[6051]),
			.S(gen[6052]),
			.SE(gen[6053]),

			.SELF(gen[5957]),
			.cell_state(gen[5957])
		); 

/******************* CELL 5958 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5958 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5862]),
			.N(gen[5863]),
			.NE(gen[5864]),

			.O(gen[5957]),
			.E(gen[5959]),

			.SO(gen[6052]),
			.S(gen[6053]),
			.SE(gen[6054]),

			.SELF(gen[5958]),
			.cell_state(gen[5958])
		); 

/******************* CELL 5959 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5959 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5863]),
			.N(gen[5864]),
			.NE(gen[5865]),

			.O(gen[5958]),
			.E(gen[5960]),

			.SO(gen[6053]),
			.S(gen[6054]),
			.SE(gen[6055]),

			.SELF(gen[5959]),
			.cell_state(gen[5959])
		); 

/******************* CELL 5960 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5960 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5864]),
			.N(gen[5865]),
			.NE(gen[5866]),

			.O(gen[5959]),
			.E(gen[5961]),

			.SO(gen[6054]),
			.S(gen[6055]),
			.SE(gen[6056]),

			.SELF(gen[5960]),
			.cell_state(gen[5960])
		); 

/******************* CELL 5961 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5961 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5865]),
			.N(gen[5866]),
			.NE(gen[5867]),

			.O(gen[5960]),
			.E(gen[5962]),

			.SO(gen[6055]),
			.S(gen[6056]),
			.SE(gen[6057]),

			.SELF(gen[5961]),
			.cell_state(gen[5961])
		); 

/******************* CELL 5962 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5962 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5866]),
			.N(gen[5867]),
			.NE(gen[5868]),

			.O(gen[5961]),
			.E(gen[5963]),

			.SO(gen[6056]),
			.S(gen[6057]),
			.SE(gen[6058]),

			.SELF(gen[5962]),
			.cell_state(gen[5962])
		); 

/******************* CELL 5963 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5963 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5867]),
			.N(gen[5868]),
			.NE(gen[5869]),

			.O(gen[5962]),
			.E(gen[5964]),

			.SO(gen[6057]),
			.S(gen[6058]),
			.SE(gen[6059]),

			.SELF(gen[5963]),
			.cell_state(gen[5963])
		); 

/******************* CELL 5964 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5964 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5868]),
			.N(gen[5869]),
			.NE(gen[5870]),

			.O(gen[5963]),
			.E(gen[5965]),

			.SO(gen[6058]),
			.S(gen[6059]),
			.SE(gen[6060]),

			.SELF(gen[5964]),
			.cell_state(gen[5964])
		); 

/******************* CELL 5965 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5965 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5869]),
			.N(gen[5870]),
			.NE(gen[5871]),

			.O(gen[5964]),
			.E(gen[5966]),

			.SO(gen[6059]),
			.S(gen[6060]),
			.SE(gen[6061]),

			.SELF(gen[5965]),
			.cell_state(gen[5965])
		); 

/******************* CELL 5966 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5966 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5870]),
			.N(gen[5871]),
			.NE(gen[5872]),

			.O(gen[5965]),
			.E(gen[5967]),

			.SO(gen[6060]),
			.S(gen[6061]),
			.SE(gen[6062]),

			.SELF(gen[5966]),
			.cell_state(gen[5966])
		); 

/******************* CELL 5967 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5967 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5871]),
			.N(gen[5872]),
			.NE(gen[5873]),

			.O(gen[5966]),
			.E(gen[5968]),

			.SO(gen[6061]),
			.S(gen[6062]),
			.SE(gen[6063]),

			.SELF(gen[5967]),
			.cell_state(gen[5967])
		); 

/******************* CELL 5968 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5968 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5872]),
			.N(gen[5873]),
			.NE(gen[5874]),

			.O(gen[5967]),
			.E(gen[5969]),

			.SO(gen[6062]),
			.S(gen[6063]),
			.SE(gen[6064]),

			.SELF(gen[5968]),
			.cell_state(gen[5968])
		); 

/******************* CELL 5969 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5969 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5873]),
			.N(gen[5874]),
			.NE(gen[5875]),

			.O(gen[5968]),
			.E(gen[5970]),

			.SO(gen[6063]),
			.S(gen[6064]),
			.SE(gen[6065]),

			.SELF(gen[5969]),
			.cell_state(gen[5969])
		); 

/******************* CELL 5970 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5970 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5874]),
			.N(gen[5875]),
			.NE(gen[5876]),

			.O(gen[5969]),
			.E(gen[5971]),

			.SO(gen[6064]),
			.S(gen[6065]),
			.SE(gen[6066]),

			.SELF(gen[5970]),
			.cell_state(gen[5970])
		); 

/******************* CELL 5971 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5971 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5875]),
			.N(gen[5876]),
			.NE(gen[5877]),

			.O(gen[5970]),
			.E(gen[5972]),

			.SO(gen[6065]),
			.S(gen[6066]),
			.SE(gen[6067]),

			.SELF(gen[5971]),
			.cell_state(gen[5971])
		); 

/******************* CELL 5972 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5972 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5876]),
			.N(gen[5877]),
			.NE(gen[5878]),

			.O(gen[5971]),
			.E(gen[5973]),

			.SO(gen[6066]),
			.S(gen[6067]),
			.SE(gen[6068]),

			.SELF(gen[5972]),
			.cell_state(gen[5972])
		); 

/******************* CELL 5973 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5973 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5877]),
			.N(gen[5878]),
			.NE(gen[5879]),

			.O(gen[5972]),
			.E(gen[5974]),

			.SO(gen[6067]),
			.S(gen[6068]),
			.SE(gen[6069]),

			.SELF(gen[5973]),
			.cell_state(gen[5973])
		); 

/******************* CELL 5974 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5974 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5878]),
			.N(gen[5879]),
			.NE(gen[5880]),

			.O(gen[5973]),
			.E(gen[5975]),

			.SO(gen[6068]),
			.S(gen[6069]),
			.SE(gen[6070]),

			.SELF(gen[5974]),
			.cell_state(gen[5974])
		); 

/******************* CELL 5975 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5975 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5879]),
			.N(gen[5880]),
			.NE(gen[5881]),

			.O(gen[5974]),
			.E(gen[5976]),

			.SO(gen[6069]),
			.S(gen[6070]),
			.SE(gen[6071]),

			.SELF(gen[5975]),
			.cell_state(gen[5975])
		); 

/******************* CELL 5976 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5976 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5880]),
			.N(gen[5881]),
			.NE(gen[5882]),

			.O(gen[5975]),
			.E(gen[5977]),

			.SO(gen[6070]),
			.S(gen[6071]),
			.SE(gen[6072]),

			.SELF(gen[5976]),
			.cell_state(gen[5976])
		); 

/******************* CELL 5977 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5977 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5881]),
			.N(gen[5882]),
			.NE(gen[5883]),

			.O(gen[5976]),
			.E(gen[5978]),

			.SO(gen[6071]),
			.S(gen[6072]),
			.SE(gen[6073]),

			.SELF(gen[5977]),
			.cell_state(gen[5977])
		); 

/******************* CELL 5978 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5978 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5882]),
			.N(gen[5883]),
			.NE(gen[5884]),

			.O(gen[5977]),
			.E(gen[5979]),

			.SO(gen[6072]),
			.S(gen[6073]),
			.SE(gen[6074]),

			.SELF(gen[5978]),
			.cell_state(gen[5978])
		); 

/******************* CELL 5979 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5979 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5883]),
			.N(gen[5884]),
			.NE(gen[5885]),

			.O(gen[5978]),
			.E(gen[5980]),

			.SO(gen[6073]),
			.S(gen[6074]),
			.SE(gen[6075]),

			.SELF(gen[5979]),
			.cell_state(gen[5979])
		); 

/******************* CELL 5980 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5980 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5884]),
			.N(gen[5885]),
			.NE(gen[5886]),

			.O(gen[5979]),
			.E(gen[5981]),

			.SO(gen[6074]),
			.S(gen[6075]),
			.SE(gen[6076]),

			.SELF(gen[5980]),
			.cell_state(gen[5980])
		); 

/******************* CELL 5981 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5981 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5885]),
			.N(gen[5886]),
			.NE(gen[5887]),

			.O(gen[5980]),
			.E(gen[5982]),

			.SO(gen[6075]),
			.S(gen[6076]),
			.SE(gen[6077]),

			.SELF(gen[5981]),
			.cell_state(gen[5981])
		); 

/******************* CELL 5982 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5982 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5886]),
			.N(gen[5887]),
			.NE(gen[5888]),

			.O(gen[5981]),
			.E(gen[5983]),

			.SO(gen[6076]),
			.S(gen[6077]),
			.SE(gen[6078]),

			.SELF(gen[5982]),
			.cell_state(gen[5982])
		); 

/******************* CELL 5983 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5983 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5887]),
			.N(gen[5888]),
			.NE(gen[5889]),

			.O(gen[5982]),
			.E(gen[5984]),

			.SO(gen[6077]),
			.S(gen[6078]),
			.SE(gen[6079]),

			.SELF(gen[5983]),
			.cell_state(gen[5983])
		); 

/******************* CELL 5984 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5984 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5888]),
			.N(gen[5889]),
			.NE(gen[5888]),

			.O(gen[5983]),
			.E(gen[5983]),

			.SO(gen[6078]),
			.S(gen[6079]),
			.SE(gen[6078]),

			.SELF(gen[5984]),
			.cell_state(gen[5984])
		); 

/******************* CELL 5985 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5985 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5891]),
			.N(gen[5890]),
			.NE(gen[5891]),

			.O(gen[5986]),
			.E(gen[5986]),

			.SO(gen[6081]),
			.S(gen[6080]),
			.SE(gen[6081]),

			.SELF(gen[5985]),
			.cell_state(gen[5985])
		); 

/******************* CELL 5986 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5986 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5890]),
			.N(gen[5891]),
			.NE(gen[5892]),

			.O(gen[5985]),
			.E(gen[5987]),

			.SO(gen[6080]),
			.S(gen[6081]),
			.SE(gen[6082]),

			.SELF(gen[5986]),
			.cell_state(gen[5986])
		); 

/******************* CELL 5987 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5987 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5891]),
			.N(gen[5892]),
			.NE(gen[5893]),

			.O(gen[5986]),
			.E(gen[5988]),

			.SO(gen[6081]),
			.S(gen[6082]),
			.SE(gen[6083]),

			.SELF(gen[5987]),
			.cell_state(gen[5987])
		); 

/******************* CELL 5988 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5988 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5892]),
			.N(gen[5893]),
			.NE(gen[5894]),

			.O(gen[5987]),
			.E(gen[5989]),

			.SO(gen[6082]),
			.S(gen[6083]),
			.SE(gen[6084]),

			.SELF(gen[5988]),
			.cell_state(gen[5988])
		); 

/******************* CELL 5989 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5989 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5893]),
			.N(gen[5894]),
			.NE(gen[5895]),

			.O(gen[5988]),
			.E(gen[5990]),

			.SO(gen[6083]),
			.S(gen[6084]),
			.SE(gen[6085]),

			.SELF(gen[5989]),
			.cell_state(gen[5989])
		); 

/******************* CELL 5990 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5990 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5894]),
			.N(gen[5895]),
			.NE(gen[5896]),

			.O(gen[5989]),
			.E(gen[5991]),

			.SO(gen[6084]),
			.S(gen[6085]),
			.SE(gen[6086]),

			.SELF(gen[5990]),
			.cell_state(gen[5990])
		); 

/******************* CELL 5991 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5991 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5895]),
			.N(gen[5896]),
			.NE(gen[5897]),

			.O(gen[5990]),
			.E(gen[5992]),

			.SO(gen[6085]),
			.S(gen[6086]),
			.SE(gen[6087]),

			.SELF(gen[5991]),
			.cell_state(gen[5991])
		); 

/******************* CELL 5992 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5992 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5896]),
			.N(gen[5897]),
			.NE(gen[5898]),

			.O(gen[5991]),
			.E(gen[5993]),

			.SO(gen[6086]),
			.S(gen[6087]),
			.SE(gen[6088]),

			.SELF(gen[5992]),
			.cell_state(gen[5992])
		); 

/******************* CELL 5993 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5993 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5897]),
			.N(gen[5898]),
			.NE(gen[5899]),

			.O(gen[5992]),
			.E(gen[5994]),

			.SO(gen[6087]),
			.S(gen[6088]),
			.SE(gen[6089]),

			.SELF(gen[5993]),
			.cell_state(gen[5993])
		); 

/******************* CELL 5994 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5994 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5898]),
			.N(gen[5899]),
			.NE(gen[5900]),

			.O(gen[5993]),
			.E(gen[5995]),

			.SO(gen[6088]),
			.S(gen[6089]),
			.SE(gen[6090]),

			.SELF(gen[5994]),
			.cell_state(gen[5994])
		); 

/******************* CELL 5995 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5995 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5899]),
			.N(gen[5900]),
			.NE(gen[5901]),

			.O(gen[5994]),
			.E(gen[5996]),

			.SO(gen[6089]),
			.S(gen[6090]),
			.SE(gen[6091]),

			.SELF(gen[5995]),
			.cell_state(gen[5995])
		); 

/******************* CELL 5996 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5996 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5900]),
			.N(gen[5901]),
			.NE(gen[5902]),

			.O(gen[5995]),
			.E(gen[5997]),

			.SO(gen[6090]),
			.S(gen[6091]),
			.SE(gen[6092]),

			.SELF(gen[5996]),
			.cell_state(gen[5996])
		); 

/******************* CELL 5997 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5997 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5901]),
			.N(gen[5902]),
			.NE(gen[5903]),

			.O(gen[5996]),
			.E(gen[5998]),

			.SO(gen[6091]),
			.S(gen[6092]),
			.SE(gen[6093]),

			.SELF(gen[5997]),
			.cell_state(gen[5997])
		); 

/******************* CELL 5998 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5998 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5902]),
			.N(gen[5903]),
			.NE(gen[5904]),

			.O(gen[5997]),
			.E(gen[5999]),

			.SO(gen[6092]),
			.S(gen[6093]),
			.SE(gen[6094]),

			.SELF(gen[5998]),
			.cell_state(gen[5998])
		); 

/******************* CELL 5999 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell5999 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5903]),
			.N(gen[5904]),
			.NE(gen[5905]),

			.O(gen[5998]),
			.E(gen[6000]),

			.SO(gen[6093]),
			.S(gen[6094]),
			.SE(gen[6095]),

			.SELF(gen[5999]),
			.cell_state(gen[5999])
		); 

/******************* CELL 6000 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6000 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5904]),
			.N(gen[5905]),
			.NE(gen[5906]),

			.O(gen[5999]),
			.E(gen[6001]),

			.SO(gen[6094]),
			.S(gen[6095]),
			.SE(gen[6096]),

			.SELF(gen[6000]),
			.cell_state(gen[6000])
		); 

/******************* CELL 6001 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6001 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5905]),
			.N(gen[5906]),
			.NE(gen[5907]),

			.O(gen[6000]),
			.E(gen[6002]),

			.SO(gen[6095]),
			.S(gen[6096]),
			.SE(gen[6097]),

			.SELF(gen[6001]),
			.cell_state(gen[6001])
		); 

/******************* CELL 6002 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6002 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5906]),
			.N(gen[5907]),
			.NE(gen[5908]),

			.O(gen[6001]),
			.E(gen[6003]),

			.SO(gen[6096]),
			.S(gen[6097]),
			.SE(gen[6098]),

			.SELF(gen[6002]),
			.cell_state(gen[6002])
		); 

/******************* CELL 6003 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6003 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5907]),
			.N(gen[5908]),
			.NE(gen[5909]),

			.O(gen[6002]),
			.E(gen[6004]),

			.SO(gen[6097]),
			.S(gen[6098]),
			.SE(gen[6099]),

			.SELF(gen[6003]),
			.cell_state(gen[6003])
		); 

/******************* CELL 6004 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6004 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5908]),
			.N(gen[5909]),
			.NE(gen[5910]),

			.O(gen[6003]),
			.E(gen[6005]),

			.SO(gen[6098]),
			.S(gen[6099]),
			.SE(gen[6100]),

			.SELF(gen[6004]),
			.cell_state(gen[6004])
		); 

/******************* CELL 6005 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6005 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5909]),
			.N(gen[5910]),
			.NE(gen[5911]),

			.O(gen[6004]),
			.E(gen[6006]),

			.SO(gen[6099]),
			.S(gen[6100]),
			.SE(gen[6101]),

			.SELF(gen[6005]),
			.cell_state(gen[6005])
		); 

/******************* CELL 6006 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6006 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5910]),
			.N(gen[5911]),
			.NE(gen[5912]),

			.O(gen[6005]),
			.E(gen[6007]),

			.SO(gen[6100]),
			.S(gen[6101]),
			.SE(gen[6102]),

			.SELF(gen[6006]),
			.cell_state(gen[6006])
		); 

/******************* CELL 6007 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6007 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5911]),
			.N(gen[5912]),
			.NE(gen[5913]),

			.O(gen[6006]),
			.E(gen[6008]),

			.SO(gen[6101]),
			.S(gen[6102]),
			.SE(gen[6103]),

			.SELF(gen[6007]),
			.cell_state(gen[6007])
		); 

/******************* CELL 6008 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6008 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5912]),
			.N(gen[5913]),
			.NE(gen[5914]),

			.O(gen[6007]),
			.E(gen[6009]),

			.SO(gen[6102]),
			.S(gen[6103]),
			.SE(gen[6104]),

			.SELF(gen[6008]),
			.cell_state(gen[6008])
		); 

/******************* CELL 6009 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6009 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5913]),
			.N(gen[5914]),
			.NE(gen[5915]),

			.O(gen[6008]),
			.E(gen[6010]),

			.SO(gen[6103]),
			.S(gen[6104]),
			.SE(gen[6105]),

			.SELF(gen[6009]),
			.cell_state(gen[6009])
		); 

/******************* CELL 6010 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6010 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5914]),
			.N(gen[5915]),
			.NE(gen[5916]),

			.O(gen[6009]),
			.E(gen[6011]),

			.SO(gen[6104]),
			.S(gen[6105]),
			.SE(gen[6106]),

			.SELF(gen[6010]),
			.cell_state(gen[6010])
		); 

/******************* CELL 6011 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6011 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5915]),
			.N(gen[5916]),
			.NE(gen[5917]),

			.O(gen[6010]),
			.E(gen[6012]),

			.SO(gen[6105]),
			.S(gen[6106]),
			.SE(gen[6107]),

			.SELF(gen[6011]),
			.cell_state(gen[6011])
		); 

/******************* CELL 6012 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6012 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5916]),
			.N(gen[5917]),
			.NE(gen[5918]),

			.O(gen[6011]),
			.E(gen[6013]),

			.SO(gen[6106]),
			.S(gen[6107]),
			.SE(gen[6108]),

			.SELF(gen[6012]),
			.cell_state(gen[6012])
		); 

/******************* CELL 6013 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6013 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5917]),
			.N(gen[5918]),
			.NE(gen[5919]),

			.O(gen[6012]),
			.E(gen[6014]),

			.SO(gen[6107]),
			.S(gen[6108]),
			.SE(gen[6109]),

			.SELF(gen[6013]),
			.cell_state(gen[6013])
		); 

/******************* CELL 6014 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6014 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5918]),
			.N(gen[5919]),
			.NE(gen[5920]),

			.O(gen[6013]),
			.E(gen[6015]),

			.SO(gen[6108]),
			.S(gen[6109]),
			.SE(gen[6110]),

			.SELF(gen[6014]),
			.cell_state(gen[6014])
		); 

/******************* CELL 6015 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6015 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5919]),
			.N(gen[5920]),
			.NE(gen[5921]),

			.O(gen[6014]),
			.E(gen[6016]),

			.SO(gen[6109]),
			.S(gen[6110]),
			.SE(gen[6111]),

			.SELF(gen[6015]),
			.cell_state(gen[6015])
		); 

/******************* CELL 6016 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6016 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5920]),
			.N(gen[5921]),
			.NE(gen[5922]),

			.O(gen[6015]),
			.E(gen[6017]),

			.SO(gen[6110]),
			.S(gen[6111]),
			.SE(gen[6112]),

			.SELF(gen[6016]),
			.cell_state(gen[6016])
		); 

/******************* CELL 6017 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6017 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5921]),
			.N(gen[5922]),
			.NE(gen[5923]),

			.O(gen[6016]),
			.E(gen[6018]),

			.SO(gen[6111]),
			.S(gen[6112]),
			.SE(gen[6113]),

			.SELF(gen[6017]),
			.cell_state(gen[6017])
		); 

/******************* CELL 6018 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6018 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5922]),
			.N(gen[5923]),
			.NE(gen[5924]),

			.O(gen[6017]),
			.E(gen[6019]),

			.SO(gen[6112]),
			.S(gen[6113]),
			.SE(gen[6114]),

			.SELF(gen[6018]),
			.cell_state(gen[6018])
		); 

/******************* CELL 6019 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6019 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5923]),
			.N(gen[5924]),
			.NE(gen[5925]),

			.O(gen[6018]),
			.E(gen[6020]),

			.SO(gen[6113]),
			.S(gen[6114]),
			.SE(gen[6115]),

			.SELF(gen[6019]),
			.cell_state(gen[6019])
		); 

/******************* CELL 6020 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6020 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5924]),
			.N(gen[5925]),
			.NE(gen[5926]),

			.O(gen[6019]),
			.E(gen[6021]),

			.SO(gen[6114]),
			.S(gen[6115]),
			.SE(gen[6116]),

			.SELF(gen[6020]),
			.cell_state(gen[6020])
		); 

/******************* CELL 6021 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6021 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5925]),
			.N(gen[5926]),
			.NE(gen[5927]),

			.O(gen[6020]),
			.E(gen[6022]),

			.SO(gen[6115]),
			.S(gen[6116]),
			.SE(gen[6117]),

			.SELF(gen[6021]),
			.cell_state(gen[6021])
		); 

/******************* CELL 6022 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6022 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5926]),
			.N(gen[5927]),
			.NE(gen[5928]),

			.O(gen[6021]),
			.E(gen[6023]),

			.SO(gen[6116]),
			.S(gen[6117]),
			.SE(gen[6118]),

			.SELF(gen[6022]),
			.cell_state(gen[6022])
		); 

/******************* CELL 6023 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6023 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5927]),
			.N(gen[5928]),
			.NE(gen[5929]),

			.O(gen[6022]),
			.E(gen[6024]),

			.SO(gen[6117]),
			.S(gen[6118]),
			.SE(gen[6119]),

			.SELF(gen[6023]),
			.cell_state(gen[6023])
		); 

/******************* CELL 6024 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6024 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5928]),
			.N(gen[5929]),
			.NE(gen[5930]),

			.O(gen[6023]),
			.E(gen[6025]),

			.SO(gen[6118]),
			.S(gen[6119]),
			.SE(gen[6120]),

			.SELF(gen[6024]),
			.cell_state(gen[6024])
		); 

/******************* CELL 6025 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6025 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5929]),
			.N(gen[5930]),
			.NE(gen[5931]),

			.O(gen[6024]),
			.E(gen[6026]),

			.SO(gen[6119]),
			.S(gen[6120]),
			.SE(gen[6121]),

			.SELF(gen[6025]),
			.cell_state(gen[6025])
		); 

/******************* CELL 6026 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6026 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5930]),
			.N(gen[5931]),
			.NE(gen[5932]),

			.O(gen[6025]),
			.E(gen[6027]),

			.SO(gen[6120]),
			.S(gen[6121]),
			.SE(gen[6122]),

			.SELF(gen[6026]),
			.cell_state(gen[6026])
		); 

/******************* CELL 6027 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6027 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5931]),
			.N(gen[5932]),
			.NE(gen[5933]),

			.O(gen[6026]),
			.E(gen[6028]),

			.SO(gen[6121]),
			.S(gen[6122]),
			.SE(gen[6123]),

			.SELF(gen[6027]),
			.cell_state(gen[6027])
		); 

/******************* CELL 6028 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6028 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5932]),
			.N(gen[5933]),
			.NE(gen[5934]),

			.O(gen[6027]),
			.E(gen[6029]),

			.SO(gen[6122]),
			.S(gen[6123]),
			.SE(gen[6124]),

			.SELF(gen[6028]),
			.cell_state(gen[6028])
		); 

/******************* CELL 6029 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6029 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5933]),
			.N(gen[5934]),
			.NE(gen[5935]),

			.O(gen[6028]),
			.E(gen[6030]),

			.SO(gen[6123]),
			.S(gen[6124]),
			.SE(gen[6125]),

			.SELF(gen[6029]),
			.cell_state(gen[6029])
		); 

/******************* CELL 6030 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6030 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5934]),
			.N(gen[5935]),
			.NE(gen[5936]),

			.O(gen[6029]),
			.E(gen[6031]),

			.SO(gen[6124]),
			.S(gen[6125]),
			.SE(gen[6126]),

			.SELF(gen[6030]),
			.cell_state(gen[6030])
		); 

/******************* CELL 6031 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6031 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5935]),
			.N(gen[5936]),
			.NE(gen[5937]),

			.O(gen[6030]),
			.E(gen[6032]),

			.SO(gen[6125]),
			.S(gen[6126]),
			.SE(gen[6127]),

			.SELF(gen[6031]),
			.cell_state(gen[6031])
		); 

/******************* CELL 6032 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6032 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5936]),
			.N(gen[5937]),
			.NE(gen[5938]),

			.O(gen[6031]),
			.E(gen[6033]),

			.SO(gen[6126]),
			.S(gen[6127]),
			.SE(gen[6128]),

			.SELF(gen[6032]),
			.cell_state(gen[6032])
		); 

/******************* CELL 6033 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6033 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5937]),
			.N(gen[5938]),
			.NE(gen[5939]),

			.O(gen[6032]),
			.E(gen[6034]),

			.SO(gen[6127]),
			.S(gen[6128]),
			.SE(gen[6129]),

			.SELF(gen[6033]),
			.cell_state(gen[6033])
		); 

/******************* CELL 6034 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6034 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5938]),
			.N(gen[5939]),
			.NE(gen[5940]),

			.O(gen[6033]),
			.E(gen[6035]),

			.SO(gen[6128]),
			.S(gen[6129]),
			.SE(gen[6130]),

			.SELF(gen[6034]),
			.cell_state(gen[6034])
		); 

/******************* CELL 6035 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6035 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5939]),
			.N(gen[5940]),
			.NE(gen[5941]),

			.O(gen[6034]),
			.E(gen[6036]),

			.SO(gen[6129]),
			.S(gen[6130]),
			.SE(gen[6131]),

			.SELF(gen[6035]),
			.cell_state(gen[6035])
		); 

/******************* CELL 6036 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6036 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5940]),
			.N(gen[5941]),
			.NE(gen[5942]),

			.O(gen[6035]),
			.E(gen[6037]),

			.SO(gen[6130]),
			.S(gen[6131]),
			.SE(gen[6132]),

			.SELF(gen[6036]),
			.cell_state(gen[6036])
		); 

/******************* CELL 6037 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6037 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5941]),
			.N(gen[5942]),
			.NE(gen[5943]),

			.O(gen[6036]),
			.E(gen[6038]),

			.SO(gen[6131]),
			.S(gen[6132]),
			.SE(gen[6133]),

			.SELF(gen[6037]),
			.cell_state(gen[6037])
		); 

/******************* CELL 6038 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6038 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5942]),
			.N(gen[5943]),
			.NE(gen[5944]),

			.O(gen[6037]),
			.E(gen[6039]),

			.SO(gen[6132]),
			.S(gen[6133]),
			.SE(gen[6134]),

			.SELF(gen[6038]),
			.cell_state(gen[6038])
		); 

/******************* CELL 6039 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6039 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5943]),
			.N(gen[5944]),
			.NE(gen[5945]),

			.O(gen[6038]),
			.E(gen[6040]),

			.SO(gen[6133]),
			.S(gen[6134]),
			.SE(gen[6135]),

			.SELF(gen[6039]),
			.cell_state(gen[6039])
		); 

/******************* CELL 6040 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6040 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5944]),
			.N(gen[5945]),
			.NE(gen[5946]),

			.O(gen[6039]),
			.E(gen[6041]),

			.SO(gen[6134]),
			.S(gen[6135]),
			.SE(gen[6136]),

			.SELF(gen[6040]),
			.cell_state(gen[6040])
		); 

/******************* CELL 6041 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6041 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5945]),
			.N(gen[5946]),
			.NE(gen[5947]),

			.O(gen[6040]),
			.E(gen[6042]),

			.SO(gen[6135]),
			.S(gen[6136]),
			.SE(gen[6137]),

			.SELF(gen[6041]),
			.cell_state(gen[6041])
		); 

/******************* CELL 6042 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6042 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5946]),
			.N(gen[5947]),
			.NE(gen[5948]),

			.O(gen[6041]),
			.E(gen[6043]),

			.SO(gen[6136]),
			.S(gen[6137]),
			.SE(gen[6138]),

			.SELF(gen[6042]),
			.cell_state(gen[6042])
		); 

/******************* CELL 6043 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6043 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5947]),
			.N(gen[5948]),
			.NE(gen[5949]),

			.O(gen[6042]),
			.E(gen[6044]),

			.SO(gen[6137]),
			.S(gen[6138]),
			.SE(gen[6139]),

			.SELF(gen[6043]),
			.cell_state(gen[6043])
		); 

/******************* CELL 6044 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6044 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5948]),
			.N(gen[5949]),
			.NE(gen[5950]),

			.O(gen[6043]),
			.E(gen[6045]),

			.SO(gen[6138]),
			.S(gen[6139]),
			.SE(gen[6140]),

			.SELF(gen[6044]),
			.cell_state(gen[6044])
		); 

/******************* CELL 6045 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6045 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5949]),
			.N(gen[5950]),
			.NE(gen[5951]),

			.O(gen[6044]),
			.E(gen[6046]),

			.SO(gen[6139]),
			.S(gen[6140]),
			.SE(gen[6141]),

			.SELF(gen[6045]),
			.cell_state(gen[6045])
		); 

/******************* CELL 6046 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6046 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5950]),
			.N(gen[5951]),
			.NE(gen[5952]),

			.O(gen[6045]),
			.E(gen[6047]),

			.SO(gen[6140]),
			.S(gen[6141]),
			.SE(gen[6142]),

			.SELF(gen[6046]),
			.cell_state(gen[6046])
		); 

/******************* CELL 6047 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6047 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5951]),
			.N(gen[5952]),
			.NE(gen[5953]),

			.O(gen[6046]),
			.E(gen[6048]),

			.SO(gen[6141]),
			.S(gen[6142]),
			.SE(gen[6143]),

			.SELF(gen[6047]),
			.cell_state(gen[6047])
		); 

/******************* CELL 6048 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6048 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5952]),
			.N(gen[5953]),
			.NE(gen[5954]),

			.O(gen[6047]),
			.E(gen[6049]),

			.SO(gen[6142]),
			.S(gen[6143]),
			.SE(gen[6144]),

			.SELF(gen[6048]),
			.cell_state(gen[6048])
		); 

/******************* CELL 6049 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6049 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5953]),
			.N(gen[5954]),
			.NE(gen[5955]),

			.O(gen[6048]),
			.E(gen[6050]),

			.SO(gen[6143]),
			.S(gen[6144]),
			.SE(gen[6145]),

			.SELF(gen[6049]),
			.cell_state(gen[6049])
		); 

/******************* CELL 6050 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6050 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5954]),
			.N(gen[5955]),
			.NE(gen[5956]),

			.O(gen[6049]),
			.E(gen[6051]),

			.SO(gen[6144]),
			.S(gen[6145]),
			.SE(gen[6146]),

			.SELF(gen[6050]),
			.cell_state(gen[6050])
		); 

/******************* CELL 6051 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6051 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5955]),
			.N(gen[5956]),
			.NE(gen[5957]),

			.O(gen[6050]),
			.E(gen[6052]),

			.SO(gen[6145]),
			.S(gen[6146]),
			.SE(gen[6147]),

			.SELF(gen[6051]),
			.cell_state(gen[6051])
		); 

/******************* CELL 6052 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6052 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5956]),
			.N(gen[5957]),
			.NE(gen[5958]),

			.O(gen[6051]),
			.E(gen[6053]),

			.SO(gen[6146]),
			.S(gen[6147]),
			.SE(gen[6148]),

			.SELF(gen[6052]),
			.cell_state(gen[6052])
		); 

/******************* CELL 6053 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6053 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5957]),
			.N(gen[5958]),
			.NE(gen[5959]),

			.O(gen[6052]),
			.E(gen[6054]),

			.SO(gen[6147]),
			.S(gen[6148]),
			.SE(gen[6149]),

			.SELF(gen[6053]),
			.cell_state(gen[6053])
		); 

/******************* CELL 6054 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6054 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5958]),
			.N(gen[5959]),
			.NE(gen[5960]),

			.O(gen[6053]),
			.E(gen[6055]),

			.SO(gen[6148]),
			.S(gen[6149]),
			.SE(gen[6150]),

			.SELF(gen[6054]),
			.cell_state(gen[6054])
		); 

/******************* CELL 6055 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6055 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5959]),
			.N(gen[5960]),
			.NE(gen[5961]),

			.O(gen[6054]),
			.E(gen[6056]),

			.SO(gen[6149]),
			.S(gen[6150]),
			.SE(gen[6151]),

			.SELF(gen[6055]),
			.cell_state(gen[6055])
		); 

/******************* CELL 6056 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6056 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5960]),
			.N(gen[5961]),
			.NE(gen[5962]),

			.O(gen[6055]),
			.E(gen[6057]),

			.SO(gen[6150]),
			.S(gen[6151]),
			.SE(gen[6152]),

			.SELF(gen[6056]),
			.cell_state(gen[6056])
		); 

/******************* CELL 6057 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6057 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5961]),
			.N(gen[5962]),
			.NE(gen[5963]),

			.O(gen[6056]),
			.E(gen[6058]),

			.SO(gen[6151]),
			.S(gen[6152]),
			.SE(gen[6153]),

			.SELF(gen[6057]),
			.cell_state(gen[6057])
		); 

/******************* CELL 6058 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6058 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5962]),
			.N(gen[5963]),
			.NE(gen[5964]),

			.O(gen[6057]),
			.E(gen[6059]),

			.SO(gen[6152]),
			.S(gen[6153]),
			.SE(gen[6154]),

			.SELF(gen[6058]),
			.cell_state(gen[6058])
		); 

/******************* CELL 6059 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6059 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5963]),
			.N(gen[5964]),
			.NE(gen[5965]),

			.O(gen[6058]),
			.E(gen[6060]),

			.SO(gen[6153]),
			.S(gen[6154]),
			.SE(gen[6155]),

			.SELF(gen[6059]),
			.cell_state(gen[6059])
		); 

/******************* CELL 6060 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6060 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5964]),
			.N(gen[5965]),
			.NE(gen[5966]),

			.O(gen[6059]),
			.E(gen[6061]),

			.SO(gen[6154]),
			.S(gen[6155]),
			.SE(gen[6156]),

			.SELF(gen[6060]),
			.cell_state(gen[6060])
		); 

/******************* CELL 6061 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6061 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5965]),
			.N(gen[5966]),
			.NE(gen[5967]),

			.O(gen[6060]),
			.E(gen[6062]),

			.SO(gen[6155]),
			.S(gen[6156]),
			.SE(gen[6157]),

			.SELF(gen[6061]),
			.cell_state(gen[6061])
		); 

/******************* CELL 6062 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6062 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5966]),
			.N(gen[5967]),
			.NE(gen[5968]),

			.O(gen[6061]),
			.E(gen[6063]),

			.SO(gen[6156]),
			.S(gen[6157]),
			.SE(gen[6158]),

			.SELF(gen[6062]),
			.cell_state(gen[6062])
		); 

/******************* CELL 6063 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6063 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5967]),
			.N(gen[5968]),
			.NE(gen[5969]),

			.O(gen[6062]),
			.E(gen[6064]),

			.SO(gen[6157]),
			.S(gen[6158]),
			.SE(gen[6159]),

			.SELF(gen[6063]),
			.cell_state(gen[6063])
		); 

/******************* CELL 6064 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6064 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5968]),
			.N(gen[5969]),
			.NE(gen[5970]),

			.O(gen[6063]),
			.E(gen[6065]),

			.SO(gen[6158]),
			.S(gen[6159]),
			.SE(gen[6160]),

			.SELF(gen[6064]),
			.cell_state(gen[6064])
		); 

/******************* CELL 6065 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6065 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5969]),
			.N(gen[5970]),
			.NE(gen[5971]),

			.O(gen[6064]),
			.E(gen[6066]),

			.SO(gen[6159]),
			.S(gen[6160]),
			.SE(gen[6161]),

			.SELF(gen[6065]),
			.cell_state(gen[6065])
		); 

/******************* CELL 6066 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6066 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5970]),
			.N(gen[5971]),
			.NE(gen[5972]),

			.O(gen[6065]),
			.E(gen[6067]),

			.SO(gen[6160]),
			.S(gen[6161]),
			.SE(gen[6162]),

			.SELF(gen[6066]),
			.cell_state(gen[6066])
		); 

/******************* CELL 6067 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6067 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5971]),
			.N(gen[5972]),
			.NE(gen[5973]),

			.O(gen[6066]),
			.E(gen[6068]),

			.SO(gen[6161]),
			.S(gen[6162]),
			.SE(gen[6163]),

			.SELF(gen[6067]),
			.cell_state(gen[6067])
		); 

/******************* CELL 6068 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6068 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5972]),
			.N(gen[5973]),
			.NE(gen[5974]),

			.O(gen[6067]),
			.E(gen[6069]),

			.SO(gen[6162]),
			.S(gen[6163]),
			.SE(gen[6164]),

			.SELF(gen[6068]),
			.cell_state(gen[6068])
		); 

/******************* CELL 6069 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6069 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5973]),
			.N(gen[5974]),
			.NE(gen[5975]),

			.O(gen[6068]),
			.E(gen[6070]),

			.SO(gen[6163]),
			.S(gen[6164]),
			.SE(gen[6165]),

			.SELF(gen[6069]),
			.cell_state(gen[6069])
		); 

/******************* CELL 6070 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6070 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5974]),
			.N(gen[5975]),
			.NE(gen[5976]),

			.O(gen[6069]),
			.E(gen[6071]),

			.SO(gen[6164]),
			.S(gen[6165]),
			.SE(gen[6166]),

			.SELF(gen[6070]),
			.cell_state(gen[6070])
		); 

/******************* CELL 6071 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6071 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5975]),
			.N(gen[5976]),
			.NE(gen[5977]),

			.O(gen[6070]),
			.E(gen[6072]),

			.SO(gen[6165]),
			.S(gen[6166]),
			.SE(gen[6167]),

			.SELF(gen[6071]),
			.cell_state(gen[6071])
		); 

/******************* CELL 6072 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6072 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5976]),
			.N(gen[5977]),
			.NE(gen[5978]),

			.O(gen[6071]),
			.E(gen[6073]),

			.SO(gen[6166]),
			.S(gen[6167]),
			.SE(gen[6168]),

			.SELF(gen[6072]),
			.cell_state(gen[6072])
		); 

/******************* CELL 6073 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6073 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5977]),
			.N(gen[5978]),
			.NE(gen[5979]),

			.O(gen[6072]),
			.E(gen[6074]),

			.SO(gen[6167]),
			.S(gen[6168]),
			.SE(gen[6169]),

			.SELF(gen[6073]),
			.cell_state(gen[6073])
		); 

/******************* CELL 6074 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6074 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5978]),
			.N(gen[5979]),
			.NE(gen[5980]),

			.O(gen[6073]),
			.E(gen[6075]),

			.SO(gen[6168]),
			.S(gen[6169]),
			.SE(gen[6170]),

			.SELF(gen[6074]),
			.cell_state(gen[6074])
		); 

/******************* CELL 6075 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6075 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5979]),
			.N(gen[5980]),
			.NE(gen[5981]),

			.O(gen[6074]),
			.E(gen[6076]),

			.SO(gen[6169]),
			.S(gen[6170]),
			.SE(gen[6171]),

			.SELF(gen[6075]),
			.cell_state(gen[6075])
		); 

/******************* CELL 6076 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6076 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5980]),
			.N(gen[5981]),
			.NE(gen[5982]),

			.O(gen[6075]),
			.E(gen[6077]),

			.SO(gen[6170]),
			.S(gen[6171]),
			.SE(gen[6172]),

			.SELF(gen[6076]),
			.cell_state(gen[6076])
		); 

/******************* CELL 6077 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6077 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5981]),
			.N(gen[5982]),
			.NE(gen[5983]),

			.O(gen[6076]),
			.E(gen[6078]),

			.SO(gen[6171]),
			.S(gen[6172]),
			.SE(gen[6173]),

			.SELF(gen[6077]),
			.cell_state(gen[6077])
		); 

/******************* CELL 6078 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6078 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5982]),
			.N(gen[5983]),
			.NE(gen[5984]),

			.O(gen[6077]),
			.E(gen[6079]),

			.SO(gen[6172]),
			.S(gen[6173]),
			.SE(gen[6174]),

			.SELF(gen[6078]),
			.cell_state(gen[6078])
		); 

/******************* CELL 6079 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6079 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5983]),
			.N(gen[5984]),
			.NE(gen[5983]),

			.O(gen[6078]),
			.E(gen[6078]),

			.SO(gen[6173]),
			.S(gen[6174]),
			.SE(gen[6173]),

			.SELF(gen[6079]),
			.cell_state(gen[6079])
		); 

/******************* CELL 6080 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6080 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5986]),
			.N(gen[5985]),
			.NE(gen[5986]),

			.O(gen[6081]),
			.E(gen[6081]),

			.SO(gen[6176]),
			.S(gen[6175]),
			.SE(gen[6176]),

			.SELF(gen[6080]),
			.cell_state(gen[6080])
		); 

/******************* CELL 6081 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6081 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5985]),
			.N(gen[5986]),
			.NE(gen[5987]),

			.O(gen[6080]),
			.E(gen[6082]),

			.SO(gen[6175]),
			.S(gen[6176]),
			.SE(gen[6177]),

			.SELF(gen[6081]),
			.cell_state(gen[6081])
		); 

/******************* CELL 6082 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6082 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5986]),
			.N(gen[5987]),
			.NE(gen[5988]),

			.O(gen[6081]),
			.E(gen[6083]),

			.SO(gen[6176]),
			.S(gen[6177]),
			.SE(gen[6178]),

			.SELF(gen[6082]),
			.cell_state(gen[6082])
		); 

/******************* CELL 6083 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6083 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5987]),
			.N(gen[5988]),
			.NE(gen[5989]),

			.O(gen[6082]),
			.E(gen[6084]),

			.SO(gen[6177]),
			.S(gen[6178]),
			.SE(gen[6179]),

			.SELF(gen[6083]),
			.cell_state(gen[6083])
		); 

/******************* CELL 6084 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6084 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5988]),
			.N(gen[5989]),
			.NE(gen[5990]),

			.O(gen[6083]),
			.E(gen[6085]),

			.SO(gen[6178]),
			.S(gen[6179]),
			.SE(gen[6180]),

			.SELF(gen[6084]),
			.cell_state(gen[6084])
		); 

/******************* CELL 6085 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6085 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5989]),
			.N(gen[5990]),
			.NE(gen[5991]),

			.O(gen[6084]),
			.E(gen[6086]),

			.SO(gen[6179]),
			.S(gen[6180]),
			.SE(gen[6181]),

			.SELF(gen[6085]),
			.cell_state(gen[6085])
		); 

/******************* CELL 6086 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6086 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5990]),
			.N(gen[5991]),
			.NE(gen[5992]),

			.O(gen[6085]),
			.E(gen[6087]),

			.SO(gen[6180]),
			.S(gen[6181]),
			.SE(gen[6182]),

			.SELF(gen[6086]),
			.cell_state(gen[6086])
		); 

/******************* CELL 6087 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6087 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5991]),
			.N(gen[5992]),
			.NE(gen[5993]),

			.O(gen[6086]),
			.E(gen[6088]),

			.SO(gen[6181]),
			.S(gen[6182]),
			.SE(gen[6183]),

			.SELF(gen[6087]),
			.cell_state(gen[6087])
		); 

/******************* CELL 6088 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6088 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5992]),
			.N(gen[5993]),
			.NE(gen[5994]),

			.O(gen[6087]),
			.E(gen[6089]),

			.SO(gen[6182]),
			.S(gen[6183]),
			.SE(gen[6184]),

			.SELF(gen[6088]),
			.cell_state(gen[6088])
		); 

/******************* CELL 6089 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6089 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5993]),
			.N(gen[5994]),
			.NE(gen[5995]),

			.O(gen[6088]),
			.E(gen[6090]),

			.SO(gen[6183]),
			.S(gen[6184]),
			.SE(gen[6185]),

			.SELF(gen[6089]),
			.cell_state(gen[6089])
		); 

/******************* CELL 6090 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6090 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5994]),
			.N(gen[5995]),
			.NE(gen[5996]),

			.O(gen[6089]),
			.E(gen[6091]),

			.SO(gen[6184]),
			.S(gen[6185]),
			.SE(gen[6186]),

			.SELF(gen[6090]),
			.cell_state(gen[6090])
		); 

/******************* CELL 6091 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6091 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5995]),
			.N(gen[5996]),
			.NE(gen[5997]),

			.O(gen[6090]),
			.E(gen[6092]),

			.SO(gen[6185]),
			.S(gen[6186]),
			.SE(gen[6187]),

			.SELF(gen[6091]),
			.cell_state(gen[6091])
		); 

/******************* CELL 6092 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6092 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5996]),
			.N(gen[5997]),
			.NE(gen[5998]),

			.O(gen[6091]),
			.E(gen[6093]),

			.SO(gen[6186]),
			.S(gen[6187]),
			.SE(gen[6188]),

			.SELF(gen[6092]),
			.cell_state(gen[6092])
		); 

/******************* CELL 6093 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6093 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5997]),
			.N(gen[5998]),
			.NE(gen[5999]),

			.O(gen[6092]),
			.E(gen[6094]),

			.SO(gen[6187]),
			.S(gen[6188]),
			.SE(gen[6189]),

			.SELF(gen[6093]),
			.cell_state(gen[6093])
		); 

/******************* CELL 6094 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6094 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5998]),
			.N(gen[5999]),
			.NE(gen[6000]),

			.O(gen[6093]),
			.E(gen[6095]),

			.SO(gen[6188]),
			.S(gen[6189]),
			.SE(gen[6190]),

			.SELF(gen[6094]),
			.cell_state(gen[6094])
		); 

/******************* CELL 6095 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6095 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5999]),
			.N(gen[6000]),
			.NE(gen[6001]),

			.O(gen[6094]),
			.E(gen[6096]),

			.SO(gen[6189]),
			.S(gen[6190]),
			.SE(gen[6191]),

			.SELF(gen[6095]),
			.cell_state(gen[6095])
		); 

/******************* CELL 6096 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6096 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6000]),
			.N(gen[6001]),
			.NE(gen[6002]),

			.O(gen[6095]),
			.E(gen[6097]),

			.SO(gen[6190]),
			.S(gen[6191]),
			.SE(gen[6192]),

			.SELF(gen[6096]),
			.cell_state(gen[6096])
		); 

/******************* CELL 6097 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6097 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6001]),
			.N(gen[6002]),
			.NE(gen[6003]),

			.O(gen[6096]),
			.E(gen[6098]),

			.SO(gen[6191]),
			.S(gen[6192]),
			.SE(gen[6193]),

			.SELF(gen[6097]),
			.cell_state(gen[6097])
		); 

/******************* CELL 6098 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6098 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6002]),
			.N(gen[6003]),
			.NE(gen[6004]),

			.O(gen[6097]),
			.E(gen[6099]),

			.SO(gen[6192]),
			.S(gen[6193]),
			.SE(gen[6194]),

			.SELF(gen[6098]),
			.cell_state(gen[6098])
		); 

/******************* CELL 6099 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6099 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6003]),
			.N(gen[6004]),
			.NE(gen[6005]),

			.O(gen[6098]),
			.E(gen[6100]),

			.SO(gen[6193]),
			.S(gen[6194]),
			.SE(gen[6195]),

			.SELF(gen[6099]),
			.cell_state(gen[6099])
		); 

/******************* CELL 6100 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6100 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6004]),
			.N(gen[6005]),
			.NE(gen[6006]),

			.O(gen[6099]),
			.E(gen[6101]),

			.SO(gen[6194]),
			.S(gen[6195]),
			.SE(gen[6196]),

			.SELF(gen[6100]),
			.cell_state(gen[6100])
		); 

/******************* CELL 6101 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6101 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6005]),
			.N(gen[6006]),
			.NE(gen[6007]),

			.O(gen[6100]),
			.E(gen[6102]),

			.SO(gen[6195]),
			.S(gen[6196]),
			.SE(gen[6197]),

			.SELF(gen[6101]),
			.cell_state(gen[6101])
		); 

/******************* CELL 6102 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6102 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6006]),
			.N(gen[6007]),
			.NE(gen[6008]),

			.O(gen[6101]),
			.E(gen[6103]),

			.SO(gen[6196]),
			.S(gen[6197]),
			.SE(gen[6198]),

			.SELF(gen[6102]),
			.cell_state(gen[6102])
		); 

/******************* CELL 6103 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6103 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6007]),
			.N(gen[6008]),
			.NE(gen[6009]),

			.O(gen[6102]),
			.E(gen[6104]),

			.SO(gen[6197]),
			.S(gen[6198]),
			.SE(gen[6199]),

			.SELF(gen[6103]),
			.cell_state(gen[6103])
		); 

/******************* CELL 6104 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6104 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6008]),
			.N(gen[6009]),
			.NE(gen[6010]),

			.O(gen[6103]),
			.E(gen[6105]),

			.SO(gen[6198]),
			.S(gen[6199]),
			.SE(gen[6200]),

			.SELF(gen[6104]),
			.cell_state(gen[6104])
		); 

/******************* CELL 6105 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6105 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6009]),
			.N(gen[6010]),
			.NE(gen[6011]),

			.O(gen[6104]),
			.E(gen[6106]),

			.SO(gen[6199]),
			.S(gen[6200]),
			.SE(gen[6201]),

			.SELF(gen[6105]),
			.cell_state(gen[6105])
		); 

/******************* CELL 6106 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6106 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6010]),
			.N(gen[6011]),
			.NE(gen[6012]),

			.O(gen[6105]),
			.E(gen[6107]),

			.SO(gen[6200]),
			.S(gen[6201]),
			.SE(gen[6202]),

			.SELF(gen[6106]),
			.cell_state(gen[6106])
		); 

/******************* CELL 6107 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6107 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6011]),
			.N(gen[6012]),
			.NE(gen[6013]),

			.O(gen[6106]),
			.E(gen[6108]),

			.SO(gen[6201]),
			.S(gen[6202]),
			.SE(gen[6203]),

			.SELF(gen[6107]),
			.cell_state(gen[6107])
		); 

/******************* CELL 6108 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6108 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6012]),
			.N(gen[6013]),
			.NE(gen[6014]),

			.O(gen[6107]),
			.E(gen[6109]),

			.SO(gen[6202]),
			.S(gen[6203]),
			.SE(gen[6204]),

			.SELF(gen[6108]),
			.cell_state(gen[6108])
		); 

/******************* CELL 6109 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6109 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6013]),
			.N(gen[6014]),
			.NE(gen[6015]),

			.O(gen[6108]),
			.E(gen[6110]),

			.SO(gen[6203]),
			.S(gen[6204]),
			.SE(gen[6205]),

			.SELF(gen[6109]),
			.cell_state(gen[6109])
		); 

/******************* CELL 6110 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6110 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6014]),
			.N(gen[6015]),
			.NE(gen[6016]),

			.O(gen[6109]),
			.E(gen[6111]),

			.SO(gen[6204]),
			.S(gen[6205]),
			.SE(gen[6206]),

			.SELF(gen[6110]),
			.cell_state(gen[6110])
		); 

/******************* CELL 6111 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6111 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6015]),
			.N(gen[6016]),
			.NE(gen[6017]),

			.O(gen[6110]),
			.E(gen[6112]),

			.SO(gen[6205]),
			.S(gen[6206]),
			.SE(gen[6207]),

			.SELF(gen[6111]),
			.cell_state(gen[6111])
		); 

/******************* CELL 6112 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6112 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6016]),
			.N(gen[6017]),
			.NE(gen[6018]),

			.O(gen[6111]),
			.E(gen[6113]),

			.SO(gen[6206]),
			.S(gen[6207]),
			.SE(gen[6208]),

			.SELF(gen[6112]),
			.cell_state(gen[6112])
		); 

/******************* CELL 6113 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6113 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6017]),
			.N(gen[6018]),
			.NE(gen[6019]),

			.O(gen[6112]),
			.E(gen[6114]),

			.SO(gen[6207]),
			.S(gen[6208]),
			.SE(gen[6209]),

			.SELF(gen[6113]),
			.cell_state(gen[6113])
		); 

/******************* CELL 6114 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6114 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6018]),
			.N(gen[6019]),
			.NE(gen[6020]),

			.O(gen[6113]),
			.E(gen[6115]),

			.SO(gen[6208]),
			.S(gen[6209]),
			.SE(gen[6210]),

			.SELF(gen[6114]),
			.cell_state(gen[6114])
		); 

/******************* CELL 6115 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6115 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6019]),
			.N(gen[6020]),
			.NE(gen[6021]),

			.O(gen[6114]),
			.E(gen[6116]),

			.SO(gen[6209]),
			.S(gen[6210]),
			.SE(gen[6211]),

			.SELF(gen[6115]),
			.cell_state(gen[6115])
		); 

/******************* CELL 6116 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6116 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6020]),
			.N(gen[6021]),
			.NE(gen[6022]),

			.O(gen[6115]),
			.E(gen[6117]),

			.SO(gen[6210]),
			.S(gen[6211]),
			.SE(gen[6212]),

			.SELF(gen[6116]),
			.cell_state(gen[6116])
		); 

/******************* CELL 6117 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6117 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6021]),
			.N(gen[6022]),
			.NE(gen[6023]),

			.O(gen[6116]),
			.E(gen[6118]),

			.SO(gen[6211]),
			.S(gen[6212]),
			.SE(gen[6213]),

			.SELF(gen[6117]),
			.cell_state(gen[6117])
		); 

/******************* CELL 6118 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6118 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6022]),
			.N(gen[6023]),
			.NE(gen[6024]),

			.O(gen[6117]),
			.E(gen[6119]),

			.SO(gen[6212]),
			.S(gen[6213]),
			.SE(gen[6214]),

			.SELF(gen[6118]),
			.cell_state(gen[6118])
		); 

/******************* CELL 6119 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6119 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6023]),
			.N(gen[6024]),
			.NE(gen[6025]),

			.O(gen[6118]),
			.E(gen[6120]),

			.SO(gen[6213]),
			.S(gen[6214]),
			.SE(gen[6215]),

			.SELF(gen[6119]),
			.cell_state(gen[6119])
		); 

/******************* CELL 6120 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6120 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6024]),
			.N(gen[6025]),
			.NE(gen[6026]),

			.O(gen[6119]),
			.E(gen[6121]),

			.SO(gen[6214]),
			.S(gen[6215]),
			.SE(gen[6216]),

			.SELF(gen[6120]),
			.cell_state(gen[6120])
		); 

/******************* CELL 6121 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6121 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6025]),
			.N(gen[6026]),
			.NE(gen[6027]),

			.O(gen[6120]),
			.E(gen[6122]),

			.SO(gen[6215]),
			.S(gen[6216]),
			.SE(gen[6217]),

			.SELF(gen[6121]),
			.cell_state(gen[6121])
		); 

/******************* CELL 6122 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6122 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6026]),
			.N(gen[6027]),
			.NE(gen[6028]),

			.O(gen[6121]),
			.E(gen[6123]),

			.SO(gen[6216]),
			.S(gen[6217]),
			.SE(gen[6218]),

			.SELF(gen[6122]),
			.cell_state(gen[6122])
		); 

/******************* CELL 6123 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6123 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6027]),
			.N(gen[6028]),
			.NE(gen[6029]),

			.O(gen[6122]),
			.E(gen[6124]),

			.SO(gen[6217]),
			.S(gen[6218]),
			.SE(gen[6219]),

			.SELF(gen[6123]),
			.cell_state(gen[6123])
		); 

/******************* CELL 6124 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6124 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6028]),
			.N(gen[6029]),
			.NE(gen[6030]),

			.O(gen[6123]),
			.E(gen[6125]),

			.SO(gen[6218]),
			.S(gen[6219]),
			.SE(gen[6220]),

			.SELF(gen[6124]),
			.cell_state(gen[6124])
		); 

/******************* CELL 6125 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6125 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6029]),
			.N(gen[6030]),
			.NE(gen[6031]),

			.O(gen[6124]),
			.E(gen[6126]),

			.SO(gen[6219]),
			.S(gen[6220]),
			.SE(gen[6221]),

			.SELF(gen[6125]),
			.cell_state(gen[6125])
		); 

/******************* CELL 6126 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6126 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6030]),
			.N(gen[6031]),
			.NE(gen[6032]),

			.O(gen[6125]),
			.E(gen[6127]),

			.SO(gen[6220]),
			.S(gen[6221]),
			.SE(gen[6222]),

			.SELF(gen[6126]),
			.cell_state(gen[6126])
		); 

/******************* CELL 6127 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6127 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6031]),
			.N(gen[6032]),
			.NE(gen[6033]),

			.O(gen[6126]),
			.E(gen[6128]),

			.SO(gen[6221]),
			.S(gen[6222]),
			.SE(gen[6223]),

			.SELF(gen[6127]),
			.cell_state(gen[6127])
		); 

/******************* CELL 6128 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6128 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6032]),
			.N(gen[6033]),
			.NE(gen[6034]),

			.O(gen[6127]),
			.E(gen[6129]),

			.SO(gen[6222]),
			.S(gen[6223]),
			.SE(gen[6224]),

			.SELF(gen[6128]),
			.cell_state(gen[6128])
		); 

/******************* CELL 6129 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6129 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6033]),
			.N(gen[6034]),
			.NE(gen[6035]),

			.O(gen[6128]),
			.E(gen[6130]),

			.SO(gen[6223]),
			.S(gen[6224]),
			.SE(gen[6225]),

			.SELF(gen[6129]),
			.cell_state(gen[6129])
		); 

/******************* CELL 6130 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6130 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6034]),
			.N(gen[6035]),
			.NE(gen[6036]),

			.O(gen[6129]),
			.E(gen[6131]),

			.SO(gen[6224]),
			.S(gen[6225]),
			.SE(gen[6226]),

			.SELF(gen[6130]),
			.cell_state(gen[6130])
		); 

/******************* CELL 6131 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6131 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6035]),
			.N(gen[6036]),
			.NE(gen[6037]),

			.O(gen[6130]),
			.E(gen[6132]),

			.SO(gen[6225]),
			.S(gen[6226]),
			.SE(gen[6227]),

			.SELF(gen[6131]),
			.cell_state(gen[6131])
		); 

/******************* CELL 6132 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6132 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6036]),
			.N(gen[6037]),
			.NE(gen[6038]),

			.O(gen[6131]),
			.E(gen[6133]),

			.SO(gen[6226]),
			.S(gen[6227]),
			.SE(gen[6228]),

			.SELF(gen[6132]),
			.cell_state(gen[6132])
		); 

/******************* CELL 6133 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6133 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6037]),
			.N(gen[6038]),
			.NE(gen[6039]),

			.O(gen[6132]),
			.E(gen[6134]),

			.SO(gen[6227]),
			.S(gen[6228]),
			.SE(gen[6229]),

			.SELF(gen[6133]),
			.cell_state(gen[6133])
		); 

/******************* CELL 6134 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6134 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6038]),
			.N(gen[6039]),
			.NE(gen[6040]),

			.O(gen[6133]),
			.E(gen[6135]),

			.SO(gen[6228]),
			.S(gen[6229]),
			.SE(gen[6230]),

			.SELF(gen[6134]),
			.cell_state(gen[6134])
		); 

/******************* CELL 6135 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6135 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6039]),
			.N(gen[6040]),
			.NE(gen[6041]),

			.O(gen[6134]),
			.E(gen[6136]),

			.SO(gen[6229]),
			.S(gen[6230]),
			.SE(gen[6231]),

			.SELF(gen[6135]),
			.cell_state(gen[6135])
		); 

/******************* CELL 6136 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6136 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6040]),
			.N(gen[6041]),
			.NE(gen[6042]),

			.O(gen[6135]),
			.E(gen[6137]),

			.SO(gen[6230]),
			.S(gen[6231]),
			.SE(gen[6232]),

			.SELF(gen[6136]),
			.cell_state(gen[6136])
		); 

/******************* CELL 6137 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6137 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6041]),
			.N(gen[6042]),
			.NE(gen[6043]),

			.O(gen[6136]),
			.E(gen[6138]),

			.SO(gen[6231]),
			.S(gen[6232]),
			.SE(gen[6233]),

			.SELF(gen[6137]),
			.cell_state(gen[6137])
		); 

/******************* CELL 6138 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6138 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6042]),
			.N(gen[6043]),
			.NE(gen[6044]),

			.O(gen[6137]),
			.E(gen[6139]),

			.SO(gen[6232]),
			.S(gen[6233]),
			.SE(gen[6234]),

			.SELF(gen[6138]),
			.cell_state(gen[6138])
		); 

/******************* CELL 6139 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6139 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6043]),
			.N(gen[6044]),
			.NE(gen[6045]),

			.O(gen[6138]),
			.E(gen[6140]),

			.SO(gen[6233]),
			.S(gen[6234]),
			.SE(gen[6235]),

			.SELF(gen[6139]),
			.cell_state(gen[6139])
		); 

/******************* CELL 6140 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6140 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6044]),
			.N(gen[6045]),
			.NE(gen[6046]),

			.O(gen[6139]),
			.E(gen[6141]),

			.SO(gen[6234]),
			.S(gen[6235]),
			.SE(gen[6236]),

			.SELF(gen[6140]),
			.cell_state(gen[6140])
		); 

/******************* CELL 6141 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6141 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6045]),
			.N(gen[6046]),
			.NE(gen[6047]),

			.O(gen[6140]),
			.E(gen[6142]),

			.SO(gen[6235]),
			.S(gen[6236]),
			.SE(gen[6237]),

			.SELF(gen[6141]),
			.cell_state(gen[6141])
		); 

/******************* CELL 6142 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6142 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6046]),
			.N(gen[6047]),
			.NE(gen[6048]),

			.O(gen[6141]),
			.E(gen[6143]),

			.SO(gen[6236]),
			.S(gen[6237]),
			.SE(gen[6238]),

			.SELF(gen[6142]),
			.cell_state(gen[6142])
		); 

/******************* CELL 6143 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6143 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6047]),
			.N(gen[6048]),
			.NE(gen[6049]),

			.O(gen[6142]),
			.E(gen[6144]),

			.SO(gen[6237]),
			.S(gen[6238]),
			.SE(gen[6239]),

			.SELF(gen[6143]),
			.cell_state(gen[6143])
		); 

/******************* CELL 6144 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6144 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6048]),
			.N(gen[6049]),
			.NE(gen[6050]),

			.O(gen[6143]),
			.E(gen[6145]),

			.SO(gen[6238]),
			.S(gen[6239]),
			.SE(gen[6240]),

			.SELF(gen[6144]),
			.cell_state(gen[6144])
		); 

/******************* CELL 6145 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6145 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6049]),
			.N(gen[6050]),
			.NE(gen[6051]),

			.O(gen[6144]),
			.E(gen[6146]),

			.SO(gen[6239]),
			.S(gen[6240]),
			.SE(gen[6241]),

			.SELF(gen[6145]),
			.cell_state(gen[6145])
		); 

/******************* CELL 6146 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6146 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6050]),
			.N(gen[6051]),
			.NE(gen[6052]),

			.O(gen[6145]),
			.E(gen[6147]),

			.SO(gen[6240]),
			.S(gen[6241]),
			.SE(gen[6242]),

			.SELF(gen[6146]),
			.cell_state(gen[6146])
		); 

/******************* CELL 6147 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6147 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6051]),
			.N(gen[6052]),
			.NE(gen[6053]),

			.O(gen[6146]),
			.E(gen[6148]),

			.SO(gen[6241]),
			.S(gen[6242]),
			.SE(gen[6243]),

			.SELF(gen[6147]),
			.cell_state(gen[6147])
		); 

/******************* CELL 6148 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6148 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6052]),
			.N(gen[6053]),
			.NE(gen[6054]),

			.O(gen[6147]),
			.E(gen[6149]),

			.SO(gen[6242]),
			.S(gen[6243]),
			.SE(gen[6244]),

			.SELF(gen[6148]),
			.cell_state(gen[6148])
		); 

/******************* CELL 6149 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6149 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6053]),
			.N(gen[6054]),
			.NE(gen[6055]),

			.O(gen[6148]),
			.E(gen[6150]),

			.SO(gen[6243]),
			.S(gen[6244]),
			.SE(gen[6245]),

			.SELF(gen[6149]),
			.cell_state(gen[6149])
		); 

/******************* CELL 6150 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6150 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6054]),
			.N(gen[6055]),
			.NE(gen[6056]),

			.O(gen[6149]),
			.E(gen[6151]),

			.SO(gen[6244]),
			.S(gen[6245]),
			.SE(gen[6246]),

			.SELF(gen[6150]),
			.cell_state(gen[6150])
		); 

/******************* CELL 6151 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6151 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6055]),
			.N(gen[6056]),
			.NE(gen[6057]),

			.O(gen[6150]),
			.E(gen[6152]),

			.SO(gen[6245]),
			.S(gen[6246]),
			.SE(gen[6247]),

			.SELF(gen[6151]),
			.cell_state(gen[6151])
		); 

/******************* CELL 6152 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6152 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6056]),
			.N(gen[6057]),
			.NE(gen[6058]),

			.O(gen[6151]),
			.E(gen[6153]),

			.SO(gen[6246]),
			.S(gen[6247]),
			.SE(gen[6248]),

			.SELF(gen[6152]),
			.cell_state(gen[6152])
		); 

/******************* CELL 6153 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6153 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6057]),
			.N(gen[6058]),
			.NE(gen[6059]),

			.O(gen[6152]),
			.E(gen[6154]),

			.SO(gen[6247]),
			.S(gen[6248]),
			.SE(gen[6249]),

			.SELF(gen[6153]),
			.cell_state(gen[6153])
		); 

/******************* CELL 6154 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6154 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6058]),
			.N(gen[6059]),
			.NE(gen[6060]),

			.O(gen[6153]),
			.E(gen[6155]),

			.SO(gen[6248]),
			.S(gen[6249]),
			.SE(gen[6250]),

			.SELF(gen[6154]),
			.cell_state(gen[6154])
		); 

/******************* CELL 6155 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6155 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6059]),
			.N(gen[6060]),
			.NE(gen[6061]),

			.O(gen[6154]),
			.E(gen[6156]),

			.SO(gen[6249]),
			.S(gen[6250]),
			.SE(gen[6251]),

			.SELF(gen[6155]),
			.cell_state(gen[6155])
		); 

/******************* CELL 6156 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6156 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6060]),
			.N(gen[6061]),
			.NE(gen[6062]),

			.O(gen[6155]),
			.E(gen[6157]),

			.SO(gen[6250]),
			.S(gen[6251]),
			.SE(gen[6252]),

			.SELF(gen[6156]),
			.cell_state(gen[6156])
		); 

/******************* CELL 6157 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6157 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6061]),
			.N(gen[6062]),
			.NE(gen[6063]),

			.O(gen[6156]),
			.E(gen[6158]),

			.SO(gen[6251]),
			.S(gen[6252]),
			.SE(gen[6253]),

			.SELF(gen[6157]),
			.cell_state(gen[6157])
		); 

/******************* CELL 6158 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6158 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6062]),
			.N(gen[6063]),
			.NE(gen[6064]),

			.O(gen[6157]),
			.E(gen[6159]),

			.SO(gen[6252]),
			.S(gen[6253]),
			.SE(gen[6254]),

			.SELF(gen[6158]),
			.cell_state(gen[6158])
		); 

/******************* CELL 6159 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6159 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6063]),
			.N(gen[6064]),
			.NE(gen[6065]),

			.O(gen[6158]),
			.E(gen[6160]),

			.SO(gen[6253]),
			.S(gen[6254]),
			.SE(gen[6255]),

			.SELF(gen[6159]),
			.cell_state(gen[6159])
		); 

/******************* CELL 6160 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6160 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6064]),
			.N(gen[6065]),
			.NE(gen[6066]),

			.O(gen[6159]),
			.E(gen[6161]),

			.SO(gen[6254]),
			.S(gen[6255]),
			.SE(gen[6256]),

			.SELF(gen[6160]),
			.cell_state(gen[6160])
		); 

/******************* CELL 6161 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6161 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6065]),
			.N(gen[6066]),
			.NE(gen[6067]),

			.O(gen[6160]),
			.E(gen[6162]),

			.SO(gen[6255]),
			.S(gen[6256]),
			.SE(gen[6257]),

			.SELF(gen[6161]),
			.cell_state(gen[6161])
		); 

/******************* CELL 6162 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6162 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6066]),
			.N(gen[6067]),
			.NE(gen[6068]),

			.O(gen[6161]),
			.E(gen[6163]),

			.SO(gen[6256]),
			.S(gen[6257]),
			.SE(gen[6258]),

			.SELF(gen[6162]),
			.cell_state(gen[6162])
		); 

/******************* CELL 6163 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6163 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6067]),
			.N(gen[6068]),
			.NE(gen[6069]),

			.O(gen[6162]),
			.E(gen[6164]),

			.SO(gen[6257]),
			.S(gen[6258]),
			.SE(gen[6259]),

			.SELF(gen[6163]),
			.cell_state(gen[6163])
		); 

/******************* CELL 6164 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6164 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6068]),
			.N(gen[6069]),
			.NE(gen[6070]),

			.O(gen[6163]),
			.E(gen[6165]),

			.SO(gen[6258]),
			.S(gen[6259]),
			.SE(gen[6260]),

			.SELF(gen[6164]),
			.cell_state(gen[6164])
		); 

/******************* CELL 6165 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6165 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6069]),
			.N(gen[6070]),
			.NE(gen[6071]),

			.O(gen[6164]),
			.E(gen[6166]),

			.SO(gen[6259]),
			.S(gen[6260]),
			.SE(gen[6261]),

			.SELF(gen[6165]),
			.cell_state(gen[6165])
		); 

/******************* CELL 6166 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6166 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6070]),
			.N(gen[6071]),
			.NE(gen[6072]),

			.O(gen[6165]),
			.E(gen[6167]),

			.SO(gen[6260]),
			.S(gen[6261]),
			.SE(gen[6262]),

			.SELF(gen[6166]),
			.cell_state(gen[6166])
		); 

/******************* CELL 6167 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6167 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6071]),
			.N(gen[6072]),
			.NE(gen[6073]),

			.O(gen[6166]),
			.E(gen[6168]),

			.SO(gen[6261]),
			.S(gen[6262]),
			.SE(gen[6263]),

			.SELF(gen[6167]),
			.cell_state(gen[6167])
		); 

/******************* CELL 6168 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6168 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6072]),
			.N(gen[6073]),
			.NE(gen[6074]),

			.O(gen[6167]),
			.E(gen[6169]),

			.SO(gen[6262]),
			.S(gen[6263]),
			.SE(gen[6264]),

			.SELF(gen[6168]),
			.cell_state(gen[6168])
		); 

/******************* CELL 6169 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6169 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6073]),
			.N(gen[6074]),
			.NE(gen[6075]),

			.O(gen[6168]),
			.E(gen[6170]),

			.SO(gen[6263]),
			.S(gen[6264]),
			.SE(gen[6265]),

			.SELF(gen[6169]),
			.cell_state(gen[6169])
		); 

/******************* CELL 6170 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6170 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6074]),
			.N(gen[6075]),
			.NE(gen[6076]),

			.O(gen[6169]),
			.E(gen[6171]),

			.SO(gen[6264]),
			.S(gen[6265]),
			.SE(gen[6266]),

			.SELF(gen[6170]),
			.cell_state(gen[6170])
		); 

/******************* CELL 6171 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6171 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6075]),
			.N(gen[6076]),
			.NE(gen[6077]),

			.O(gen[6170]),
			.E(gen[6172]),

			.SO(gen[6265]),
			.S(gen[6266]),
			.SE(gen[6267]),

			.SELF(gen[6171]),
			.cell_state(gen[6171])
		); 

/******************* CELL 6172 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6172 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6076]),
			.N(gen[6077]),
			.NE(gen[6078]),

			.O(gen[6171]),
			.E(gen[6173]),

			.SO(gen[6266]),
			.S(gen[6267]),
			.SE(gen[6268]),

			.SELF(gen[6172]),
			.cell_state(gen[6172])
		); 

/******************* CELL 6173 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6173 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6077]),
			.N(gen[6078]),
			.NE(gen[6079]),

			.O(gen[6172]),
			.E(gen[6174]),

			.SO(gen[6267]),
			.S(gen[6268]),
			.SE(gen[6269]),

			.SELF(gen[6173]),
			.cell_state(gen[6173])
		); 

/******************* CELL 6174 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6174 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6078]),
			.N(gen[6079]),
			.NE(gen[6078]),

			.O(gen[6173]),
			.E(gen[6173]),

			.SO(gen[6268]),
			.S(gen[6269]),
			.SE(gen[6268]),

			.SELF(gen[6174]),
			.cell_state(gen[6174])
		); 

/******************* CELL 6175 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6175 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6081]),
			.N(gen[6080]),
			.NE(gen[6081]),

			.O(gen[6176]),
			.E(gen[6176]),

			.SO(gen[6271]),
			.S(gen[6270]),
			.SE(gen[6271]),

			.SELF(gen[6175]),
			.cell_state(gen[6175])
		); 

/******************* CELL 6176 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6176 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6080]),
			.N(gen[6081]),
			.NE(gen[6082]),

			.O(gen[6175]),
			.E(gen[6177]),

			.SO(gen[6270]),
			.S(gen[6271]),
			.SE(gen[6272]),

			.SELF(gen[6176]),
			.cell_state(gen[6176])
		); 

/******************* CELL 6177 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6177 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6081]),
			.N(gen[6082]),
			.NE(gen[6083]),

			.O(gen[6176]),
			.E(gen[6178]),

			.SO(gen[6271]),
			.S(gen[6272]),
			.SE(gen[6273]),

			.SELF(gen[6177]),
			.cell_state(gen[6177])
		); 

/******************* CELL 6178 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6178 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6082]),
			.N(gen[6083]),
			.NE(gen[6084]),

			.O(gen[6177]),
			.E(gen[6179]),

			.SO(gen[6272]),
			.S(gen[6273]),
			.SE(gen[6274]),

			.SELF(gen[6178]),
			.cell_state(gen[6178])
		); 

/******************* CELL 6179 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6179 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6083]),
			.N(gen[6084]),
			.NE(gen[6085]),

			.O(gen[6178]),
			.E(gen[6180]),

			.SO(gen[6273]),
			.S(gen[6274]),
			.SE(gen[6275]),

			.SELF(gen[6179]),
			.cell_state(gen[6179])
		); 

/******************* CELL 6180 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6180 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6084]),
			.N(gen[6085]),
			.NE(gen[6086]),

			.O(gen[6179]),
			.E(gen[6181]),

			.SO(gen[6274]),
			.S(gen[6275]),
			.SE(gen[6276]),

			.SELF(gen[6180]),
			.cell_state(gen[6180])
		); 

/******************* CELL 6181 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6181 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6085]),
			.N(gen[6086]),
			.NE(gen[6087]),

			.O(gen[6180]),
			.E(gen[6182]),

			.SO(gen[6275]),
			.S(gen[6276]),
			.SE(gen[6277]),

			.SELF(gen[6181]),
			.cell_state(gen[6181])
		); 

/******************* CELL 6182 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6182 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6086]),
			.N(gen[6087]),
			.NE(gen[6088]),

			.O(gen[6181]),
			.E(gen[6183]),

			.SO(gen[6276]),
			.S(gen[6277]),
			.SE(gen[6278]),

			.SELF(gen[6182]),
			.cell_state(gen[6182])
		); 

/******************* CELL 6183 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6183 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6087]),
			.N(gen[6088]),
			.NE(gen[6089]),

			.O(gen[6182]),
			.E(gen[6184]),

			.SO(gen[6277]),
			.S(gen[6278]),
			.SE(gen[6279]),

			.SELF(gen[6183]),
			.cell_state(gen[6183])
		); 

/******************* CELL 6184 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6184 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6088]),
			.N(gen[6089]),
			.NE(gen[6090]),

			.O(gen[6183]),
			.E(gen[6185]),

			.SO(gen[6278]),
			.S(gen[6279]),
			.SE(gen[6280]),

			.SELF(gen[6184]),
			.cell_state(gen[6184])
		); 

/******************* CELL 6185 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6185 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6089]),
			.N(gen[6090]),
			.NE(gen[6091]),

			.O(gen[6184]),
			.E(gen[6186]),

			.SO(gen[6279]),
			.S(gen[6280]),
			.SE(gen[6281]),

			.SELF(gen[6185]),
			.cell_state(gen[6185])
		); 

/******************* CELL 6186 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6186 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6090]),
			.N(gen[6091]),
			.NE(gen[6092]),

			.O(gen[6185]),
			.E(gen[6187]),

			.SO(gen[6280]),
			.S(gen[6281]),
			.SE(gen[6282]),

			.SELF(gen[6186]),
			.cell_state(gen[6186])
		); 

/******************* CELL 6187 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6187 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6091]),
			.N(gen[6092]),
			.NE(gen[6093]),

			.O(gen[6186]),
			.E(gen[6188]),

			.SO(gen[6281]),
			.S(gen[6282]),
			.SE(gen[6283]),

			.SELF(gen[6187]),
			.cell_state(gen[6187])
		); 

/******************* CELL 6188 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6188 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6092]),
			.N(gen[6093]),
			.NE(gen[6094]),

			.O(gen[6187]),
			.E(gen[6189]),

			.SO(gen[6282]),
			.S(gen[6283]),
			.SE(gen[6284]),

			.SELF(gen[6188]),
			.cell_state(gen[6188])
		); 

/******************* CELL 6189 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6189 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6093]),
			.N(gen[6094]),
			.NE(gen[6095]),

			.O(gen[6188]),
			.E(gen[6190]),

			.SO(gen[6283]),
			.S(gen[6284]),
			.SE(gen[6285]),

			.SELF(gen[6189]),
			.cell_state(gen[6189])
		); 

/******************* CELL 6190 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6190 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6094]),
			.N(gen[6095]),
			.NE(gen[6096]),

			.O(gen[6189]),
			.E(gen[6191]),

			.SO(gen[6284]),
			.S(gen[6285]),
			.SE(gen[6286]),

			.SELF(gen[6190]),
			.cell_state(gen[6190])
		); 

/******************* CELL 6191 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6191 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6095]),
			.N(gen[6096]),
			.NE(gen[6097]),

			.O(gen[6190]),
			.E(gen[6192]),

			.SO(gen[6285]),
			.S(gen[6286]),
			.SE(gen[6287]),

			.SELF(gen[6191]),
			.cell_state(gen[6191])
		); 

/******************* CELL 6192 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6192 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6096]),
			.N(gen[6097]),
			.NE(gen[6098]),

			.O(gen[6191]),
			.E(gen[6193]),

			.SO(gen[6286]),
			.S(gen[6287]),
			.SE(gen[6288]),

			.SELF(gen[6192]),
			.cell_state(gen[6192])
		); 

/******************* CELL 6193 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6193 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6097]),
			.N(gen[6098]),
			.NE(gen[6099]),

			.O(gen[6192]),
			.E(gen[6194]),

			.SO(gen[6287]),
			.S(gen[6288]),
			.SE(gen[6289]),

			.SELF(gen[6193]),
			.cell_state(gen[6193])
		); 

/******************* CELL 6194 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6194 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6098]),
			.N(gen[6099]),
			.NE(gen[6100]),

			.O(gen[6193]),
			.E(gen[6195]),

			.SO(gen[6288]),
			.S(gen[6289]),
			.SE(gen[6290]),

			.SELF(gen[6194]),
			.cell_state(gen[6194])
		); 

/******************* CELL 6195 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6195 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6099]),
			.N(gen[6100]),
			.NE(gen[6101]),

			.O(gen[6194]),
			.E(gen[6196]),

			.SO(gen[6289]),
			.S(gen[6290]),
			.SE(gen[6291]),

			.SELF(gen[6195]),
			.cell_state(gen[6195])
		); 

/******************* CELL 6196 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6196 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6100]),
			.N(gen[6101]),
			.NE(gen[6102]),

			.O(gen[6195]),
			.E(gen[6197]),

			.SO(gen[6290]),
			.S(gen[6291]),
			.SE(gen[6292]),

			.SELF(gen[6196]),
			.cell_state(gen[6196])
		); 

/******************* CELL 6197 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6197 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6101]),
			.N(gen[6102]),
			.NE(gen[6103]),

			.O(gen[6196]),
			.E(gen[6198]),

			.SO(gen[6291]),
			.S(gen[6292]),
			.SE(gen[6293]),

			.SELF(gen[6197]),
			.cell_state(gen[6197])
		); 

/******************* CELL 6198 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6198 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6102]),
			.N(gen[6103]),
			.NE(gen[6104]),

			.O(gen[6197]),
			.E(gen[6199]),

			.SO(gen[6292]),
			.S(gen[6293]),
			.SE(gen[6294]),

			.SELF(gen[6198]),
			.cell_state(gen[6198])
		); 

/******************* CELL 6199 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6199 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6103]),
			.N(gen[6104]),
			.NE(gen[6105]),

			.O(gen[6198]),
			.E(gen[6200]),

			.SO(gen[6293]),
			.S(gen[6294]),
			.SE(gen[6295]),

			.SELF(gen[6199]),
			.cell_state(gen[6199])
		); 

/******************* CELL 6200 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6200 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6104]),
			.N(gen[6105]),
			.NE(gen[6106]),

			.O(gen[6199]),
			.E(gen[6201]),

			.SO(gen[6294]),
			.S(gen[6295]),
			.SE(gen[6296]),

			.SELF(gen[6200]),
			.cell_state(gen[6200])
		); 

/******************* CELL 6201 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6201 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6105]),
			.N(gen[6106]),
			.NE(gen[6107]),

			.O(gen[6200]),
			.E(gen[6202]),

			.SO(gen[6295]),
			.S(gen[6296]),
			.SE(gen[6297]),

			.SELF(gen[6201]),
			.cell_state(gen[6201])
		); 

/******************* CELL 6202 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6202 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6106]),
			.N(gen[6107]),
			.NE(gen[6108]),

			.O(gen[6201]),
			.E(gen[6203]),

			.SO(gen[6296]),
			.S(gen[6297]),
			.SE(gen[6298]),

			.SELF(gen[6202]),
			.cell_state(gen[6202])
		); 

/******************* CELL 6203 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6203 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6107]),
			.N(gen[6108]),
			.NE(gen[6109]),

			.O(gen[6202]),
			.E(gen[6204]),

			.SO(gen[6297]),
			.S(gen[6298]),
			.SE(gen[6299]),

			.SELF(gen[6203]),
			.cell_state(gen[6203])
		); 

/******************* CELL 6204 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6204 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6108]),
			.N(gen[6109]),
			.NE(gen[6110]),

			.O(gen[6203]),
			.E(gen[6205]),

			.SO(gen[6298]),
			.S(gen[6299]),
			.SE(gen[6300]),

			.SELF(gen[6204]),
			.cell_state(gen[6204])
		); 

/******************* CELL 6205 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6205 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6109]),
			.N(gen[6110]),
			.NE(gen[6111]),

			.O(gen[6204]),
			.E(gen[6206]),

			.SO(gen[6299]),
			.S(gen[6300]),
			.SE(gen[6301]),

			.SELF(gen[6205]),
			.cell_state(gen[6205])
		); 

/******************* CELL 6206 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6206 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6110]),
			.N(gen[6111]),
			.NE(gen[6112]),

			.O(gen[6205]),
			.E(gen[6207]),

			.SO(gen[6300]),
			.S(gen[6301]),
			.SE(gen[6302]),

			.SELF(gen[6206]),
			.cell_state(gen[6206])
		); 

/******************* CELL 6207 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6207 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6111]),
			.N(gen[6112]),
			.NE(gen[6113]),

			.O(gen[6206]),
			.E(gen[6208]),

			.SO(gen[6301]),
			.S(gen[6302]),
			.SE(gen[6303]),

			.SELF(gen[6207]),
			.cell_state(gen[6207])
		); 

/******************* CELL 6208 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6208 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6112]),
			.N(gen[6113]),
			.NE(gen[6114]),

			.O(gen[6207]),
			.E(gen[6209]),

			.SO(gen[6302]),
			.S(gen[6303]),
			.SE(gen[6304]),

			.SELF(gen[6208]),
			.cell_state(gen[6208])
		); 

/******************* CELL 6209 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6209 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6113]),
			.N(gen[6114]),
			.NE(gen[6115]),

			.O(gen[6208]),
			.E(gen[6210]),

			.SO(gen[6303]),
			.S(gen[6304]),
			.SE(gen[6305]),

			.SELF(gen[6209]),
			.cell_state(gen[6209])
		); 

/******************* CELL 6210 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6210 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6114]),
			.N(gen[6115]),
			.NE(gen[6116]),

			.O(gen[6209]),
			.E(gen[6211]),

			.SO(gen[6304]),
			.S(gen[6305]),
			.SE(gen[6306]),

			.SELF(gen[6210]),
			.cell_state(gen[6210])
		); 

/******************* CELL 6211 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6211 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6115]),
			.N(gen[6116]),
			.NE(gen[6117]),

			.O(gen[6210]),
			.E(gen[6212]),

			.SO(gen[6305]),
			.S(gen[6306]),
			.SE(gen[6307]),

			.SELF(gen[6211]),
			.cell_state(gen[6211])
		); 

/******************* CELL 6212 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6212 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6116]),
			.N(gen[6117]),
			.NE(gen[6118]),

			.O(gen[6211]),
			.E(gen[6213]),

			.SO(gen[6306]),
			.S(gen[6307]),
			.SE(gen[6308]),

			.SELF(gen[6212]),
			.cell_state(gen[6212])
		); 

/******************* CELL 6213 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6213 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6117]),
			.N(gen[6118]),
			.NE(gen[6119]),

			.O(gen[6212]),
			.E(gen[6214]),

			.SO(gen[6307]),
			.S(gen[6308]),
			.SE(gen[6309]),

			.SELF(gen[6213]),
			.cell_state(gen[6213])
		); 

/******************* CELL 6214 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6214 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6118]),
			.N(gen[6119]),
			.NE(gen[6120]),

			.O(gen[6213]),
			.E(gen[6215]),

			.SO(gen[6308]),
			.S(gen[6309]),
			.SE(gen[6310]),

			.SELF(gen[6214]),
			.cell_state(gen[6214])
		); 

/******************* CELL 6215 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6215 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6119]),
			.N(gen[6120]),
			.NE(gen[6121]),

			.O(gen[6214]),
			.E(gen[6216]),

			.SO(gen[6309]),
			.S(gen[6310]),
			.SE(gen[6311]),

			.SELF(gen[6215]),
			.cell_state(gen[6215])
		); 

/******************* CELL 6216 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6216 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6120]),
			.N(gen[6121]),
			.NE(gen[6122]),

			.O(gen[6215]),
			.E(gen[6217]),

			.SO(gen[6310]),
			.S(gen[6311]),
			.SE(gen[6312]),

			.SELF(gen[6216]),
			.cell_state(gen[6216])
		); 

/******************* CELL 6217 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6217 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6121]),
			.N(gen[6122]),
			.NE(gen[6123]),

			.O(gen[6216]),
			.E(gen[6218]),

			.SO(gen[6311]),
			.S(gen[6312]),
			.SE(gen[6313]),

			.SELF(gen[6217]),
			.cell_state(gen[6217])
		); 

/******************* CELL 6218 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6218 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6122]),
			.N(gen[6123]),
			.NE(gen[6124]),

			.O(gen[6217]),
			.E(gen[6219]),

			.SO(gen[6312]),
			.S(gen[6313]),
			.SE(gen[6314]),

			.SELF(gen[6218]),
			.cell_state(gen[6218])
		); 

/******************* CELL 6219 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6219 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6123]),
			.N(gen[6124]),
			.NE(gen[6125]),

			.O(gen[6218]),
			.E(gen[6220]),

			.SO(gen[6313]),
			.S(gen[6314]),
			.SE(gen[6315]),

			.SELF(gen[6219]),
			.cell_state(gen[6219])
		); 

/******************* CELL 6220 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6220 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6124]),
			.N(gen[6125]),
			.NE(gen[6126]),

			.O(gen[6219]),
			.E(gen[6221]),

			.SO(gen[6314]),
			.S(gen[6315]),
			.SE(gen[6316]),

			.SELF(gen[6220]),
			.cell_state(gen[6220])
		); 

/******************* CELL 6221 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6221 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6125]),
			.N(gen[6126]),
			.NE(gen[6127]),

			.O(gen[6220]),
			.E(gen[6222]),

			.SO(gen[6315]),
			.S(gen[6316]),
			.SE(gen[6317]),

			.SELF(gen[6221]),
			.cell_state(gen[6221])
		); 

/******************* CELL 6222 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6222 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6126]),
			.N(gen[6127]),
			.NE(gen[6128]),

			.O(gen[6221]),
			.E(gen[6223]),

			.SO(gen[6316]),
			.S(gen[6317]),
			.SE(gen[6318]),

			.SELF(gen[6222]),
			.cell_state(gen[6222])
		); 

/******************* CELL 6223 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6223 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6127]),
			.N(gen[6128]),
			.NE(gen[6129]),

			.O(gen[6222]),
			.E(gen[6224]),

			.SO(gen[6317]),
			.S(gen[6318]),
			.SE(gen[6319]),

			.SELF(gen[6223]),
			.cell_state(gen[6223])
		); 

/******************* CELL 6224 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6224 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6128]),
			.N(gen[6129]),
			.NE(gen[6130]),

			.O(gen[6223]),
			.E(gen[6225]),

			.SO(gen[6318]),
			.S(gen[6319]),
			.SE(gen[6320]),

			.SELF(gen[6224]),
			.cell_state(gen[6224])
		); 

/******************* CELL 6225 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6225 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6129]),
			.N(gen[6130]),
			.NE(gen[6131]),

			.O(gen[6224]),
			.E(gen[6226]),

			.SO(gen[6319]),
			.S(gen[6320]),
			.SE(gen[6321]),

			.SELF(gen[6225]),
			.cell_state(gen[6225])
		); 

/******************* CELL 6226 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6226 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6130]),
			.N(gen[6131]),
			.NE(gen[6132]),

			.O(gen[6225]),
			.E(gen[6227]),

			.SO(gen[6320]),
			.S(gen[6321]),
			.SE(gen[6322]),

			.SELF(gen[6226]),
			.cell_state(gen[6226])
		); 

/******************* CELL 6227 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6227 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6131]),
			.N(gen[6132]),
			.NE(gen[6133]),

			.O(gen[6226]),
			.E(gen[6228]),

			.SO(gen[6321]),
			.S(gen[6322]),
			.SE(gen[6323]),

			.SELF(gen[6227]),
			.cell_state(gen[6227])
		); 

/******************* CELL 6228 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6228 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6132]),
			.N(gen[6133]),
			.NE(gen[6134]),

			.O(gen[6227]),
			.E(gen[6229]),

			.SO(gen[6322]),
			.S(gen[6323]),
			.SE(gen[6324]),

			.SELF(gen[6228]),
			.cell_state(gen[6228])
		); 

/******************* CELL 6229 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6229 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6133]),
			.N(gen[6134]),
			.NE(gen[6135]),

			.O(gen[6228]),
			.E(gen[6230]),

			.SO(gen[6323]),
			.S(gen[6324]),
			.SE(gen[6325]),

			.SELF(gen[6229]),
			.cell_state(gen[6229])
		); 

/******************* CELL 6230 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6230 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6134]),
			.N(gen[6135]),
			.NE(gen[6136]),

			.O(gen[6229]),
			.E(gen[6231]),

			.SO(gen[6324]),
			.S(gen[6325]),
			.SE(gen[6326]),

			.SELF(gen[6230]),
			.cell_state(gen[6230])
		); 

/******************* CELL 6231 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6231 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6135]),
			.N(gen[6136]),
			.NE(gen[6137]),

			.O(gen[6230]),
			.E(gen[6232]),

			.SO(gen[6325]),
			.S(gen[6326]),
			.SE(gen[6327]),

			.SELF(gen[6231]),
			.cell_state(gen[6231])
		); 

/******************* CELL 6232 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6232 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6136]),
			.N(gen[6137]),
			.NE(gen[6138]),

			.O(gen[6231]),
			.E(gen[6233]),

			.SO(gen[6326]),
			.S(gen[6327]),
			.SE(gen[6328]),

			.SELF(gen[6232]),
			.cell_state(gen[6232])
		); 

/******************* CELL 6233 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6233 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6137]),
			.N(gen[6138]),
			.NE(gen[6139]),

			.O(gen[6232]),
			.E(gen[6234]),

			.SO(gen[6327]),
			.S(gen[6328]),
			.SE(gen[6329]),

			.SELF(gen[6233]),
			.cell_state(gen[6233])
		); 

/******************* CELL 6234 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6234 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6138]),
			.N(gen[6139]),
			.NE(gen[6140]),

			.O(gen[6233]),
			.E(gen[6235]),

			.SO(gen[6328]),
			.S(gen[6329]),
			.SE(gen[6330]),

			.SELF(gen[6234]),
			.cell_state(gen[6234])
		); 

/******************* CELL 6235 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6235 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6139]),
			.N(gen[6140]),
			.NE(gen[6141]),

			.O(gen[6234]),
			.E(gen[6236]),

			.SO(gen[6329]),
			.S(gen[6330]),
			.SE(gen[6331]),

			.SELF(gen[6235]),
			.cell_state(gen[6235])
		); 

/******************* CELL 6236 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6236 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6140]),
			.N(gen[6141]),
			.NE(gen[6142]),

			.O(gen[6235]),
			.E(gen[6237]),

			.SO(gen[6330]),
			.S(gen[6331]),
			.SE(gen[6332]),

			.SELF(gen[6236]),
			.cell_state(gen[6236])
		); 

/******************* CELL 6237 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6237 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6141]),
			.N(gen[6142]),
			.NE(gen[6143]),

			.O(gen[6236]),
			.E(gen[6238]),

			.SO(gen[6331]),
			.S(gen[6332]),
			.SE(gen[6333]),

			.SELF(gen[6237]),
			.cell_state(gen[6237])
		); 

/******************* CELL 6238 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6238 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6142]),
			.N(gen[6143]),
			.NE(gen[6144]),

			.O(gen[6237]),
			.E(gen[6239]),

			.SO(gen[6332]),
			.S(gen[6333]),
			.SE(gen[6334]),

			.SELF(gen[6238]),
			.cell_state(gen[6238])
		); 

/******************* CELL 6239 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6239 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6143]),
			.N(gen[6144]),
			.NE(gen[6145]),

			.O(gen[6238]),
			.E(gen[6240]),

			.SO(gen[6333]),
			.S(gen[6334]),
			.SE(gen[6335]),

			.SELF(gen[6239]),
			.cell_state(gen[6239])
		); 

/******************* CELL 6240 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6240 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6144]),
			.N(gen[6145]),
			.NE(gen[6146]),

			.O(gen[6239]),
			.E(gen[6241]),

			.SO(gen[6334]),
			.S(gen[6335]),
			.SE(gen[6336]),

			.SELF(gen[6240]),
			.cell_state(gen[6240])
		); 

/******************* CELL 6241 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6241 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6145]),
			.N(gen[6146]),
			.NE(gen[6147]),

			.O(gen[6240]),
			.E(gen[6242]),

			.SO(gen[6335]),
			.S(gen[6336]),
			.SE(gen[6337]),

			.SELF(gen[6241]),
			.cell_state(gen[6241])
		); 

/******************* CELL 6242 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6242 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6146]),
			.N(gen[6147]),
			.NE(gen[6148]),

			.O(gen[6241]),
			.E(gen[6243]),

			.SO(gen[6336]),
			.S(gen[6337]),
			.SE(gen[6338]),

			.SELF(gen[6242]),
			.cell_state(gen[6242])
		); 

/******************* CELL 6243 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6243 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6147]),
			.N(gen[6148]),
			.NE(gen[6149]),

			.O(gen[6242]),
			.E(gen[6244]),

			.SO(gen[6337]),
			.S(gen[6338]),
			.SE(gen[6339]),

			.SELF(gen[6243]),
			.cell_state(gen[6243])
		); 

/******************* CELL 6244 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6244 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6148]),
			.N(gen[6149]),
			.NE(gen[6150]),

			.O(gen[6243]),
			.E(gen[6245]),

			.SO(gen[6338]),
			.S(gen[6339]),
			.SE(gen[6340]),

			.SELF(gen[6244]),
			.cell_state(gen[6244])
		); 

/******************* CELL 6245 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6245 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6149]),
			.N(gen[6150]),
			.NE(gen[6151]),

			.O(gen[6244]),
			.E(gen[6246]),

			.SO(gen[6339]),
			.S(gen[6340]),
			.SE(gen[6341]),

			.SELF(gen[6245]),
			.cell_state(gen[6245])
		); 

/******************* CELL 6246 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6246 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6150]),
			.N(gen[6151]),
			.NE(gen[6152]),

			.O(gen[6245]),
			.E(gen[6247]),

			.SO(gen[6340]),
			.S(gen[6341]),
			.SE(gen[6342]),

			.SELF(gen[6246]),
			.cell_state(gen[6246])
		); 

/******************* CELL 6247 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6247 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6151]),
			.N(gen[6152]),
			.NE(gen[6153]),

			.O(gen[6246]),
			.E(gen[6248]),

			.SO(gen[6341]),
			.S(gen[6342]),
			.SE(gen[6343]),

			.SELF(gen[6247]),
			.cell_state(gen[6247])
		); 

/******************* CELL 6248 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6248 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6152]),
			.N(gen[6153]),
			.NE(gen[6154]),

			.O(gen[6247]),
			.E(gen[6249]),

			.SO(gen[6342]),
			.S(gen[6343]),
			.SE(gen[6344]),

			.SELF(gen[6248]),
			.cell_state(gen[6248])
		); 

/******************* CELL 6249 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6249 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6153]),
			.N(gen[6154]),
			.NE(gen[6155]),

			.O(gen[6248]),
			.E(gen[6250]),

			.SO(gen[6343]),
			.S(gen[6344]),
			.SE(gen[6345]),

			.SELF(gen[6249]),
			.cell_state(gen[6249])
		); 

/******************* CELL 6250 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6250 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6154]),
			.N(gen[6155]),
			.NE(gen[6156]),

			.O(gen[6249]),
			.E(gen[6251]),

			.SO(gen[6344]),
			.S(gen[6345]),
			.SE(gen[6346]),

			.SELF(gen[6250]),
			.cell_state(gen[6250])
		); 

/******************* CELL 6251 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6251 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6155]),
			.N(gen[6156]),
			.NE(gen[6157]),

			.O(gen[6250]),
			.E(gen[6252]),

			.SO(gen[6345]),
			.S(gen[6346]),
			.SE(gen[6347]),

			.SELF(gen[6251]),
			.cell_state(gen[6251])
		); 

/******************* CELL 6252 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6252 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6156]),
			.N(gen[6157]),
			.NE(gen[6158]),

			.O(gen[6251]),
			.E(gen[6253]),

			.SO(gen[6346]),
			.S(gen[6347]),
			.SE(gen[6348]),

			.SELF(gen[6252]),
			.cell_state(gen[6252])
		); 

/******************* CELL 6253 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6253 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6157]),
			.N(gen[6158]),
			.NE(gen[6159]),

			.O(gen[6252]),
			.E(gen[6254]),

			.SO(gen[6347]),
			.S(gen[6348]),
			.SE(gen[6349]),

			.SELF(gen[6253]),
			.cell_state(gen[6253])
		); 

/******************* CELL 6254 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6254 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6158]),
			.N(gen[6159]),
			.NE(gen[6160]),

			.O(gen[6253]),
			.E(gen[6255]),

			.SO(gen[6348]),
			.S(gen[6349]),
			.SE(gen[6350]),

			.SELF(gen[6254]),
			.cell_state(gen[6254])
		); 

/******************* CELL 6255 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6255 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6159]),
			.N(gen[6160]),
			.NE(gen[6161]),

			.O(gen[6254]),
			.E(gen[6256]),

			.SO(gen[6349]),
			.S(gen[6350]),
			.SE(gen[6351]),

			.SELF(gen[6255]),
			.cell_state(gen[6255])
		); 

/******************* CELL 6256 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6256 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6160]),
			.N(gen[6161]),
			.NE(gen[6162]),

			.O(gen[6255]),
			.E(gen[6257]),

			.SO(gen[6350]),
			.S(gen[6351]),
			.SE(gen[6352]),

			.SELF(gen[6256]),
			.cell_state(gen[6256])
		); 

/******************* CELL 6257 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6257 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6161]),
			.N(gen[6162]),
			.NE(gen[6163]),

			.O(gen[6256]),
			.E(gen[6258]),

			.SO(gen[6351]),
			.S(gen[6352]),
			.SE(gen[6353]),

			.SELF(gen[6257]),
			.cell_state(gen[6257])
		); 

/******************* CELL 6258 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6258 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6162]),
			.N(gen[6163]),
			.NE(gen[6164]),

			.O(gen[6257]),
			.E(gen[6259]),

			.SO(gen[6352]),
			.S(gen[6353]),
			.SE(gen[6354]),

			.SELF(gen[6258]),
			.cell_state(gen[6258])
		); 

/******************* CELL 6259 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6259 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6163]),
			.N(gen[6164]),
			.NE(gen[6165]),

			.O(gen[6258]),
			.E(gen[6260]),

			.SO(gen[6353]),
			.S(gen[6354]),
			.SE(gen[6355]),

			.SELF(gen[6259]),
			.cell_state(gen[6259])
		); 

/******************* CELL 6260 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6260 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6164]),
			.N(gen[6165]),
			.NE(gen[6166]),

			.O(gen[6259]),
			.E(gen[6261]),

			.SO(gen[6354]),
			.S(gen[6355]),
			.SE(gen[6356]),

			.SELF(gen[6260]),
			.cell_state(gen[6260])
		); 

/******************* CELL 6261 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6261 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6165]),
			.N(gen[6166]),
			.NE(gen[6167]),

			.O(gen[6260]),
			.E(gen[6262]),

			.SO(gen[6355]),
			.S(gen[6356]),
			.SE(gen[6357]),

			.SELF(gen[6261]),
			.cell_state(gen[6261])
		); 

/******************* CELL 6262 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6262 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6166]),
			.N(gen[6167]),
			.NE(gen[6168]),

			.O(gen[6261]),
			.E(gen[6263]),

			.SO(gen[6356]),
			.S(gen[6357]),
			.SE(gen[6358]),

			.SELF(gen[6262]),
			.cell_state(gen[6262])
		); 

/******************* CELL 6263 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6263 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6167]),
			.N(gen[6168]),
			.NE(gen[6169]),

			.O(gen[6262]),
			.E(gen[6264]),

			.SO(gen[6357]),
			.S(gen[6358]),
			.SE(gen[6359]),

			.SELF(gen[6263]),
			.cell_state(gen[6263])
		); 

/******************* CELL 6264 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6264 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6168]),
			.N(gen[6169]),
			.NE(gen[6170]),

			.O(gen[6263]),
			.E(gen[6265]),

			.SO(gen[6358]),
			.S(gen[6359]),
			.SE(gen[6360]),

			.SELF(gen[6264]),
			.cell_state(gen[6264])
		); 

/******************* CELL 6265 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6265 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6169]),
			.N(gen[6170]),
			.NE(gen[6171]),

			.O(gen[6264]),
			.E(gen[6266]),

			.SO(gen[6359]),
			.S(gen[6360]),
			.SE(gen[6361]),

			.SELF(gen[6265]),
			.cell_state(gen[6265])
		); 

/******************* CELL 6266 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6266 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6170]),
			.N(gen[6171]),
			.NE(gen[6172]),

			.O(gen[6265]),
			.E(gen[6267]),

			.SO(gen[6360]),
			.S(gen[6361]),
			.SE(gen[6362]),

			.SELF(gen[6266]),
			.cell_state(gen[6266])
		); 

/******************* CELL 6267 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6267 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6171]),
			.N(gen[6172]),
			.NE(gen[6173]),

			.O(gen[6266]),
			.E(gen[6268]),

			.SO(gen[6361]),
			.S(gen[6362]),
			.SE(gen[6363]),

			.SELF(gen[6267]),
			.cell_state(gen[6267])
		); 

/******************* CELL 6268 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6268 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6172]),
			.N(gen[6173]),
			.NE(gen[6174]),

			.O(gen[6267]),
			.E(gen[6269]),

			.SO(gen[6362]),
			.S(gen[6363]),
			.SE(gen[6364]),

			.SELF(gen[6268]),
			.cell_state(gen[6268])
		); 

/******************* CELL 6269 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6269 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6173]),
			.N(gen[6174]),
			.NE(gen[6173]),

			.O(gen[6268]),
			.E(gen[6268]),

			.SO(gen[6363]),
			.S(gen[6364]),
			.SE(gen[6363]),

			.SELF(gen[6269]),
			.cell_state(gen[6269])
		); 

/******************* CELL 6270 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6270 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6176]),
			.N(gen[6175]),
			.NE(gen[6176]),

			.O(gen[6271]),
			.E(gen[6271]),

			.SO(gen[6366]),
			.S(gen[6365]),
			.SE(gen[6366]),

			.SELF(gen[6270]),
			.cell_state(gen[6270])
		); 

/******************* CELL 6271 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6271 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6175]),
			.N(gen[6176]),
			.NE(gen[6177]),

			.O(gen[6270]),
			.E(gen[6272]),

			.SO(gen[6365]),
			.S(gen[6366]),
			.SE(gen[6367]),

			.SELF(gen[6271]),
			.cell_state(gen[6271])
		); 

/******************* CELL 6272 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6272 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6176]),
			.N(gen[6177]),
			.NE(gen[6178]),

			.O(gen[6271]),
			.E(gen[6273]),

			.SO(gen[6366]),
			.S(gen[6367]),
			.SE(gen[6368]),

			.SELF(gen[6272]),
			.cell_state(gen[6272])
		); 

/******************* CELL 6273 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6273 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6177]),
			.N(gen[6178]),
			.NE(gen[6179]),

			.O(gen[6272]),
			.E(gen[6274]),

			.SO(gen[6367]),
			.S(gen[6368]),
			.SE(gen[6369]),

			.SELF(gen[6273]),
			.cell_state(gen[6273])
		); 

/******************* CELL 6274 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6274 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6178]),
			.N(gen[6179]),
			.NE(gen[6180]),

			.O(gen[6273]),
			.E(gen[6275]),

			.SO(gen[6368]),
			.S(gen[6369]),
			.SE(gen[6370]),

			.SELF(gen[6274]),
			.cell_state(gen[6274])
		); 

/******************* CELL 6275 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6275 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6179]),
			.N(gen[6180]),
			.NE(gen[6181]),

			.O(gen[6274]),
			.E(gen[6276]),

			.SO(gen[6369]),
			.S(gen[6370]),
			.SE(gen[6371]),

			.SELF(gen[6275]),
			.cell_state(gen[6275])
		); 

/******************* CELL 6276 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6276 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6180]),
			.N(gen[6181]),
			.NE(gen[6182]),

			.O(gen[6275]),
			.E(gen[6277]),

			.SO(gen[6370]),
			.S(gen[6371]),
			.SE(gen[6372]),

			.SELF(gen[6276]),
			.cell_state(gen[6276])
		); 

/******************* CELL 6277 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6277 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6181]),
			.N(gen[6182]),
			.NE(gen[6183]),

			.O(gen[6276]),
			.E(gen[6278]),

			.SO(gen[6371]),
			.S(gen[6372]),
			.SE(gen[6373]),

			.SELF(gen[6277]),
			.cell_state(gen[6277])
		); 

/******************* CELL 6278 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6278 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6182]),
			.N(gen[6183]),
			.NE(gen[6184]),

			.O(gen[6277]),
			.E(gen[6279]),

			.SO(gen[6372]),
			.S(gen[6373]),
			.SE(gen[6374]),

			.SELF(gen[6278]),
			.cell_state(gen[6278])
		); 

/******************* CELL 6279 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6279 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6183]),
			.N(gen[6184]),
			.NE(gen[6185]),

			.O(gen[6278]),
			.E(gen[6280]),

			.SO(gen[6373]),
			.S(gen[6374]),
			.SE(gen[6375]),

			.SELF(gen[6279]),
			.cell_state(gen[6279])
		); 

/******************* CELL 6280 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6280 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6184]),
			.N(gen[6185]),
			.NE(gen[6186]),

			.O(gen[6279]),
			.E(gen[6281]),

			.SO(gen[6374]),
			.S(gen[6375]),
			.SE(gen[6376]),

			.SELF(gen[6280]),
			.cell_state(gen[6280])
		); 

/******************* CELL 6281 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6281 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6185]),
			.N(gen[6186]),
			.NE(gen[6187]),

			.O(gen[6280]),
			.E(gen[6282]),

			.SO(gen[6375]),
			.S(gen[6376]),
			.SE(gen[6377]),

			.SELF(gen[6281]),
			.cell_state(gen[6281])
		); 

/******************* CELL 6282 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6282 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6186]),
			.N(gen[6187]),
			.NE(gen[6188]),

			.O(gen[6281]),
			.E(gen[6283]),

			.SO(gen[6376]),
			.S(gen[6377]),
			.SE(gen[6378]),

			.SELF(gen[6282]),
			.cell_state(gen[6282])
		); 

/******************* CELL 6283 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6283 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6187]),
			.N(gen[6188]),
			.NE(gen[6189]),

			.O(gen[6282]),
			.E(gen[6284]),

			.SO(gen[6377]),
			.S(gen[6378]),
			.SE(gen[6379]),

			.SELF(gen[6283]),
			.cell_state(gen[6283])
		); 

/******************* CELL 6284 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6284 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6188]),
			.N(gen[6189]),
			.NE(gen[6190]),

			.O(gen[6283]),
			.E(gen[6285]),

			.SO(gen[6378]),
			.S(gen[6379]),
			.SE(gen[6380]),

			.SELF(gen[6284]),
			.cell_state(gen[6284])
		); 

/******************* CELL 6285 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6285 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6189]),
			.N(gen[6190]),
			.NE(gen[6191]),

			.O(gen[6284]),
			.E(gen[6286]),

			.SO(gen[6379]),
			.S(gen[6380]),
			.SE(gen[6381]),

			.SELF(gen[6285]),
			.cell_state(gen[6285])
		); 

/******************* CELL 6286 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6286 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6190]),
			.N(gen[6191]),
			.NE(gen[6192]),

			.O(gen[6285]),
			.E(gen[6287]),

			.SO(gen[6380]),
			.S(gen[6381]),
			.SE(gen[6382]),

			.SELF(gen[6286]),
			.cell_state(gen[6286])
		); 

/******************* CELL 6287 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6287 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6191]),
			.N(gen[6192]),
			.NE(gen[6193]),

			.O(gen[6286]),
			.E(gen[6288]),

			.SO(gen[6381]),
			.S(gen[6382]),
			.SE(gen[6383]),

			.SELF(gen[6287]),
			.cell_state(gen[6287])
		); 

/******************* CELL 6288 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6288 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6192]),
			.N(gen[6193]),
			.NE(gen[6194]),

			.O(gen[6287]),
			.E(gen[6289]),

			.SO(gen[6382]),
			.S(gen[6383]),
			.SE(gen[6384]),

			.SELF(gen[6288]),
			.cell_state(gen[6288])
		); 

/******************* CELL 6289 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6289 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6193]),
			.N(gen[6194]),
			.NE(gen[6195]),

			.O(gen[6288]),
			.E(gen[6290]),

			.SO(gen[6383]),
			.S(gen[6384]),
			.SE(gen[6385]),

			.SELF(gen[6289]),
			.cell_state(gen[6289])
		); 

/******************* CELL 6290 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6290 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6194]),
			.N(gen[6195]),
			.NE(gen[6196]),

			.O(gen[6289]),
			.E(gen[6291]),

			.SO(gen[6384]),
			.S(gen[6385]),
			.SE(gen[6386]),

			.SELF(gen[6290]),
			.cell_state(gen[6290])
		); 

/******************* CELL 6291 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6291 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6195]),
			.N(gen[6196]),
			.NE(gen[6197]),

			.O(gen[6290]),
			.E(gen[6292]),

			.SO(gen[6385]),
			.S(gen[6386]),
			.SE(gen[6387]),

			.SELF(gen[6291]),
			.cell_state(gen[6291])
		); 

/******************* CELL 6292 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6292 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6196]),
			.N(gen[6197]),
			.NE(gen[6198]),

			.O(gen[6291]),
			.E(gen[6293]),

			.SO(gen[6386]),
			.S(gen[6387]),
			.SE(gen[6388]),

			.SELF(gen[6292]),
			.cell_state(gen[6292])
		); 

/******************* CELL 6293 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6293 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6197]),
			.N(gen[6198]),
			.NE(gen[6199]),

			.O(gen[6292]),
			.E(gen[6294]),

			.SO(gen[6387]),
			.S(gen[6388]),
			.SE(gen[6389]),

			.SELF(gen[6293]),
			.cell_state(gen[6293])
		); 

/******************* CELL 6294 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6294 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6198]),
			.N(gen[6199]),
			.NE(gen[6200]),

			.O(gen[6293]),
			.E(gen[6295]),

			.SO(gen[6388]),
			.S(gen[6389]),
			.SE(gen[6390]),

			.SELF(gen[6294]),
			.cell_state(gen[6294])
		); 

/******************* CELL 6295 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6295 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6199]),
			.N(gen[6200]),
			.NE(gen[6201]),

			.O(gen[6294]),
			.E(gen[6296]),

			.SO(gen[6389]),
			.S(gen[6390]),
			.SE(gen[6391]),

			.SELF(gen[6295]),
			.cell_state(gen[6295])
		); 

/******************* CELL 6296 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6296 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6200]),
			.N(gen[6201]),
			.NE(gen[6202]),

			.O(gen[6295]),
			.E(gen[6297]),

			.SO(gen[6390]),
			.S(gen[6391]),
			.SE(gen[6392]),

			.SELF(gen[6296]),
			.cell_state(gen[6296])
		); 

/******************* CELL 6297 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6297 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6201]),
			.N(gen[6202]),
			.NE(gen[6203]),

			.O(gen[6296]),
			.E(gen[6298]),

			.SO(gen[6391]),
			.S(gen[6392]),
			.SE(gen[6393]),

			.SELF(gen[6297]),
			.cell_state(gen[6297])
		); 

/******************* CELL 6298 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6298 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6202]),
			.N(gen[6203]),
			.NE(gen[6204]),

			.O(gen[6297]),
			.E(gen[6299]),

			.SO(gen[6392]),
			.S(gen[6393]),
			.SE(gen[6394]),

			.SELF(gen[6298]),
			.cell_state(gen[6298])
		); 

/******************* CELL 6299 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6299 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6203]),
			.N(gen[6204]),
			.NE(gen[6205]),

			.O(gen[6298]),
			.E(gen[6300]),

			.SO(gen[6393]),
			.S(gen[6394]),
			.SE(gen[6395]),

			.SELF(gen[6299]),
			.cell_state(gen[6299])
		); 

/******************* CELL 6300 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6300 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6204]),
			.N(gen[6205]),
			.NE(gen[6206]),

			.O(gen[6299]),
			.E(gen[6301]),

			.SO(gen[6394]),
			.S(gen[6395]),
			.SE(gen[6396]),

			.SELF(gen[6300]),
			.cell_state(gen[6300])
		); 

/******************* CELL 6301 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6301 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6205]),
			.N(gen[6206]),
			.NE(gen[6207]),

			.O(gen[6300]),
			.E(gen[6302]),

			.SO(gen[6395]),
			.S(gen[6396]),
			.SE(gen[6397]),

			.SELF(gen[6301]),
			.cell_state(gen[6301])
		); 

/******************* CELL 6302 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6302 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6206]),
			.N(gen[6207]),
			.NE(gen[6208]),

			.O(gen[6301]),
			.E(gen[6303]),

			.SO(gen[6396]),
			.S(gen[6397]),
			.SE(gen[6398]),

			.SELF(gen[6302]),
			.cell_state(gen[6302])
		); 

/******************* CELL 6303 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6303 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6207]),
			.N(gen[6208]),
			.NE(gen[6209]),

			.O(gen[6302]),
			.E(gen[6304]),

			.SO(gen[6397]),
			.S(gen[6398]),
			.SE(gen[6399]),

			.SELF(gen[6303]),
			.cell_state(gen[6303])
		); 

/******************* CELL 6304 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6304 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6208]),
			.N(gen[6209]),
			.NE(gen[6210]),

			.O(gen[6303]),
			.E(gen[6305]),

			.SO(gen[6398]),
			.S(gen[6399]),
			.SE(gen[6400]),

			.SELF(gen[6304]),
			.cell_state(gen[6304])
		); 

/******************* CELL 6305 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6305 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6209]),
			.N(gen[6210]),
			.NE(gen[6211]),

			.O(gen[6304]),
			.E(gen[6306]),

			.SO(gen[6399]),
			.S(gen[6400]),
			.SE(gen[6401]),

			.SELF(gen[6305]),
			.cell_state(gen[6305])
		); 

/******************* CELL 6306 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6306 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6210]),
			.N(gen[6211]),
			.NE(gen[6212]),

			.O(gen[6305]),
			.E(gen[6307]),

			.SO(gen[6400]),
			.S(gen[6401]),
			.SE(gen[6402]),

			.SELF(gen[6306]),
			.cell_state(gen[6306])
		); 

/******************* CELL 6307 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6307 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6211]),
			.N(gen[6212]),
			.NE(gen[6213]),

			.O(gen[6306]),
			.E(gen[6308]),

			.SO(gen[6401]),
			.S(gen[6402]),
			.SE(gen[6403]),

			.SELF(gen[6307]),
			.cell_state(gen[6307])
		); 

/******************* CELL 6308 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6308 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6212]),
			.N(gen[6213]),
			.NE(gen[6214]),

			.O(gen[6307]),
			.E(gen[6309]),

			.SO(gen[6402]),
			.S(gen[6403]),
			.SE(gen[6404]),

			.SELF(gen[6308]),
			.cell_state(gen[6308])
		); 

/******************* CELL 6309 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6309 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6213]),
			.N(gen[6214]),
			.NE(gen[6215]),

			.O(gen[6308]),
			.E(gen[6310]),

			.SO(gen[6403]),
			.S(gen[6404]),
			.SE(gen[6405]),

			.SELF(gen[6309]),
			.cell_state(gen[6309])
		); 

/******************* CELL 6310 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6310 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6214]),
			.N(gen[6215]),
			.NE(gen[6216]),

			.O(gen[6309]),
			.E(gen[6311]),

			.SO(gen[6404]),
			.S(gen[6405]),
			.SE(gen[6406]),

			.SELF(gen[6310]),
			.cell_state(gen[6310])
		); 

/******************* CELL 6311 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6311 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6215]),
			.N(gen[6216]),
			.NE(gen[6217]),

			.O(gen[6310]),
			.E(gen[6312]),

			.SO(gen[6405]),
			.S(gen[6406]),
			.SE(gen[6407]),

			.SELF(gen[6311]),
			.cell_state(gen[6311])
		); 

/******************* CELL 6312 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6312 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6216]),
			.N(gen[6217]),
			.NE(gen[6218]),

			.O(gen[6311]),
			.E(gen[6313]),

			.SO(gen[6406]),
			.S(gen[6407]),
			.SE(gen[6408]),

			.SELF(gen[6312]),
			.cell_state(gen[6312])
		); 

/******************* CELL 6313 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6313 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6217]),
			.N(gen[6218]),
			.NE(gen[6219]),

			.O(gen[6312]),
			.E(gen[6314]),

			.SO(gen[6407]),
			.S(gen[6408]),
			.SE(gen[6409]),

			.SELF(gen[6313]),
			.cell_state(gen[6313])
		); 

/******************* CELL 6314 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6314 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6218]),
			.N(gen[6219]),
			.NE(gen[6220]),

			.O(gen[6313]),
			.E(gen[6315]),

			.SO(gen[6408]),
			.S(gen[6409]),
			.SE(gen[6410]),

			.SELF(gen[6314]),
			.cell_state(gen[6314])
		); 

/******************* CELL 6315 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6315 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6219]),
			.N(gen[6220]),
			.NE(gen[6221]),

			.O(gen[6314]),
			.E(gen[6316]),

			.SO(gen[6409]),
			.S(gen[6410]),
			.SE(gen[6411]),

			.SELF(gen[6315]),
			.cell_state(gen[6315])
		); 

/******************* CELL 6316 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6316 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6220]),
			.N(gen[6221]),
			.NE(gen[6222]),

			.O(gen[6315]),
			.E(gen[6317]),

			.SO(gen[6410]),
			.S(gen[6411]),
			.SE(gen[6412]),

			.SELF(gen[6316]),
			.cell_state(gen[6316])
		); 

/******************* CELL 6317 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6317 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6221]),
			.N(gen[6222]),
			.NE(gen[6223]),

			.O(gen[6316]),
			.E(gen[6318]),

			.SO(gen[6411]),
			.S(gen[6412]),
			.SE(gen[6413]),

			.SELF(gen[6317]),
			.cell_state(gen[6317])
		); 

/******************* CELL 6318 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6318 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6222]),
			.N(gen[6223]),
			.NE(gen[6224]),

			.O(gen[6317]),
			.E(gen[6319]),

			.SO(gen[6412]),
			.S(gen[6413]),
			.SE(gen[6414]),

			.SELF(gen[6318]),
			.cell_state(gen[6318])
		); 

/******************* CELL 6319 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6319 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6223]),
			.N(gen[6224]),
			.NE(gen[6225]),

			.O(gen[6318]),
			.E(gen[6320]),

			.SO(gen[6413]),
			.S(gen[6414]),
			.SE(gen[6415]),

			.SELF(gen[6319]),
			.cell_state(gen[6319])
		); 

/******************* CELL 6320 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6320 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6224]),
			.N(gen[6225]),
			.NE(gen[6226]),

			.O(gen[6319]),
			.E(gen[6321]),

			.SO(gen[6414]),
			.S(gen[6415]),
			.SE(gen[6416]),

			.SELF(gen[6320]),
			.cell_state(gen[6320])
		); 

/******************* CELL 6321 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6321 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6225]),
			.N(gen[6226]),
			.NE(gen[6227]),

			.O(gen[6320]),
			.E(gen[6322]),

			.SO(gen[6415]),
			.S(gen[6416]),
			.SE(gen[6417]),

			.SELF(gen[6321]),
			.cell_state(gen[6321])
		); 

/******************* CELL 6322 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6322 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6226]),
			.N(gen[6227]),
			.NE(gen[6228]),

			.O(gen[6321]),
			.E(gen[6323]),

			.SO(gen[6416]),
			.S(gen[6417]),
			.SE(gen[6418]),

			.SELF(gen[6322]),
			.cell_state(gen[6322])
		); 

/******************* CELL 6323 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6323 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6227]),
			.N(gen[6228]),
			.NE(gen[6229]),

			.O(gen[6322]),
			.E(gen[6324]),

			.SO(gen[6417]),
			.S(gen[6418]),
			.SE(gen[6419]),

			.SELF(gen[6323]),
			.cell_state(gen[6323])
		); 

/******************* CELL 6324 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6324 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6228]),
			.N(gen[6229]),
			.NE(gen[6230]),

			.O(gen[6323]),
			.E(gen[6325]),

			.SO(gen[6418]),
			.S(gen[6419]),
			.SE(gen[6420]),

			.SELF(gen[6324]),
			.cell_state(gen[6324])
		); 

/******************* CELL 6325 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6325 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6229]),
			.N(gen[6230]),
			.NE(gen[6231]),

			.O(gen[6324]),
			.E(gen[6326]),

			.SO(gen[6419]),
			.S(gen[6420]),
			.SE(gen[6421]),

			.SELF(gen[6325]),
			.cell_state(gen[6325])
		); 

/******************* CELL 6326 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6326 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6230]),
			.N(gen[6231]),
			.NE(gen[6232]),

			.O(gen[6325]),
			.E(gen[6327]),

			.SO(gen[6420]),
			.S(gen[6421]),
			.SE(gen[6422]),

			.SELF(gen[6326]),
			.cell_state(gen[6326])
		); 

/******************* CELL 6327 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6327 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6231]),
			.N(gen[6232]),
			.NE(gen[6233]),

			.O(gen[6326]),
			.E(gen[6328]),

			.SO(gen[6421]),
			.S(gen[6422]),
			.SE(gen[6423]),

			.SELF(gen[6327]),
			.cell_state(gen[6327])
		); 

/******************* CELL 6328 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6328 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6232]),
			.N(gen[6233]),
			.NE(gen[6234]),

			.O(gen[6327]),
			.E(gen[6329]),

			.SO(gen[6422]),
			.S(gen[6423]),
			.SE(gen[6424]),

			.SELF(gen[6328]),
			.cell_state(gen[6328])
		); 

/******************* CELL 6329 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6329 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6233]),
			.N(gen[6234]),
			.NE(gen[6235]),

			.O(gen[6328]),
			.E(gen[6330]),

			.SO(gen[6423]),
			.S(gen[6424]),
			.SE(gen[6425]),

			.SELF(gen[6329]),
			.cell_state(gen[6329])
		); 

/******************* CELL 6330 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6330 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6234]),
			.N(gen[6235]),
			.NE(gen[6236]),

			.O(gen[6329]),
			.E(gen[6331]),

			.SO(gen[6424]),
			.S(gen[6425]),
			.SE(gen[6426]),

			.SELF(gen[6330]),
			.cell_state(gen[6330])
		); 

/******************* CELL 6331 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6331 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6235]),
			.N(gen[6236]),
			.NE(gen[6237]),

			.O(gen[6330]),
			.E(gen[6332]),

			.SO(gen[6425]),
			.S(gen[6426]),
			.SE(gen[6427]),

			.SELF(gen[6331]),
			.cell_state(gen[6331])
		); 

/******************* CELL 6332 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6332 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6236]),
			.N(gen[6237]),
			.NE(gen[6238]),

			.O(gen[6331]),
			.E(gen[6333]),

			.SO(gen[6426]),
			.S(gen[6427]),
			.SE(gen[6428]),

			.SELF(gen[6332]),
			.cell_state(gen[6332])
		); 

/******************* CELL 6333 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6333 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6237]),
			.N(gen[6238]),
			.NE(gen[6239]),

			.O(gen[6332]),
			.E(gen[6334]),

			.SO(gen[6427]),
			.S(gen[6428]),
			.SE(gen[6429]),

			.SELF(gen[6333]),
			.cell_state(gen[6333])
		); 

/******************* CELL 6334 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6334 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6238]),
			.N(gen[6239]),
			.NE(gen[6240]),

			.O(gen[6333]),
			.E(gen[6335]),

			.SO(gen[6428]),
			.S(gen[6429]),
			.SE(gen[6430]),

			.SELF(gen[6334]),
			.cell_state(gen[6334])
		); 

/******************* CELL 6335 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6335 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6239]),
			.N(gen[6240]),
			.NE(gen[6241]),

			.O(gen[6334]),
			.E(gen[6336]),

			.SO(gen[6429]),
			.S(gen[6430]),
			.SE(gen[6431]),

			.SELF(gen[6335]),
			.cell_state(gen[6335])
		); 

/******************* CELL 6336 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6336 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6240]),
			.N(gen[6241]),
			.NE(gen[6242]),

			.O(gen[6335]),
			.E(gen[6337]),

			.SO(gen[6430]),
			.S(gen[6431]),
			.SE(gen[6432]),

			.SELF(gen[6336]),
			.cell_state(gen[6336])
		); 

/******************* CELL 6337 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6337 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6241]),
			.N(gen[6242]),
			.NE(gen[6243]),

			.O(gen[6336]),
			.E(gen[6338]),

			.SO(gen[6431]),
			.S(gen[6432]),
			.SE(gen[6433]),

			.SELF(gen[6337]),
			.cell_state(gen[6337])
		); 

/******************* CELL 6338 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6338 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6242]),
			.N(gen[6243]),
			.NE(gen[6244]),

			.O(gen[6337]),
			.E(gen[6339]),

			.SO(gen[6432]),
			.S(gen[6433]),
			.SE(gen[6434]),

			.SELF(gen[6338]),
			.cell_state(gen[6338])
		); 

/******************* CELL 6339 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6339 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6243]),
			.N(gen[6244]),
			.NE(gen[6245]),

			.O(gen[6338]),
			.E(gen[6340]),

			.SO(gen[6433]),
			.S(gen[6434]),
			.SE(gen[6435]),

			.SELF(gen[6339]),
			.cell_state(gen[6339])
		); 

/******************* CELL 6340 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6340 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6244]),
			.N(gen[6245]),
			.NE(gen[6246]),

			.O(gen[6339]),
			.E(gen[6341]),

			.SO(gen[6434]),
			.S(gen[6435]),
			.SE(gen[6436]),

			.SELF(gen[6340]),
			.cell_state(gen[6340])
		); 

/******************* CELL 6341 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6341 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6245]),
			.N(gen[6246]),
			.NE(gen[6247]),

			.O(gen[6340]),
			.E(gen[6342]),

			.SO(gen[6435]),
			.S(gen[6436]),
			.SE(gen[6437]),

			.SELF(gen[6341]),
			.cell_state(gen[6341])
		); 

/******************* CELL 6342 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6342 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6246]),
			.N(gen[6247]),
			.NE(gen[6248]),

			.O(gen[6341]),
			.E(gen[6343]),

			.SO(gen[6436]),
			.S(gen[6437]),
			.SE(gen[6438]),

			.SELF(gen[6342]),
			.cell_state(gen[6342])
		); 

/******************* CELL 6343 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6343 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6247]),
			.N(gen[6248]),
			.NE(gen[6249]),

			.O(gen[6342]),
			.E(gen[6344]),

			.SO(gen[6437]),
			.S(gen[6438]),
			.SE(gen[6439]),

			.SELF(gen[6343]),
			.cell_state(gen[6343])
		); 

/******************* CELL 6344 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6344 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6248]),
			.N(gen[6249]),
			.NE(gen[6250]),

			.O(gen[6343]),
			.E(gen[6345]),

			.SO(gen[6438]),
			.S(gen[6439]),
			.SE(gen[6440]),

			.SELF(gen[6344]),
			.cell_state(gen[6344])
		); 

/******************* CELL 6345 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6345 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6249]),
			.N(gen[6250]),
			.NE(gen[6251]),

			.O(gen[6344]),
			.E(gen[6346]),

			.SO(gen[6439]),
			.S(gen[6440]),
			.SE(gen[6441]),

			.SELF(gen[6345]),
			.cell_state(gen[6345])
		); 

/******************* CELL 6346 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6346 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6250]),
			.N(gen[6251]),
			.NE(gen[6252]),

			.O(gen[6345]),
			.E(gen[6347]),

			.SO(gen[6440]),
			.S(gen[6441]),
			.SE(gen[6442]),

			.SELF(gen[6346]),
			.cell_state(gen[6346])
		); 

/******************* CELL 6347 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6347 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6251]),
			.N(gen[6252]),
			.NE(gen[6253]),

			.O(gen[6346]),
			.E(gen[6348]),

			.SO(gen[6441]),
			.S(gen[6442]),
			.SE(gen[6443]),

			.SELF(gen[6347]),
			.cell_state(gen[6347])
		); 

/******************* CELL 6348 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6348 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6252]),
			.N(gen[6253]),
			.NE(gen[6254]),

			.O(gen[6347]),
			.E(gen[6349]),

			.SO(gen[6442]),
			.S(gen[6443]),
			.SE(gen[6444]),

			.SELF(gen[6348]),
			.cell_state(gen[6348])
		); 

/******************* CELL 6349 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6349 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6253]),
			.N(gen[6254]),
			.NE(gen[6255]),

			.O(gen[6348]),
			.E(gen[6350]),

			.SO(gen[6443]),
			.S(gen[6444]),
			.SE(gen[6445]),

			.SELF(gen[6349]),
			.cell_state(gen[6349])
		); 

/******************* CELL 6350 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6350 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6254]),
			.N(gen[6255]),
			.NE(gen[6256]),

			.O(gen[6349]),
			.E(gen[6351]),

			.SO(gen[6444]),
			.S(gen[6445]),
			.SE(gen[6446]),

			.SELF(gen[6350]),
			.cell_state(gen[6350])
		); 

/******************* CELL 6351 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6351 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6255]),
			.N(gen[6256]),
			.NE(gen[6257]),

			.O(gen[6350]),
			.E(gen[6352]),

			.SO(gen[6445]),
			.S(gen[6446]),
			.SE(gen[6447]),

			.SELF(gen[6351]),
			.cell_state(gen[6351])
		); 

/******************* CELL 6352 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6352 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6256]),
			.N(gen[6257]),
			.NE(gen[6258]),

			.O(gen[6351]),
			.E(gen[6353]),

			.SO(gen[6446]),
			.S(gen[6447]),
			.SE(gen[6448]),

			.SELF(gen[6352]),
			.cell_state(gen[6352])
		); 

/******************* CELL 6353 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6353 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6257]),
			.N(gen[6258]),
			.NE(gen[6259]),

			.O(gen[6352]),
			.E(gen[6354]),

			.SO(gen[6447]),
			.S(gen[6448]),
			.SE(gen[6449]),

			.SELF(gen[6353]),
			.cell_state(gen[6353])
		); 

/******************* CELL 6354 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6354 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6258]),
			.N(gen[6259]),
			.NE(gen[6260]),

			.O(gen[6353]),
			.E(gen[6355]),

			.SO(gen[6448]),
			.S(gen[6449]),
			.SE(gen[6450]),

			.SELF(gen[6354]),
			.cell_state(gen[6354])
		); 

/******************* CELL 6355 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6355 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6259]),
			.N(gen[6260]),
			.NE(gen[6261]),

			.O(gen[6354]),
			.E(gen[6356]),

			.SO(gen[6449]),
			.S(gen[6450]),
			.SE(gen[6451]),

			.SELF(gen[6355]),
			.cell_state(gen[6355])
		); 

/******************* CELL 6356 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6356 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6260]),
			.N(gen[6261]),
			.NE(gen[6262]),

			.O(gen[6355]),
			.E(gen[6357]),

			.SO(gen[6450]),
			.S(gen[6451]),
			.SE(gen[6452]),

			.SELF(gen[6356]),
			.cell_state(gen[6356])
		); 

/******************* CELL 6357 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6357 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6261]),
			.N(gen[6262]),
			.NE(gen[6263]),

			.O(gen[6356]),
			.E(gen[6358]),

			.SO(gen[6451]),
			.S(gen[6452]),
			.SE(gen[6453]),

			.SELF(gen[6357]),
			.cell_state(gen[6357])
		); 

/******************* CELL 6358 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6358 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6262]),
			.N(gen[6263]),
			.NE(gen[6264]),

			.O(gen[6357]),
			.E(gen[6359]),

			.SO(gen[6452]),
			.S(gen[6453]),
			.SE(gen[6454]),

			.SELF(gen[6358]),
			.cell_state(gen[6358])
		); 

/******************* CELL 6359 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6359 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6263]),
			.N(gen[6264]),
			.NE(gen[6265]),

			.O(gen[6358]),
			.E(gen[6360]),

			.SO(gen[6453]),
			.S(gen[6454]),
			.SE(gen[6455]),

			.SELF(gen[6359]),
			.cell_state(gen[6359])
		); 

/******************* CELL 6360 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6360 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6264]),
			.N(gen[6265]),
			.NE(gen[6266]),

			.O(gen[6359]),
			.E(gen[6361]),

			.SO(gen[6454]),
			.S(gen[6455]),
			.SE(gen[6456]),

			.SELF(gen[6360]),
			.cell_state(gen[6360])
		); 

/******************* CELL 6361 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6361 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6265]),
			.N(gen[6266]),
			.NE(gen[6267]),

			.O(gen[6360]),
			.E(gen[6362]),

			.SO(gen[6455]),
			.S(gen[6456]),
			.SE(gen[6457]),

			.SELF(gen[6361]),
			.cell_state(gen[6361])
		); 

/******************* CELL 6362 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6362 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6266]),
			.N(gen[6267]),
			.NE(gen[6268]),

			.O(gen[6361]),
			.E(gen[6363]),

			.SO(gen[6456]),
			.S(gen[6457]),
			.SE(gen[6458]),

			.SELF(gen[6362]),
			.cell_state(gen[6362])
		); 

/******************* CELL 6363 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6363 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6267]),
			.N(gen[6268]),
			.NE(gen[6269]),

			.O(gen[6362]),
			.E(gen[6364]),

			.SO(gen[6457]),
			.S(gen[6458]),
			.SE(gen[6459]),

			.SELF(gen[6363]),
			.cell_state(gen[6363])
		); 

/******************* CELL 6364 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6364 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6268]),
			.N(gen[6269]),
			.NE(gen[6268]),

			.O(gen[6363]),
			.E(gen[6363]),

			.SO(gen[6458]),
			.S(gen[6459]),
			.SE(gen[6458]),

			.SELF(gen[6364]),
			.cell_state(gen[6364])
		); 

/******************* CELL 6365 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6365 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6271]),
			.N(gen[6270]),
			.NE(gen[6271]),

			.O(gen[6366]),
			.E(gen[6366]),

			.SO(gen[6461]),
			.S(gen[6460]),
			.SE(gen[6461]),

			.SELF(gen[6365]),
			.cell_state(gen[6365])
		); 

/******************* CELL 6366 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6366 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6270]),
			.N(gen[6271]),
			.NE(gen[6272]),

			.O(gen[6365]),
			.E(gen[6367]),

			.SO(gen[6460]),
			.S(gen[6461]),
			.SE(gen[6462]),

			.SELF(gen[6366]),
			.cell_state(gen[6366])
		); 

/******************* CELL 6367 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6367 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6271]),
			.N(gen[6272]),
			.NE(gen[6273]),

			.O(gen[6366]),
			.E(gen[6368]),

			.SO(gen[6461]),
			.S(gen[6462]),
			.SE(gen[6463]),

			.SELF(gen[6367]),
			.cell_state(gen[6367])
		); 

/******************* CELL 6368 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6368 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6272]),
			.N(gen[6273]),
			.NE(gen[6274]),

			.O(gen[6367]),
			.E(gen[6369]),

			.SO(gen[6462]),
			.S(gen[6463]),
			.SE(gen[6464]),

			.SELF(gen[6368]),
			.cell_state(gen[6368])
		); 

/******************* CELL 6369 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6369 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6273]),
			.N(gen[6274]),
			.NE(gen[6275]),

			.O(gen[6368]),
			.E(gen[6370]),

			.SO(gen[6463]),
			.S(gen[6464]),
			.SE(gen[6465]),

			.SELF(gen[6369]),
			.cell_state(gen[6369])
		); 

/******************* CELL 6370 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6370 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6274]),
			.N(gen[6275]),
			.NE(gen[6276]),

			.O(gen[6369]),
			.E(gen[6371]),

			.SO(gen[6464]),
			.S(gen[6465]),
			.SE(gen[6466]),

			.SELF(gen[6370]),
			.cell_state(gen[6370])
		); 

/******************* CELL 6371 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6371 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6275]),
			.N(gen[6276]),
			.NE(gen[6277]),

			.O(gen[6370]),
			.E(gen[6372]),

			.SO(gen[6465]),
			.S(gen[6466]),
			.SE(gen[6467]),

			.SELF(gen[6371]),
			.cell_state(gen[6371])
		); 

/******************* CELL 6372 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6372 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6276]),
			.N(gen[6277]),
			.NE(gen[6278]),

			.O(gen[6371]),
			.E(gen[6373]),

			.SO(gen[6466]),
			.S(gen[6467]),
			.SE(gen[6468]),

			.SELF(gen[6372]),
			.cell_state(gen[6372])
		); 

/******************* CELL 6373 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6373 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6277]),
			.N(gen[6278]),
			.NE(gen[6279]),

			.O(gen[6372]),
			.E(gen[6374]),

			.SO(gen[6467]),
			.S(gen[6468]),
			.SE(gen[6469]),

			.SELF(gen[6373]),
			.cell_state(gen[6373])
		); 

/******************* CELL 6374 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6374 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6278]),
			.N(gen[6279]),
			.NE(gen[6280]),

			.O(gen[6373]),
			.E(gen[6375]),

			.SO(gen[6468]),
			.S(gen[6469]),
			.SE(gen[6470]),

			.SELF(gen[6374]),
			.cell_state(gen[6374])
		); 

/******************* CELL 6375 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6375 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6279]),
			.N(gen[6280]),
			.NE(gen[6281]),

			.O(gen[6374]),
			.E(gen[6376]),

			.SO(gen[6469]),
			.S(gen[6470]),
			.SE(gen[6471]),

			.SELF(gen[6375]),
			.cell_state(gen[6375])
		); 

/******************* CELL 6376 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6376 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6280]),
			.N(gen[6281]),
			.NE(gen[6282]),

			.O(gen[6375]),
			.E(gen[6377]),

			.SO(gen[6470]),
			.S(gen[6471]),
			.SE(gen[6472]),

			.SELF(gen[6376]),
			.cell_state(gen[6376])
		); 

/******************* CELL 6377 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6377 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6281]),
			.N(gen[6282]),
			.NE(gen[6283]),

			.O(gen[6376]),
			.E(gen[6378]),

			.SO(gen[6471]),
			.S(gen[6472]),
			.SE(gen[6473]),

			.SELF(gen[6377]),
			.cell_state(gen[6377])
		); 

/******************* CELL 6378 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6378 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6282]),
			.N(gen[6283]),
			.NE(gen[6284]),

			.O(gen[6377]),
			.E(gen[6379]),

			.SO(gen[6472]),
			.S(gen[6473]),
			.SE(gen[6474]),

			.SELF(gen[6378]),
			.cell_state(gen[6378])
		); 

/******************* CELL 6379 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6379 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6283]),
			.N(gen[6284]),
			.NE(gen[6285]),

			.O(gen[6378]),
			.E(gen[6380]),

			.SO(gen[6473]),
			.S(gen[6474]),
			.SE(gen[6475]),

			.SELF(gen[6379]),
			.cell_state(gen[6379])
		); 

/******************* CELL 6380 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6380 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6284]),
			.N(gen[6285]),
			.NE(gen[6286]),

			.O(gen[6379]),
			.E(gen[6381]),

			.SO(gen[6474]),
			.S(gen[6475]),
			.SE(gen[6476]),

			.SELF(gen[6380]),
			.cell_state(gen[6380])
		); 

/******************* CELL 6381 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6381 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6285]),
			.N(gen[6286]),
			.NE(gen[6287]),

			.O(gen[6380]),
			.E(gen[6382]),

			.SO(gen[6475]),
			.S(gen[6476]),
			.SE(gen[6477]),

			.SELF(gen[6381]),
			.cell_state(gen[6381])
		); 

/******************* CELL 6382 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6382 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6286]),
			.N(gen[6287]),
			.NE(gen[6288]),

			.O(gen[6381]),
			.E(gen[6383]),

			.SO(gen[6476]),
			.S(gen[6477]),
			.SE(gen[6478]),

			.SELF(gen[6382]),
			.cell_state(gen[6382])
		); 

/******************* CELL 6383 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6383 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6287]),
			.N(gen[6288]),
			.NE(gen[6289]),

			.O(gen[6382]),
			.E(gen[6384]),

			.SO(gen[6477]),
			.S(gen[6478]),
			.SE(gen[6479]),

			.SELF(gen[6383]),
			.cell_state(gen[6383])
		); 

/******************* CELL 6384 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6384 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6288]),
			.N(gen[6289]),
			.NE(gen[6290]),

			.O(gen[6383]),
			.E(gen[6385]),

			.SO(gen[6478]),
			.S(gen[6479]),
			.SE(gen[6480]),

			.SELF(gen[6384]),
			.cell_state(gen[6384])
		); 

/******************* CELL 6385 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6385 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6289]),
			.N(gen[6290]),
			.NE(gen[6291]),

			.O(gen[6384]),
			.E(gen[6386]),

			.SO(gen[6479]),
			.S(gen[6480]),
			.SE(gen[6481]),

			.SELF(gen[6385]),
			.cell_state(gen[6385])
		); 

/******************* CELL 6386 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6386 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6290]),
			.N(gen[6291]),
			.NE(gen[6292]),

			.O(gen[6385]),
			.E(gen[6387]),

			.SO(gen[6480]),
			.S(gen[6481]),
			.SE(gen[6482]),

			.SELF(gen[6386]),
			.cell_state(gen[6386])
		); 

/******************* CELL 6387 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6387 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6291]),
			.N(gen[6292]),
			.NE(gen[6293]),

			.O(gen[6386]),
			.E(gen[6388]),

			.SO(gen[6481]),
			.S(gen[6482]),
			.SE(gen[6483]),

			.SELF(gen[6387]),
			.cell_state(gen[6387])
		); 

/******************* CELL 6388 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6388 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6292]),
			.N(gen[6293]),
			.NE(gen[6294]),

			.O(gen[6387]),
			.E(gen[6389]),

			.SO(gen[6482]),
			.S(gen[6483]),
			.SE(gen[6484]),

			.SELF(gen[6388]),
			.cell_state(gen[6388])
		); 

/******************* CELL 6389 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6389 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6293]),
			.N(gen[6294]),
			.NE(gen[6295]),

			.O(gen[6388]),
			.E(gen[6390]),

			.SO(gen[6483]),
			.S(gen[6484]),
			.SE(gen[6485]),

			.SELF(gen[6389]),
			.cell_state(gen[6389])
		); 

/******************* CELL 6390 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6390 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6294]),
			.N(gen[6295]),
			.NE(gen[6296]),

			.O(gen[6389]),
			.E(gen[6391]),

			.SO(gen[6484]),
			.S(gen[6485]),
			.SE(gen[6486]),

			.SELF(gen[6390]),
			.cell_state(gen[6390])
		); 

/******************* CELL 6391 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6391 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6295]),
			.N(gen[6296]),
			.NE(gen[6297]),

			.O(gen[6390]),
			.E(gen[6392]),

			.SO(gen[6485]),
			.S(gen[6486]),
			.SE(gen[6487]),

			.SELF(gen[6391]),
			.cell_state(gen[6391])
		); 

/******************* CELL 6392 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6392 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6296]),
			.N(gen[6297]),
			.NE(gen[6298]),

			.O(gen[6391]),
			.E(gen[6393]),

			.SO(gen[6486]),
			.S(gen[6487]),
			.SE(gen[6488]),

			.SELF(gen[6392]),
			.cell_state(gen[6392])
		); 

/******************* CELL 6393 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6393 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6297]),
			.N(gen[6298]),
			.NE(gen[6299]),

			.O(gen[6392]),
			.E(gen[6394]),

			.SO(gen[6487]),
			.S(gen[6488]),
			.SE(gen[6489]),

			.SELF(gen[6393]),
			.cell_state(gen[6393])
		); 

/******************* CELL 6394 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6394 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6298]),
			.N(gen[6299]),
			.NE(gen[6300]),

			.O(gen[6393]),
			.E(gen[6395]),

			.SO(gen[6488]),
			.S(gen[6489]),
			.SE(gen[6490]),

			.SELF(gen[6394]),
			.cell_state(gen[6394])
		); 

/******************* CELL 6395 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6395 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6299]),
			.N(gen[6300]),
			.NE(gen[6301]),

			.O(gen[6394]),
			.E(gen[6396]),

			.SO(gen[6489]),
			.S(gen[6490]),
			.SE(gen[6491]),

			.SELF(gen[6395]),
			.cell_state(gen[6395])
		); 

/******************* CELL 6396 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6396 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6300]),
			.N(gen[6301]),
			.NE(gen[6302]),

			.O(gen[6395]),
			.E(gen[6397]),

			.SO(gen[6490]),
			.S(gen[6491]),
			.SE(gen[6492]),

			.SELF(gen[6396]),
			.cell_state(gen[6396])
		); 

/******************* CELL 6397 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6397 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6301]),
			.N(gen[6302]),
			.NE(gen[6303]),

			.O(gen[6396]),
			.E(gen[6398]),

			.SO(gen[6491]),
			.S(gen[6492]),
			.SE(gen[6493]),

			.SELF(gen[6397]),
			.cell_state(gen[6397])
		); 

/******************* CELL 6398 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6398 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6302]),
			.N(gen[6303]),
			.NE(gen[6304]),

			.O(gen[6397]),
			.E(gen[6399]),

			.SO(gen[6492]),
			.S(gen[6493]),
			.SE(gen[6494]),

			.SELF(gen[6398]),
			.cell_state(gen[6398])
		); 

/******************* CELL 6399 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6399 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6303]),
			.N(gen[6304]),
			.NE(gen[6305]),

			.O(gen[6398]),
			.E(gen[6400]),

			.SO(gen[6493]),
			.S(gen[6494]),
			.SE(gen[6495]),

			.SELF(gen[6399]),
			.cell_state(gen[6399])
		); 

/******************* CELL 6400 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6400 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6304]),
			.N(gen[6305]),
			.NE(gen[6306]),

			.O(gen[6399]),
			.E(gen[6401]),

			.SO(gen[6494]),
			.S(gen[6495]),
			.SE(gen[6496]),

			.SELF(gen[6400]),
			.cell_state(gen[6400])
		); 

/******************* CELL 6401 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6401 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6305]),
			.N(gen[6306]),
			.NE(gen[6307]),

			.O(gen[6400]),
			.E(gen[6402]),

			.SO(gen[6495]),
			.S(gen[6496]),
			.SE(gen[6497]),

			.SELF(gen[6401]),
			.cell_state(gen[6401])
		); 

/******************* CELL 6402 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6402 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6306]),
			.N(gen[6307]),
			.NE(gen[6308]),

			.O(gen[6401]),
			.E(gen[6403]),

			.SO(gen[6496]),
			.S(gen[6497]),
			.SE(gen[6498]),

			.SELF(gen[6402]),
			.cell_state(gen[6402])
		); 

/******************* CELL 6403 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6403 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6307]),
			.N(gen[6308]),
			.NE(gen[6309]),

			.O(gen[6402]),
			.E(gen[6404]),

			.SO(gen[6497]),
			.S(gen[6498]),
			.SE(gen[6499]),

			.SELF(gen[6403]),
			.cell_state(gen[6403])
		); 

/******************* CELL 6404 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6404 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6308]),
			.N(gen[6309]),
			.NE(gen[6310]),

			.O(gen[6403]),
			.E(gen[6405]),

			.SO(gen[6498]),
			.S(gen[6499]),
			.SE(gen[6500]),

			.SELF(gen[6404]),
			.cell_state(gen[6404])
		); 

/******************* CELL 6405 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6405 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6309]),
			.N(gen[6310]),
			.NE(gen[6311]),

			.O(gen[6404]),
			.E(gen[6406]),

			.SO(gen[6499]),
			.S(gen[6500]),
			.SE(gen[6501]),

			.SELF(gen[6405]),
			.cell_state(gen[6405])
		); 

/******************* CELL 6406 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6406 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6310]),
			.N(gen[6311]),
			.NE(gen[6312]),

			.O(gen[6405]),
			.E(gen[6407]),

			.SO(gen[6500]),
			.S(gen[6501]),
			.SE(gen[6502]),

			.SELF(gen[6406]),
			.cell_state(gen[6406])
		); 

/******************* CELL 6407 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6407 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6311]),
			.N(gen[6312]),
			.NE(gen[6313]),

			.O(gen[6406]),
			.E(gen[6408]),

			.SO(gen[6501]),
			.S(gen[6502]),
			.SE(gen[6503]),

			.SELF(gen[6407]),
			.cell_state(gen[6407])
		); 

/******************* CELL 6408 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6408 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6312]),
			.N(gen[6313]),
			.NE(gen[6314]),

			.O(gen[6407]),
			.E(gen[6409]),

			.SO(gen[6502]),
			.S(gen[6503]),
			.SE(gen[6504]),

			.SELF(gen[6408]),
			.cell_state(gen[6408])
		); 

/******************* CELL 6409 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6409 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6313]),
			.N(gen[6314]),
			.NE(gen[6315]),

			.O(gen[6408]),
			.E(gen[6410]),

			.SO(gen[6503]),
			.S(gen[6504]),
			.SE(gen[6505]),

			.SELF(gen[6409]),
			.cell_state(gen[6409])
		); 

/******************* CELL 6410 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6410 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6314]),
			.N(gen[6315]),
			.NE(gen[6316]),

			.O(gen[6409]),
			.E(gen[6411]),

			.SO(gen[6504]),
			.S(gen[6505]),
			.SE(gen[6506]),

			.SELF(gen[6410]),
			.cell_state(gen[6410])
		); 

/******************* CELL 6411 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6411 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6315]),
			.N(gen[6316]),
			.NE(gen[6317]),

			.O(gen[6410]),
			.E(gen[6412]),

			.SO(gen[6505]),
			.S(gen[6506]),
			.SE(gen[6507]),

			.SELF(gen[6411]),
			.cell_state(gen[6411])
		); 

/******************* CELL 6412 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6412 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6316]),
			.N(gen[6317]),
			.NE(gen[6318]),

			.O(gen[6411]),
			.E(gen[6413]),

			.SO(gen[6506]),
			.S(gen[6507]),
			.SE(gen[6508]),

			.SELF(gen[6412]),
			.cell_state(gen[6412])
		); 

/******************* CELL 6413 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6413 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6317]),
			.N(gen[6318]),
			.NE(gen[6319]),

			.O(gen[6412]),
			.E(gen[6414]),

			.SO(gen[6507]),
			.S(gen[6508]),
			.SE(gen[6509]),

			.SELF(gen[6413]),
			.cell_state(gen[6413])
		); 

/******************* CELL 6414 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6414 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6318]),
			.N(gen[6319]),
			.NE(gen[6320]),

			.O(gen[6413]),
			.E(gen[6415]),

			.SO(gen[6508]),
			.S(gen[6509]),
			.SE(gen[6510]),

			.SELF(gen[6414]),
			.cell_state(gen[6414])
		); 

/******************* CELL 6415 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6415 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6319]),
			.N(gen[6320]),
			.NE(gen[6321]),

			.O(gen[6414]),
			.E(gen[6416]),

			.SO(gen[6509]),
			.S(gen[6510]),
			.SE(gen[6511]),

			.SELF(gen[6415]),
			.cell_state(gen[6415])
		); 

/******************* CELL 6416 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6416 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6320]),
			.N(gen[6321]),
			.NE(gen[6322]),

			.O(gen[6415]),
			.E(gen[6417]),

			.SO(gen[6510]),
			.S(gen[6511]),
			.SE(gen[6512]),

			.SELF(gen[6416]),
			.cell_state(gen[6416])
		); 

/******************* CELL 6417 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6417 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6321]),
			.N(gen[6322]),
			.NE(gen[6323]),

			.O(gen[6416]),
			.E(gen[6418]),

			.SO(gen[6511]),
			.S(gen[6512]),
			.SE(gen[6513]),

			.SELF(gen[6417]),
			.cell_state(gen[6417])
		); 

/******************* CELL 6418 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6418 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6322]),
			.N(gen[6323]),
			.NE(gen[6324]),

			.O(gen[6417]),
			.E(gen[6419]),

			.SO(gen[6512]),
			.S(gen[6513]),
			.SE(gen[6514]),

			.SELF(gen[6418]),
			.cell_state(gen[6418])
		); 

/******************* CELL 6419 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6419 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6323]),
			.N(gen[6324]),
			.NE(gen[6325]),

			.O(gen[6418]),
			.E(gen[6420]),

			.SO(gen[6513]),
			.S(gen[6514]),
			.SE(gen[6515]),

			.SELF(gen[6419]),
			.cell_state(gen[6419])
		); 

/******************* CELL 6420 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6420 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6324]),
			.N(gen[6325]),
			.NE(gen[6326]),

			.O(gen[6419]),
			.E(gen[6421]),

			.SO(gen[6514]),
			.S(gen[6515]),
			.SE(gen[6516]),

			.SELF(gen[6420]),
			.cell_state(gen[6420])
		); 

/******************* CELL 6421 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6421 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6325]),
			.N(gen[6326]),
			.NE(gen[6327]),

			.O(gen[6420]),
			.E(gen[6422]),

			.SO(gen[6515]),
			.S(gen[6516]),
			.SE(gen[6517]),

			.SELF(gen[6421]),
			.cell_state(gen[6421])
		); 

/******************* CELL 6422 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6422 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6326]),
			.N(gen[6327]),
			.NE(gen[6328]),

			.O(gen[6421]),
			.E(gen[6423]),

			.SO(gen[6516]),
			.S(gen[6517]),
			.SE(gen[6518]),

			.SELF(gen[6422]),
			.cell_state(gen[6422])
		); 

/******************* CELL 6423 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6423 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6327]),
			.N(gen[6328]),
			.NE(gen[6329]),

			.O(gen[6422]),
			.E(gen[6424]),

			.SO(gen[6517]),
			.S(gen[6518]),
			.SE(gen[6519]),

			.SELF(gen[6423]),
			.cell_state(gen[6423])
		); 

/******************* CELL 6424 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6424 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6328]),
			.N(gen[6329]),
			.NE(gen[6330]),

			.O(gen[6423]),
			.E(gen[6425]),

			.SO(gen[6518]),
			.S(gen[6519]),
			.SE(gen[6520]),

			.SELF(gen[6424]),
			.cell_state(gen[6424])
		); 

/******************* CELL 6425 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6425 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6329]),
			.N(gen[6330]),
			.NE(gen[6331]),

			.O(gen[6424]),
			.E(gen[6426]),

			.SO(gen[6519]),
			.S(gen[6520]),
			.SE(gen[6521]),

			.SELF(gen[6425]),
			.cell_state(gen[6425])
		); 

/******************* CELL 6426 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6426 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6330]),
			.N(gen[6331]),
			.NE(gen[6332]),

			.O(gen[6425]),
			.E(gen[6427]),

			.SO(gen[6520]),
			.S(gen[6521]),
			.SE(gen[6522]),

			.SELF(gen[6426]),
			.cell_state(gen[6426])
		); 

/******************* CELL 6427 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6427 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6331]),
			.N(gen[6332]),
			.NE(gen[6333]),

			.O(gen[6426]),
			.E(gen[6428]),

			.SO(gen[6521]),
			.S(gen[6522]),
			.SE(gen[6523]),

			.SELF(gen[6427]),
			.cell_state(gen[6427])
		); 

/******************* CELL 6428 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6428 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6332]),
			.N(gen[6333]),
			.NE(gen[6334]),

			.O(gen[6427]),
			.E(gen[6429]),

			.SO(gen[6522]),
			.S(gen[6523]),
			.SE(gen[6524]),

			.SELF(gen[6428]),
			.cell_state(gen[6428])
		); 

/******************* CELL 6429 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6429 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6333]),
			.N(gen[6334]),
			.NE(gen[6335]),

			.O(gen[6428]),
			.E(gen[6430]),

			.SO(gen[6523]),
			.S(gen[6524]),
			.SE(gen[6525]),

			.SELF(gen[6429]),
			.cell_state(gen[6429])
		); 

/******************* CELL 6430 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6430 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6334]),
			.N(gen[6335]),
			.NE(gen[6336]),

			.O(gen[6429]),
			.E(gen[6431]),

			.SO(gen[6524]),
			.S(gen[6525]),
			.SE(gen[6526]),

			.SELF(gen[6430]),
			.cell_state(gen[6430])
		); 

/******************* CELL 6431 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6431 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6335]),
			.N(gen[6336]),
			.NE(gen[6337]),

			.O(gen[6430]),
			.E(gen[6432]),

			.SO(gen[6525]),
			.S(gen[6526]),
			.SE(gen[6527]),

			.SELF(gen[6431]),
			.cell_state(gen[6431])
		); 

/******************* CELL 6432 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6432 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6336]),
			.N(gen[6337]),
			.NE(gen[6338]),

			.O(gen[6431]),
			.E(gen[6433]),

			.SO(gen[6526]),
			.S(gen[6527]),
			.SE(gen[6528]),

			.SELF(gen[6432]),
			.cell_state(gen[6432])
		); 

/******************* CELL 6433 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6433 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6337]),
			.N(gen[6338]),
			.NE(gen[6339]),

			.O(gen[6432]),
			.E(gen[6434]),

			.SO(gen[6527]),
			.S(gen[6528]),
			.SE(gen[6529]),

			.SELF(gen[6433]),
			.cell_state(gen[6433])
		); 

/******************* CELL 6434 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6434 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6338]),
			.N(gen[6339]),
			.NE(gen[6340]),

			.O(gen[6433]),
			.E(gen[6435]),

			.SO(gen[6528]),
			.S(gen[6529]),
			.SE(gen[6530]),

			.SELF(gen[6434]),
			.cell_state(gen[6434])
		); 

/******************* CELL 6435 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6435 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6339]),
			.N(gen[6340]),
			.NE(gen[6341]),

			.O(gen[6434]),
			.E(gen[6436]),

			.SO(gen[6529]),
			.S(gen[6530]),
			.SE(gen[6531]),

			.SELF(gen[6435]),
			.cell_state(gen[6435])
		); 

/******************* CELL 6436 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6436 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6340]),
			.N(gen[6341]),
			.NE(gen[6342]),

			.O(gen[6435]),
			.E(gen[6437]),

			.SO(gen[6530]),
			.S(gen[6531]),
			.SE(gen[6532]),

			.SELF(gen[6436]),
			.cell_state(gen[6436])
		); 

/******************* CELL 6437 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6437 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6341]),
			.N(gen[6342]),
			.NE(gen[6343]),

			.O(gen[6436]),
			.E(gen[6438]),

			.SO(gen[6531]),
			.S(gen[6532]),
			.SE(gen[6533]),

			.SELF(gen[6437]),
			.cell_state(gen[6437])
		); 

/******************* CELL 6438 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6438 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6342]),
			.N(gen[6343]),
			.NE(gen[6344]),

			.O(gen[6437]),
			.E(gen[6439]),

			.SO(gen[6532]),
			.S(gen[6533]),
			.SE(gen[6534]),

			.SELF(gen[6438]),
			.cell_state(gen[6438])
		); 

/******************* CELL 6439 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6439 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6343]),
			.N(gen[6344]),
			.NE(gen[6345]),

			.O(gen[6438]),
			.E(gen[6440]),

			.SO(gen[6533]),
			.S(gen[6534]),
			.SE(gen[6535]),

			.SELF(gen[6439]),
			.cell_state(gen[6439])
		); 

/******************* CELL 6440 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6440 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6344]),
			.N(gen[6345]),
			.NE(gen[6346]),

			.O(gen[6439]),
			.E(gen[6441]),

			.SO(gen[6534]),
			.S(gen[6535]),
			.SE(gen[6536]),

			.SELF(gen[6440]),
			.cell_state(gen[6440])
		); 

/******************* CELL 6441 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6441 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6345]),
			.N(gen[6346]),
			.NE(gen[6347]),

			.O(gen[6440]),
			.E(gen[6442]),

			.SO(gen[6535]),
			.S(gen[6536]),
			.SE(gen[6537]),

			.SELF(gen[6441]),
			.cell_state(gen[6441])
		); 

/******************* CELL 6442 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6442 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6346]),
			.N(gen[6347]),
			.NE(gen[6348]),

			.O(gen[6441]),
			.E(gen[6443]),

			.SO(gen[6536]),
			.S(gen[6537]),
			.SE(gen[6538]),

			.SELF(gen[6442]),
			.cell_state(gen[6442])
		); 

/******************* CELL 6443 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6443 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6347]),
			.N(gen[6348]),
			.NE(gen[6349]),

			.O(gen[6442]),
			.E(gen[6444]),

			.SO(gen[6537]),
			.S(gen[6538]),
			.SE(gen[6539]),

			.SELF(gen[6443]),
			.cell_state(gen[6443])
		); 

/******************* CELL 6444 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6444 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6348]),
			.N(gen[6349]),
			.NE(gen[6350]),

			.O(gen[6443]),
			.E(gen[6445]),

			.SO(gen[6538]),
			.S(gen[6539]),
			.SE(gen[6540]),

			.SELF(gen[6444]),
			.cell_state(gen[6444])
		); 

/******************* CELL 6445 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6445 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6349]),
			.N(gen[6350]),
			.NE(gen[6351]),

			.O(gen[6444]),
			.E(gen[6446]),

			.SO(gen[6539]),
			.S(gen[6540]),
			.SE(gen[6541]),

			.SELF(gen[6445]),
			.cell_state(gen[6445])
		); 

/******************* CELL 6446 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6446 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6350]),
			.N(gen[6351]),
			.NE(gen[6352]),

			.O(gen[6445]),
			.E(gen[6447]),

			.SO(gen[6540]),
			.S(gen[6541]),
			.SE(gen[6542]),

			.SELF(gen[6446]),
			.cell_state(gen[6446])
		); 

/******************* CELL 6447 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6447 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6351]),
			.N(gen[6352]),
			.NE(gen[6353]),

			.O(gen[6446]),
			.E(gen[6448]),

			.SO(gen[6541]),
			.S(gen[6542]),
			.SE(gen[6543]),

			.SELF(gen[6447]),
			.cell_state(gen[6447])
		); 

/******************* CELL 6448 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6448 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6352]),
			.N(gen[6353]),
			.NE(gen[6354]),

			.O(gen[6447]),
			.E(gen[6449]),

			.SO(gen[6542]),
			.S(gen[6543]),
			.SE(gen[6544]),

			.SELF(gen[6448]),
			.cell_state(gen[6448])
		); 

/******************* CELL 6449 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6449 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6353]),
			.N(gen[6354]),
			.NE(gen[6355]),

			.O(gen[6448]),
			.E(gen[6450]),

			.SO(gen[6543]),
			.S(gen[6544]),
			.SE(gen[6545]),

			.SELF(gen[6449]),
			.cell_state(gen[6449])
		); 

/******************* CELL 6450 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6450 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6354]),
			.N(gen[6355]),
			.NE(gen[6356]),

			.O(gen[6449]),
			.E(gen[6451]),

			.SO(gen[6544]),
			.S(gen[6545]),
			.SE(gen[6546]),

			.SELF(gen[6450]),
			.cell_state(gen[6450])
		); 

/******************* CELL 6451 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6451 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6355]),
			.N(gen[6356]),
			.NE(gen[6357]),

			.O(gen[6450]),
			.E(gen[6452]),

			.SO(gen[6545]),
			.S(gen[6546]),
			.SE(gen[6547]),

			.SELF(gen[6451]),
			.cell_state(gen[6451])
		); 

/******************* CELL 6452 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6452 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6356]),
			.N(gen[6357]),
			.NE(gen[6358]),

			.O(gen[6451]),
			.E(gen[6453]),

			.SO(gen[6546]),
			.S(gen[6547]),
			.SE(gen[6548]),

			.SELF(gen[6452]),
			.cell_state(gen[6452])
		); 

/******************* CELL 6453 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6453 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6357]),
			.N(gen[6358]),
			.NE(gen[6359]),

			.O(gen[6452]),
			.E(gen[6454]),

			.SO(gen[6547]),
			.S(gen[6548]),
			.SE(gen[6549]),

			.SELF(gen[6453]),
			.cell_state(gen[6453])
		); 

/******************* CELL 6454 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6454 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6358]),
			.N(gen[6359]),
			.NE(gen[6360]),

			.O(gen[6453]),
			.E(gen[6455]),

			.SO(gen[6548]),
			.S(gen[6549]),
			.SE(gen[6550]),

			.SELF(gen[6454]),
			.cell_state(gen[6454])
		); 

/******************* CELL 6455 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6455 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6359]),
			.N(gen[6360]),
			.NE(gen[6361]),

			.O(gen[6454]),
			.E(gen[6456]),

			.SO(gen[6549]),
			.S(gen[6550]),
			.SE(gen[6551]),

			.SELF(gen[6455]),
			.cell_state(gen[6455])
		); 

/******************* CELL 6456 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6456 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6360]),
			.N(gen[6361]),
			.NE(gen[6362]),

			.O(gen[6455]),
			.E(gen[6457]),

			.SO(gen[6550]),
			.S(gen[6551]),
			.SE(gen[6552]),

			.SELF(gen[6456]),
			.cell_state(gen[6456])
		); 

/******************* CELL 6457 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6457 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6361]),
			.N(gen[6362]),
			.NE(gen[6363]),

			.O(gen[6456]),
			.E(gen[6458]),

			.SO(gen[6551]),
			.S(gen[6552]),
			.SE(gen[6553]),

			.SELF(gen[6457]),
			.cell_state(gen[6457])
		); 

/******************* CELL 6458 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6458 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6362]),
			.N(gen[6363]),
			.NE(gen[6364]),

			.O(gen[6457]),
			.E(gen[6459]),

			.SO(gen[6552]),
			.S(gen[6553]),
			.SE(gen[6554]),

			.SELF(gen[6458]),
			.cell_state(gen[6458])
		); 

/******************* CELL 6459 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6459 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6363]),
			.N(gen[6364]),
			.NE(gen[6363]),

			.O(gen[6458]),
			.E(gen[6458]),

			.SO(gen[6553]),
			.S(gen[6554]),
			.SE(gen[6553]),

			.SELF(gen[6459]),
			.cell_state(gen[6459])
		); 

/******************* CELL 6460 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6460 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6366]),
			.N(gen[6365]),
			.NE(gen[6366]),

			.O(gen[6461]),
			.E(gen[6461]),

			.SO(gen[6556]),
			.S(gen[6555]),
			.SE(gen[6556]),

			.SELF(gen[6460]),
			.cell_state(gen[6460])
		); 

/******************* CELL 6461 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6461 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6365]),
			.N(gen[6366]),
			.NE(gen[6367]),

			.O(gen[6460]),
			.E(gen[6462]),

			.SO(gen[6555]),
			.S(gen[6556]),
			.SE(gen[6557]),

			.SELF(gen[6461]),
			.cell_state(gen[6461])
		); 

/******************* CELL 6462 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6462 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6366]),
			.N(gen[6367]),
			.NE(gen[6368]),

			.O(gen[6461]),
			.E(gen[6463]),

			.SO(gen[6556]),
			.S(gen[6557]),
			.SE(gen[6558]),

			.SELF(gen[6462]),
			.cell_state(gen[6462])
		); 

/******************* CELL 6463 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6463 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6367]),
			.N(gen[6368]),
			.NE(gen[6369]),

			.O(gen[6462]),
			.E(gen[6464]),

			.SO(gen[6557]),
			.S(gen[6558]),
			.SE(gen[6559]),

			.SELF(gen[6463]),
			.cell_state(gen[6463])
		); 

/******************* CELL 6464 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6464 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6368]),
			.N(gen[6369]),
			.NE(gen[6370]),

			.O(gen[6463]),
			.E(gen[6465]),

			.SO(gen[6558]),
			.S(gen[6559]),
			.SE(gen[6560]),

			.SELF(gen[6464]),
			.cell_state(gen[6464])
		); 

/******************* CELL 6465 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6465 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6369]),
			.N(gen[6370]),
			.NE(gen[6371]),

			.O(gen[6464]),
			.E(gen[6466]),

			.SO(gen[6559]),
			.S(gen[6560]),
			.SE(gen[6561]),

			.SELF(gen[6465]),
			.cell_state(gen[6465])
		); 

/******************* CELL 6466 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6466 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6370]),
			.N(gen[6371]),
			.NE(gen[6372]),

			.O(gen[6465]),
			.E(gen[6467]),

			.SO(gen[6560]),
			.S(gen[6561]),
			.SE(gen[6562]),

			.SELF(gen[6466]),
			.cell_state(gen[6466])
		); 

/******************* CELL 6467 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6467 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6371]),
			.N(gen[6372]),
			.NE(gen[6373]),

			.O(gen[6466]),
			.E(gen[6468]),

			.SO(gen[6561]),
			.S(gen[6562]),
			.SE(gen[6563]),

			.SELF(gen[6467]),
			.cell_state(gen[6467])
		); 

/******************* CELL 6468 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6468 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6372]),
			.N(gen[6373]),
			.NE(gen[6374]),

			.O(gen[6467]),
			.E(gen[6469]),

			.SO(gen[6562]),
			.S(gen[6563]),
			.SE(gen[6564]),

			.SELF(gen[6468]),
			.cell_state(gen[6468])
		); 

/******************* CELL 6469 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6469 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6373]),
			.N(gen[6374]),
			.NE(gen[6375]),

			.O(gen[6468]),
			.E(gen[6470]),

			.SO(gen[6563]),
			.S(gen[6564]),
			.SE(gen[6565]),

			.SELF(gen[6469]),
			.cell_state(gen[6469])
		); 

/******************* CELL 6470 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6470 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6374]),
			.N(gen[6375]),
			.NE(gen[6376]),

			.O(gen[6469]),
			.E(gen[6471]),

			.SO(gen[6564]),
			.S(gen[6565]),
			.SE(gen[6566]),

			.SELF(gen[6470]),
			.cell_state(gen[6470])
		); 

/******************* CELL 6471 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6471 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6375]),
			.N(gen[6376]),
			.NE(gen[6377]),

			.O(gen[6470]),
			.E(gen[6472]),

			.SO(gen[6565]),
			.S(gen[6566]),
			.SE(gen[6567]),

			.SELF(gen[6471]),
			.cell_state(gen[6471])
		); 

/******************* CELL 6472 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6472 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6376]),
			.N(gen[6377]),
			.NE(gen[6378]),

			.O(gen[6471]),
			.E(gen[6473]),

			.SO(gen[6566]),
			.S(gen[6567]),
			.SE(gen[6568]),

			.SELF(gen[6472]),
			.cell_state(gen[6472])
		); 

/******************* CELL 6473 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6473 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6377]),
			.N(gen[6378]),
			.NE(gen[6379]),

			.O(gen[6472]),
			.E(gen[6474]),

			.SO(gen[6567]),
			.S(gen[6568]),
			.SE(gen[6569]),

			.SELF(gen[6473]),
			.cell_state(gen[6473])
		); 

/******************* CELL 6474 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6474 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6378]),
			.N(gen[6379]),
			.NE(gen[6380]),

			.O(gen[6473]),
			.E(gen[6475]),

			.SO(gen[6568]),
			.S(gen[6569]),
			.SE(gen[6570]),

			.SELF(gen[6474]),
			.cell_state(gen[6474])
		); 

/******************* CELL 6475 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6475 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6379]),
			.N(gen[6380]),
			.NE(gen[6381]),

			.O(gen[6474]),
			.E(gen[6476]),

			.SO(gen[6569]),
			.S(gen[6570]),
			.SE(gen[6571]),

			.SELF(gen[6475]),
			.cell_state(gen[6475])
		); 

/******************* CELL 6476 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6476 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6380]),
			.N(gen[6381]),
			.NE(gen[6382]),

			.O(gen[6475]),
			.E(gen[6477]),

			.SO(gen[6570]),
			.S(gen[6571]),
			.SE(gen[6572]),

			.SELF(gen[6476]),
			.cell_state(gen[6476])
		); 

/******************* CELL 6477 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6477 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6381]),
			.N(gen[6382]),
			.NE(gen[6383]),

			.O(gen[6476]),
			.E(gen[6478]),

			.SO(gen[6571]),
			.S(gen[6572]),
			.SE(gen[6573]),

			.SELF(gen[6477]),
			.cell_state(gen[6477])
		); 

/******************* CELL 6478 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6478 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6382]),
			.N(gen[6383]),
			.NE(gen[6384]),

			.O(gen[6477]),
			.E(gen[6479]),

			.SO(gen[6572]),
			.S(gen[6573]),
			.SE(gen[6574]),

			.SELF(gen[6478]),
			.cell_state(gen[6478])
		); 

/******************* CELL 6479 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6479 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6383]),
			.N(gen[6384]),
			.NE(gen[6385]),

			.O(gen[6478]),
			.E(gen[6480]),

			.SO(gen[6573]),
			.S(gen[6574]),
			.SE(gen[6575]),

			.SELF(gen[6479]),
			.cell_state(gen[6479])
		); 

/******************* CELL 6480 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6480 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6384]),
			.N(gen[6385]),
			.NE(gen[6386]),

			.O(gen[6479]),
			.E(gen[6481]),

			.SO(gen[6574]),
			.S(gen[6575]),
			.SE(gen[6576]),

			.SELF(gen[6480]),
			.cell_state(gen[6480])
		); 

/******************* CELL 6481 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6481 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6385]),
			.N(gen[6386]),
			.NE(gen[6387]),

			.O(gen[6480]),
			.E(gen[6482]),

			.SO(gen[6575]),
			.S(gen[6576]),
			.SE(gen[6577]),

			.SELF(gen[6481]),
			.cell_state(gen[6481])
		); 

/******************* CELL 6482 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6482 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6386]),
			.N(gen[6387]),
			.NE(gen[6388]),

			.O(gen[6481]),
			.E(gen[6483]),

			.SO(gen[6576]),
			.S(gen[6577]),
			.SE(gen[6578]),

			.SELF(gen[6482]),
			.cell_state(gen[6482])
		); 

/******************* CELL 6483 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6483 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6387]),
			.N(gen[6388]),
			.NE(gen[6389]),

			.O(gen[6482]),
			.E(gen[6484]),

			.SO(gen[6577]),
			.S(gen[6578]),
			.SE(gen[6579]),

			.SELF(gen[6483]),
			.cell_state(gen[6483])
		); 

/******************* CELL 6484 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6484 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6388]),
			.N(gen[6389]),
			.NE(gen[6390]),

			.O(gen[6483]),
			.E(gen[6485]),

			.SO(gen[6578]),
			.S(gen[6579]),
			.SE(gen[6580]),

			.SELF(gen[6484]),
			.cell_state(gen[6484])
		); 

/******************* CELL 6485 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6485 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6389]),
			.N(gen[6390]),
			.NE(gen[6391]),

			.O(gen[6484]),
			.E(gen[6486]),

			.SO(gen[6579]),
			.S(gen[6580]),
			.SE(gen[6581]),

			.SELF(gen[6485]),
			.cell_state(gen[6485])
		); 

/******************* CELL 6486 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6486 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6390]),
			.N(gen[6391]),
			.NE(gen[6392]),

			.O(gen[6485]),
			.E(gen[6487]),

			.SO(gen[6580]),
			.S(gen[6581]),
			.SE(gen[6582]),

			.SELF(gen[6486]),
			.cell_state(gen[6486])
		); 

/******************* CELL 6487 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6487 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6391]),
			.N(gen[6392]),
			.NE(gen[6393]),

			.O(gen[6486]),
			.E(gen[6488]),

			.SO(gen[6581]),
			.S(gen[6582]),
			.SE(gen[6583]),

			.SELF(gen[6487]),
			.cell_state(gen[6487])
		); 

/******************* CELL 6488 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6488 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6392]),
			.N(gen[6393]),
			.NE(gen[6394]),

			.O(gen[6487]),
			.E(gen[6489]),

			.SO(gen[6582]),
			.S(gen[6583]),
			.SE(gen[6584]),

			.SELF(gen[6488]),
			.cell_state(gen[6488])
		); 

/******************* CELL 6489 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6489 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6393]),
			.N(gen[6394]),
			.NE(gen[6395]),

			.O(gen[6488]),
			.E(gen[6490]),

			.SO(gen[6583]),
			.S(gen[6584]),
			.SE(gen[6585]),

			.SELF(gen[6489]),
			.cell_state(gen[6489])
		); 

/******************* CELL 6490 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6490 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6394]),
			.N(gen[6395]),
			.NE(gen[6396]),

			.O(gen[6489]),
			.E(gen[6491]),

			.SO(gen[6584]),
			.S(gen[6585]),
			.SE(gen[6586]),

			.SELF(gen[6490]),
			.cell_state(gen[6490])
		); 

/******************* CELL 6491 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6491 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6395]),
			.N(gen[6396]),
			.NE(gen[6397]),

			.O(gen[6490]),
			.E(gen[6492]),

			.SO(gen[6585]),
			.S(gen[6586]),
			.SE(gen[6587]),

			.SELF(gen[6491]),
			.cell_state(gen[6491])
		); 

/******************* CELL 6492 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6492 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6396]),
			.N(gen[6397]),
			.NE(gen[6398]),

			.O(gen[6491]),
			.E(gen[6493]),

			.SO(gen[6586]),
			.S(gen[6587]),
			.SE(gen[6588]),

			.SELF(gen[6492]),
			.cell_state(gen[6492])
		); 

/******************* CELL 6493 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6493 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6397]),
			.N(gen[6398]),
			.NE(gen[6399]),

			.O(gen[6492]),
			.E(gen[6494]),

			.SO(gen[6587]),
			.S(gen[6588]),
			.SE(gen[6589]),

			.SELF(gen[6493]),
			.cell_state(gen[6493])
		); 

/******************* CELL 6494 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6494 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6398]),
			.N(gen[6399]),
			.NE(gen[6400]),

			.O(gen[6493]),
			.E(gen[6495]),

			.SO(gen[6588]),
			.S(gen[6589]),
			.SE(gen[6590]),

			.SELF(gen[6494]),
			.cell_state(gen[6494])
		); 

/******************* CELL 6495 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6495 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6399]),
			.N(gen[6400]),
			.NE(gen[6401]),

			.O(gen[6494]),
			.E(gen[6496]),

			.SO(gen[6589]),
			.S(gen[6590]),
			.SE(gen[6591]),

			.SELF(gen[6495]),
			.cell_state(gen[6495])
		); 

/******************* CELL 6496 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6496 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6400]),
			.N(gen[6401]),
			.NE(gen[6402]),

			.O(gen[6495]),
			.E(gen[6497]),

			.SO(gen[6590]),
			.S(gen[6591]),
			.SE(gen[6592]),

			.SELF(gen[6496]),
			.cell_state(gen[6496])
		); 

/******************* CELL 6497 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6497 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6401]),
			.N(gen[6402]),
			.NE(gen[6403]),

			.O(gen[6496]),
			.E(gen[6498]),

			.SO(gen[6591]),
			.S(gen[6592]),
			.SE(gen[6593]),

			.SELF(gen[6497]),
			.cell_state(gen[6497])
		); 

/******************* CELL 6498 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6498 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6402]),
			.N(gen[6403]),
			.NE(gen[6404]),

			.O(gen[6497]),
			.E(gen[6499]),

			.SO(gen[6592]),
			.S(gen[6593]),
			.SE(gen[6594]),

			.SELF(gen[6498]),
			.cell_state(gen[6498])
		); 

/******************* CELL 6499 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6499 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6403]),
			.N(gen[6404]),
			.NE(gen[6405]),

			.O(gen[6498]),
			.E(gen[6500]),

			.SO(gen[6593]),
			.S(gen[6594]),
			.SE(gen[6595]),

			.SELF(gen[6499]),
			.cell_state(gen[6499])
		); 

/******************* CELL 6500 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6500 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6404]),
			.N(gen[6405]),
			.NE(gen[6406]),

			.O(gen[6499]),
			.E(gen[6501]),

			.SO(gen[6594]),
			.S(gen[6595]),
			.SE(gen[6596]),

			.SELF(gen[6500]),
			.cell_state(gen[6500])
		); 

/******************* CELL 6501 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6501 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6405]),
			.N(gen[6406]),
			.NE(gen[6407]),

			.O(gen[6500]),
			.E(gen[6502]),

			.SO(gen[6595]),
			.S(gen[6596]),
			.SE(gen[6597]),

			.SELF(gen[6501]),
			.cell_state(gen[6501])
		); 

/******************* CELL 6502 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6502 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6406]),
			.N(gen[6407]),
			.NE(gen[6408]),

			.O(gen[6501]),
			.E(gen[6503]),

			.SO(gen[6596]),
			.S(gen[6597]),
			.SE(gen[6598]),

			.SELF(gen[6502]),
			.cell_state(gen[6502])
		); 

/******************* CELL 6503 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6503 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6407]),
			.N(gen[6408]),
			.NE(gen[6409]),

			.O(gen[6502]),
			.E(gen[6504]),

			.SO(gen[6597]),
			.S(gen[6598]),
			.SE(gen[6599]),

			.SELF(gen[6503]),
			.cell_state(gen[6503])
		); 

/******************* CELL 6504 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6504 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6408]),
			.N(gen[6409]),
			.NE(gen[6410]),

			.O(gen[6503]),
			.E(gen[6505]),

			.SO(gen[6598]),
			.S(gen[6599]),
			.SE(gen[6600]),

			.SELF(gen[6504]),
			.cell_state(gen[6504])
		); 

/******************* CELL 6505 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6505 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6409]),
			.N(gen[6410]),
			.NE(gen[6411]),

			.O(gen[6504]),
			.E(gen[6506]),

			.SO(gen[6599]),
			.S(gen[6600]),
			.SE(gen[6601]),

			.SELF(gen[6505]),
			.cell_state(gen[6505])
		); 

/******************* CELL 6506 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6506 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6410]),
			.N(gen[6411]),
			.NE(gen[6412]),

			.O(gen[6505]),
			.E(gen[6507]),

			.SO(gen[6600]),
			.S(gen[6601]),
			.SE(gen[6602]),

			.SELF(gen[6506]),
			.cell_state(gen[6506])
		); 

/******************* CELL 6507 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6507 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6411]),
			.N(gen[6412]),
			.NE(gen[6413]),

			.O(gen[6506]),
			.E(gen[6508]),

			.SO(gen[6601]),
			.S(gen[6602]),
			.SE(gen[6603]),

			.SELF(gen[6507]),
			.cell_state(gen[6507])
		); 

/******************* CELL 6508 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6508 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6412]),
			.N(gen[6413]),
			.NE(gen[6414]),

			.O(gen[6507]),
			.E(gen[6509]),

			.SO(gen[6602]),
			.S(gen[6603]),
			.SE(gen[6604]),

			.SELF(gen[6508]),
			.cell_state(gen[6508])
		); 

/******************* CELL 6509 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6509 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6413]),
			.N(gen[6414]),
			.NE(gen[6415]),

			.O(gen[6508]),
			.E(gen[6510]),

			.SO(gen[6603]),
			.S(gen[6604]),
			.SE(gen[6605]),

			.SELF(gen[6509]),
			.cell_state(gen[6509])
		); 

/******************* CELL 6510 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6510 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6414]),
			.N(gen[6415]),
			.NE(gen[6416]),

			.O(gen[6509]),
			.E(gen[6511]),

			.SO(gen[6604]),
			.S(gen[6605]),
			.SE(gen[6606]),

			.SELF(gen[6510]),
			.cell_state(gen[6510])
		); 

/******************* CELL 6511 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6511 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6415]),
			.N(gen[6416]),
			.NE(gen[6417]),

			.O(gen[6510]),
			.E(gen[6512]),

			.SO(gen[6605]),
			.S(gen[6606]),
			.SE(gen[6607]),

			.SELF(gen[6511]),
			.cell_state(gen[6511])
		); 

/******************* CELL 6512 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6512 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6416]),
			.N(gen[6417]),
			.NE(gen[6418]),

			.O(gen[6511]),
			.E(gen[6513]),

			.SO(gen[6606]),
			.S(gen[6607]),
			.SE(gen[6608]),

			.SELF(gen[6512]),
			.cell_state(gen[6512])
		); 

/******************* CELL 6513 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6513 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6417]),
			.N(gen[6418]),
			.NE(gen[6419]),

			.O(gen[6512]),
			.E(gen[6514]),

			.SO(gen[6607]),
			.S(gen[6608]),
			.SE(gen[6609]),

			.SELF(gen[6513]),
			.cell_state(gen[6513])
		); 

/******************* CELL 6514 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6514 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6418]),
			.N(gen[6419]),
			.NE(gen[6420]),

			.O(gen[6513]),
			.E(gen[6515]),

			.SO(gen[6608]),
			.S(gen[6609]),
			.SE(gen[6610]),

			.SELF(gen[6514]),
			.cell_state(gen[6514])
		); 

/******************* CELL 6515 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6515 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6419]),
			.N(gen[6420]),
			.NE(gen[6421]),

			.O(gen[6514]),
			.E(gen[6516]),

			.SO(gen[6609]),
			.S(gen[6610]),
			.SE(gen[6611]),

			.SELF(gen[6515]),
			.cell_state(gen[6515])
		); 

/******************* CELL 6516 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6516 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6420]),
			.N(gen[6421]),
			.NE(gen[6422]),

			.O(gen[6515]),
			.E(gen[6517]),

			.SO(gen[6610]),
			.S(gen[6611]),
			.SE(gen[6612]),

			.SELF(gen[6516]),
			.cell_state(gen[6516])
		); 

/******************* CELL 6517 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6517 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6421]),
			.N(gen[6422]),
			.NE(gen[6423]),

			.O(gen[6516]),
			.E(gen[6518]),

			.SO(gen[6611]),
			.S(gen[6612]),
			.SE(gen[6613]),

			.SELF(gen[6517]),
			.cell_state(gen[6517])
		); 

/******************* CELL 6518 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6518 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6422]),
			.N(gen[6423]),
			.NE(gen[6424]),

			.O(gen[6517]),
			.E(gen[6519]),

			.SO(gen[6612]),
			.S(gen[6613]),
			.SE(gen[6614]),

			.SELF(gen[6518]),
			.cell_state(gen[6518])
		); 

/******************* CELL 6519 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6519 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6423]),
			.N(gen[6424]),
			.NE(gen[6425]),

			.O(gen[6518]),
			.E(gen[6520]),

			.SO(gen[6613]),
			.S(gen[6614]),
			.SE(gen[6615]),

			.SELF(gen[6519]),
			.cell_state(gen[6519])
		); 

/******************* CELL 6520 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6520 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6424]),
			.N(gen[6425]),
			.NE(gen[6426]),

			.O(gen[6519]),
			.E(gen[6521]),

			.SO(gen[6614]),
			.S(gen[6615]),
			.SE(gen[6616]),

			.SELF(gen[6520]),
			.cell_state(gen[6520])
		); 

/******************* CELL 6521 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6521 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6425]),
			.N(gen[6426]),
			.NE(gen[6427]),

			.O(gen[6520]),
			.E(gen[6522]),

			.SO(gen[6615]),
			.S(gen[6616]),
			.SE(gen[6617]),

			.SELF(gen[6521]),
			.cell_state(gen[6521])
		); 

/******************* CELL 6522 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6522 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6426]),
			.N(gen[6427]),
			.NE(gen[6428]),

			.O(gen[6521]),
			.E(gen[6523]),

			.SO(gen[6616]),
			.S(gen[6617]),
			.SE(gen[6618]),

			.SELF(gen[6522]),
			.cell_state(gen[6522])
		); 

/******************* CELL 6523 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6523 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6427]),
			.N(gen[6428]),
			.NE(gen[6429]),

			.O(gen[6522]),
			.E(gen[6524]),

			.SO(gen[6617]),
			.S(gen[6618]),
			.SE(gen[6619]),

			.SELF(gen[6523]),
			.cell_state(gen[6523])
		); 

/******************* CELL 6524 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6524 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6428]),
			.N(gen[6429]),
			.NE(gen[6430]),

			.O(gen[6523]),
			.E(gen[6525]),

			.SO(gen[6618]),
			.S(gen[6619]),
			.SE(gen[6620]),

			.SELF(gen[6524]),
			.cell_state(gen[6524])
		); 

/******************* CELL 6525 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6525 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6429]),
			.N(gen[6430]),
			.NE(gen[6431]),

			.O(gen[6524]),
			.E(gen[6526]),

			.SO(gen[6619]),
			.S(gen[6620]),
			.SE(gen[6621]),

			.SELF(gen[6525]),
			.cell_state(gen[6525])
		); 

/******************* CELL 6526 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6526 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6430]),
			.N(gen[6431]),
			.NE(gen[6432]),

			.O(gen[6525]),
			.E(gen[6527]),

			.SO(gen[6620]),
			.S(gen[6621]),
			.SE(gen[6622]),

			.SELF(gen[6526]),
			.cell_state(gen[6526])
		); 

/******************* CELL 6527 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6527 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6431]),
			.N(gen[6432]),
			.NE(gen[6433]),

			.O(gen[6526]),
			.E(gen[6528]),

			.SO(gen[6621]),
			.S(gen[6622]),
			.SE(gen[6623]),

			.SELF(gen[6527]),
			.cell_state(gen[6527])
		); 

/******************* CELL 6528 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6528 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6432]),
			.N(gen[6433]),
			.NE(gen[6434]),

			.O(gen[6527]),
			.E(gen[6529]),

			.SO(gen[6622]),
			.S(gen[6623]),
			.SE(gen[6624]),

			.SELF(gen[6528]),
			.cell_state(gen[6528])
		); 

/******************* CELL 6529 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6529 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6433]),
			.N(gen[6434]),
			.NE(gen[6435]),

			.O(gen[6528]),
			.E(gen[6530]),

			.SO(gen[6623]),
			.S(gen[6624]),
			.SE(gen[6625]),

			.SELF(gen[6529]),
			.cell_state(gen[6529])
		); 

/******************* CELL 6530 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6530 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6434]),
			.N(gen[6435]),
			.NE(gen[6436]),

			.O(gen[6529]),
			.E(gen[6531]),

			.SO(gen[6624]),
			.S(gen[6625]),
			.SE(gen[6626]),

			.SELF(gen[6530]),
			.cell_state(gen[6530])
		); 

/******************* CELL 6531 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6531 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6435]),
			.N(gen[6436]),
			.NE(gen[6437]),

			.O(gen[6530]),
			.E(gen[6532]),

			.SO(gen[6625]),
			.S(gen[6626]),
			.SE(gen[6627]),

			.SELF(gen[6531]),
			.cell_state(gen[6531])
		); 

/******************* CELL 6532 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6532 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6436]),
			.N(gen[6437]),
			.NE(gen[6438]),

			.O(gen[6531]),
			.E(gen[6533]),

			.SO(gen[6626]),
			.S(gen[6627]),
			.SE(gen[6628]),

			.SELF(gen[6532]),
			.cell_state(gen[6532])
		); 

/******************* CELL 6533 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6533 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6437]),
			.N(gen[6438]),
			.NE(gen[6439]),

			.O(gen[6532]),
			.E(gen[6534]),

			.SO(gen[6627]),
			.S(gen[6628]),
			.SE(gen[6629]),

			.SELF(gen[6533]),
			.cell_state(gen[6533])
		); 

/******************* CELL 6534 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6534 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6438]),
			.N(gen[6439]),
			.NE(gen[6440]),

			.O(gen[6533]),
			.E(gen[6535]),

			.SO(gen[6628]),
			.S(gen[6629]),
			.SE(gen[6630]),

			.SELF(gen[6534]),
			.cell_state(gen[6534])
		); 

/******************* CELL 6535 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6535 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6439]),
			.N(gen[6440]),
			.NE(gen[6441]),

			.O(gen[6534]),
			.E(gen[6536]),

			.SO(gen[6629]),
			.S(gen[6630]),
			.SE(gen[6631]),

			.SELF(gen[6535]),
			.cell_state(gen[6535])
		); 

/******************* CELL 6536 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6536 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6440]),
			.N(gen[6441]),
			.NE(gen[6442]),

			.O(gen[6535]),
			.E(gen[6537]),

			.SO(gen[6630]),
			.S(gen[6631]),
			.SE(gen[6632]),

			.SELF(gen[6536]),
			.cell_state(gen[6536])
		); 

/******************* CELL 6537 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6537 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6441]),
			.N(gen[6442]),
			.NE(gen[6443]),

			.O(gen[6536]),
			.E(gen[6538]),

			.SO(gen[6631]),
			.S(gen[6632]),
			.SE(gen[6633]),

			.SELF(gen[6537]),
			.cell_state(gen[6537])
		); 

/******************* CELL 6538 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6538 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6442]),
			.N(gen[6443]),
			.NE(gen[6444]),

			.O(gen[6537]),
			.E(gen[6539]),

			.SO(gen[6632]),
			.S(gen[6633]),
			.SE(gen[6634]),

			.SELF(gen[6538]),
			.cell_state(gen[6538])
		); 

/******************* CELL 6539 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6539 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6443]),
			.N(gen[6444]),
			.NE(gen[6445]),

			.O(gen[6538]),
			.E(gen[6540]),

			.SO(gen[6633]),
			.S(gen[6634]),
			.SE(gen[6635]),

			.SELF(gen[6539]),
			.cell_state(gen[6539])
		); 

/******************* CELL 6540 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6540 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6444]),
			.N(gen[6445]),
			.NE(gen[6446]),

			.O(gen[6539]),
			.E(gen[6541]),

			.SO(gen[6634]),
			.S(gen[6635]),
			.SE(gen[6636]),

			.SELF(gen[6540]),
			.cell_state(gen[6540])
		); 

/******************* CELL 6541 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6541 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6445]),
			.N(gen[6446]),
			.NE(gen[6447]),

			.O(gen[6540]),
			.E(gen[6542]),

			.SO(gen[6635]),
			.S(gen[6636]),
			.SE(gen[6637]),

			.SELF(gen[6541]),
			.cell_state(gen[6541])
		); 

/******************* CELL 6542 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6542 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6446]),
			.N(gen[6447]),
			.NE(gen[6448]),

			.O(gen[6541]),
			.E(gen[6543]),

			.SO(gen[6636]),
			.S(gen[6637]),
			.SE(gen[6638]),

			.SELF(gen[6542]),
			.cell_state(gen[6542])
		); 

/******************* CELL 6543 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6543 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6447]),
			.N(gen[6448]),
			.NE(gen[6449]),

			.O(gen[6542]),
			.E(gen[6544]),

			.SO(gen[6637]),
			.S(gen[6638]),
			.SE(gen[6639]),

			.SELF(gen[6543]),
			.cell_state(gen[6543])
		); 

/******************* CELL 6544 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6544 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6448]),
			.N(gen[6449]),
			.NE(gen[6450]),

			.O(gen[6543]),
			.E(gen[6545]),

			.SO(gen[6638]),
			.S(gen[6639]),
			.SE(gen[6640]),

			.SELF(gen[6544]),
			.cell_state(gen[6544])
		); 

/******************* CELL 6545 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6545 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6449]),
			.N(gen[6450]),
			.NE(gen[6451]),

			.O(gen[6544]),
			.E(gen[6546]),

			.SO(gen[6639]),
			.S(gen[6640]),
			.SE(gen[6641]),

			.SELF(gen[6545]),
			.cell_state(gen[6545])
		); 

/******************* CELL 6546 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6546 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6450]),
			.N(gen[6451]),
			.NE(gen[6452]),

			.O(gen[6545]),
			.E(gen[6547]),

			.SO(gen[6640]),
			.S(gen[6641]),
			.SE(gen[6642]),

			.SELF(gen[6546]),
			.cell_state(gen[6546])
		); 

/******************* CELL 6547 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6547 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6451]),
			.N(gen[6452]),
			.NE(gen[6453]),

			.O(gen[6546]),
			.E(gen[6548]),

			.SO(gen[6641]),
			.S(gen[6642]),
			.SE(gen[6643]),

			.SELF(gen[6547]),
			.cell_state(gen[6547])
		); 

/******************* CELL 6548 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6548 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6452]),
			.N(gen[6453]),
			.NE(gen[6454]),

			.O(gen[6547]),
			.E(gen[6549]),

			.SO(gen[6642]),
			.S(gen[6643]),
			.SE(gen[6644]),

			.SELF(gen[6548]),
			.cell_state(gen[6548])
		); 

/******************* CELL 6549 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6549 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6453]),
			.N(gen[6454]),
			.NE(gen[6455]),

			.O(gen[6548]),
			.E(gen[6550]),

			.SO(gen[6643]),
			.S(gen[6644]),
			.SE(gen[6645]),

			.SELF(gen[6549]),
			.cell_state(gen[6549])
		); 

/******************* CELL 6550 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6550 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6454]),
			.N(gen[6455]),
			.NE(gen[6456]),

			.O(gen[6549]),
			.E(gen[6551]),

			.SO(gen[6644]),
			.S(gen[6645]),
			.SE(gen[6646]),

			.SELF(gen[6550]),
			.cell_state(gen[6550])
		); 

/******************* CELL 6551 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6551 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6455]),
			.N(gen[6456]),
			.NE(gen[6457]),

			.O(gen[6550]),
			.E(gen[6552]),

			.SO(gen[6645]),
			.S(gen[6646]),
			.SE(gen[6647]),

			.SELF(gen[6551]),
			.cell_state(gen[6551])
		); 

/******************* CELL 6552 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6552 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6456]),
			.N(gen[6457]),
			.NE(gen[6458]),

			.O(gen[6551]),
			.E(gen[6553]),

			.SO(gen[6646]),
			.S(gen[6647]),
			.SE(gen[6648]),

			.SELF(gen[6552]),
			.cell_state(gen[6552])
		); 

/******************* CELL 6553 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6553 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6457]),
			.N(gen[6458]),
			.NE(gen[6459]),

			.O(gen[6552]),
			.E(gen[6554]),

			.SO(gen[6647]),
			.S(gen[6648]),
			.SE(gen[6649]),

			.SELF(gen[6553]),
			.cell_state(gen[6553])
		); 

/******************* CELL 6554 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6554 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6458]),
			.N(gen[6459]),
			.NE(gen[6458]),

			.O(gen[6553]),
			.E(gen[6553]),

			.SO(gen[6648]),
			.S(gen[6649]),
			.SE(gen[6648]),

			.SELF(gen[6554]),
			.cell_state(gen[6554])
		); 

/******************* CELL 6555 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6555 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6461]),
			.N(gen[6460]),
			.NE(gen[6461]),

			.O(gen[6556]),
			.E(gen[6556]),

			.SO(gen[6651]),
			.S(gen[6650]),
			.SE(gen[6651]),

			.SELF(gen[6555]),
			.cell_state(gen[6555])
		); 

/******************* CELL 6556 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6556 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6460]),
			.N(gen[6461]),
			.NE(gen[6462]),

			.O(gen[6555]),
			.E(gen[6557]),

			.SO(gen[6650]),
			.S(gen[6651]),
			.SE(gen[6652]),

			.SELF(gen[6556]),
			.cell_state(gen[6556])
		); 

/******************* CELL 6557 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6557 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6461]),
			.N(gen[6462]),
			.NE(gen[6463]),

			.O(gen[6556]),
			.E(gen[6558]),

			.SO(gen[6651]),
			.S(gen[6652]),
			.SE(gen[6653]),

			.SELF(gen[6557]),
			.cell_state(gen[6557])
		); 

/******************* CELL 6558 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6558 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6462]),
			.N(gen[6463]),
			.NE(gen[6464]),

			.O(gen[6557]),
			.E(gen[6559]),

			.SO(gen[6652]),
			.S(gen[6653]),
			.SE(gen[6654]),

			.SELF(gen[6558]),
			.cell_state(gen[6558])
		); 

/******************* CELL 6559 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6559 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6463]),
			.N(gen[6464]),
			.NE(gen[6465]),

			.O(gen[6558]),
			.E(gen[6560]),

			.SO(gen[6653]),
			.S(gen[6654]),
			.SE(gen[6655]),

			.SELF(gen[6559]),
			.cell_state(gen[6559])
		); 

/******************* CELL 6560 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6560 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6464]),
			.N(gen[6465]),
			.NE(gen[6466]),

			.O(gen[6559]),
			.E(gen[6561]),

			.SO(gen[6654]),
			.S(gen[6655]),
			.SE(gen[6656]),

			.SELF(gen[6560]),
			.cell_state(gen[6560])
		); 

/******************* CELL 6561 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6561 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6465]),
			.N(gen[6466]),
			.NE(gen[6467]),

			.O(gen[6560]),
			.E(gen[6562]),

			.SO(gen[6655]),
			.S(gen[6656]),
			.SE(gen[6657]),

			.SELF(gen[6561]),
			.cell_state(gen[6561])
		); 

/******************* CELL 6562 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6562 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6466]),
			.N(gen[6467]),
			.NE(gen[6468]),

			.O(gen[6561]),
			.E(gen[6563]),

			.SO(gen[6656]),
			.S(gen[6657]),
			.SE(gen[6658]),

			.SELF(gen[6562]),
			.cell_state(gen[6562])
		); 

/******************* CELL 6563 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6563 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6467]),
			.N(gen[6468]),
			.NE(gen[6469]),

			.O(gen[6562]),
			.E(gen[6564]),

			.SO(gen[6657]),
			.S(gen[6658]),
			.SE(gen[6659]),

			.SELF(gen[6563]),
			.cell_state(gen[6563])
		); 

/******************* CELL 6564 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6564 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6468]),
			.N(gen[6469]),
			.NE(gen[6470]),

			.O(gen[6563]),
			.E(gen[6565]),

			.SO(gen[6658]),
			.S(gen[6659]),
			.SE(gen[6660]),

			.SELF(gen[6564]),
			.cell_state(gen[6564])
		); 

/******************* CELL 6565 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6565 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6469]),
			.N(gen[6470]),
			.NE(gen[6471]),

			.O(gen[6564]),
			.E(gen[6566]),

			.SO(gen[6659]),
			.S(gen[6660]),
			.SE(gen[6661]),

			.SELF(gen[6565]),
			.cell_state(gen[6565])
		); 

/******************* CELL 6566 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6566 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6470]),
			.N(gen[6471]),
			.NE(gen[6472]),

			.O(gen[6565]),
			.E(gen[6567]),

			.SO(gen[6660]),
			.S(gen[6661]),
			.SE(gen[6662]),

			.SELF(gen[6566]),
			.cell_state(gen[6566])
		); 

/******************* CELL 6567 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6567 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6471]),
			.N(gen[6472]),
			.NE(gen[6473]),

			.O(gen[6566]),
			.E(gen[6568]),

			.SO(gen[6661]),
			.S(gen[6662]),
			.SE(gen[6663]),

			.SELF(gen[6567]),
			.cell_state(gen[6567])
		); 

/******************* CELL 6568 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6568 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6472]),
			.N(gen[6473]),
			.NE(gen[6474]),

			.O(gen[6567]),
			.E(gen[6569]),

			.SO(gen[6662]),
			.S(gen[6663]),
			.SE(gen[6664]),

			.SELF(gen[6568]),
			.cell_state(gen[6568])
		); 

/******************* CELL 6569 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6569 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6473]),
			.N(gen[6474]),
			.NE(gen[6475]),

			.O(gen[6568]),
			.E(gen[6570]),

			.SO(gen[6663]),
			.S(gen[6664]),
			.SE(gen[6665]),

			.SELF(gen[6569]),
			.cell_state(gen[6569])
		); 

/******************* CELL 6570 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6570 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6474]),
			.N(gen[6475]),
			.NE(gen[6476]),

			.O(gen[6569]),
			.E(gen[6571]),

			.SO(gen[6664]),
			.S(gen[6665]),
			.SE(gen[6666]),

			.SELF(gen[6570]),
			.cell_state(gen[6570])
		); 

/******************* CELL 6571 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6571 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6475]),
			.N(gen[6476]),
			.NE(gen[6477]),

			.O(gen[6570]),
			.E(gen[6572]),

			.SO(gen[6665]),
			.S(gen[6666]),
			.SE(gen[6667]),

			.SELF(gen[6571]),
			.cell_state(gen[6571])
		); 

/******************* CELL 6572 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6572 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6476]),
			.N(gen[6477]),
			.NE(gen[6478]),

			.O(gen[6571]),
			.E(gen[6573]),

			.SO(gen[6666]),
			.S(gen[6667]),
			.SE(gen[6668]),

			.SELF(gen[6572]),
			.cell_state(gen[6572])
		); 

/******************* CELL 6573 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6573 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6477]),
			.N(gen[6478]),
			.NE(gen[6479]),

			.O(gen[6572]),
			.E(gen[6574]),

			.SO(gen[6667]),
			.S(gen[6668]),
			.SE(gen[6669]),

			.SELF(gen[6573]),
			.cell_state(gen[6573])
		); 

/******************* CELL 6574 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6574 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6478]),
			.N(gen[6479]),
			.NE(gen[6480]),

			.O(gen[6573]),
			.E(gen[6575]),

			.SO(gen[6668]),
			.S(gen[6669]),
			.SE(gen[6670]),

			.SELF(gen[6574]),
			.cell_state(gen[6574])
		); 

/******************* CELL 6575 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6575 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6479]),
			.N(gen[6480]),
			.NE(gen[6481]),

			.O(gen[6574]),
			.E(gen[6576]),

			.SO(gen[6669]),
			.S(gen[6670]),
			.SE(gen[6671]),

			.SELF(gen[6575]),
			.cell_state(gen[6575])
		); 

/******************* CELL 6576 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6576 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6480]),
			.N(gen[6481]),
			.NE(gen[6482]),

			.O(gen[6575]),
			.E(gen[6577]),

			.SO(gen[6670]),
			.S(gen[6671]),
			.SE(gen[6672]),

			.SELF(gen[6576]),
			.cell_state(gen[6576])
		); 

/******************* CELL 6577 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6577 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6481]),
			.N(gen[6482]),
			.NE(gen[6483]),

			.O(gen[6576]),
			.E(gen[6578]),

			.SO(gen[6671]),
			.S(gen[6672]),
			.SE(gen[6673]),

			.SELF(gen[6577]),
			.cell_state(gen[6577])
		); 

/******************* CELL 6578 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6578 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6482]),
			.N(gen[6483]),
			.NE(gen[6484]),

			.O(gen[6577]),
			.E(gen[6579]),

			.SO(gen[6672]),
			.S(gen[6673]),
			.SE(gen[6674]),

			.SELF(gen[6578]),
			.cell_state(gen[6578])
		); 

/******************* CELL 6579 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6579 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6483]),
			.N(gen[6484]),
			.NE(gen[6485]),

			.O(gen[6578]),
			.E(gen[6580]),

			.SO(gen[6673]),
			.S(gen[6674]),
			.SE(gen[6675]),

			.SELF(gen[6579]),
			.cell_state(gen[6579])
		); 

/******************* CELL 6580 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6580 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6484]),
			.N(gen[6485]),
			.NE(gen[6486]),

			.O(gen[6579]),
			.E(gen[6581]),

			.SO(gen[6674]),
			.S(gen[6675]),
			.SE(gen[6676]),

			.SELF(gen[6580]),
			.cell_state(gen[6580])
		); 

/******************* CELL 6581 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6581 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6485]),
			.N(gen[6486]),
			.NE(gen[6487]),

			.O(gen[6580]),
			.E(gen[6582]),

			.SO(gen[6675]),
			.S(gen[6676]),
			.SE(gen[6677]),

			.SELF(gen[6581]),
			.cell_state(gen[6581])
		); 

/******************* CELL 6582 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6582 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6486]),
			.N(gen[6487]),
			.NE(gen[6488]),

			.O(gen[6581]),
			.E(gen[6583]),

			.SO(gen[6676]),
			.S(gen[6677]),
			.SE(gen[6678]),

			.SELF(gen[6582]),
			.cell_state(gen[6582])
		); 

/******************* CELL 6583 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6583 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6487]),
			.N(gen[6488]),
			.NE(gen[6489]),

			.O(gen[6582]),
			.E(gen[6584]),

			.SO(gen[6677]),
			.S(gen[6678]),
			.SE(gen[6679]),

			.SELF(gen[6583]),
			.cell_state(gen[6583])
		); 

/******************* CELL 6584 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6584 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6488]),
			.N(gen[6489]),
			.NE(gen[6490]),

			.O(gen[6583]),
			.E(gen[6585]),

			.SO(gen[6678]),
			.S(gen[6679]),
			.SE(gen[6680]),

			.SELF(gen[6584]),
			.cell_state(gen[6584])
		); 

/******************* CELL 6585 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6585 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6489]),
			.N(gen[6490]),
			.NE(gen[6491]),

			.O(gen[6584]),
			.E(gen[6586]),

			.SO(gen[6679]),
			.S(gen[6680]),
			.SE(gen[6681]),

			.SELF(gen[6585]),
			.cell_state(gen[6585])
		); 

/******************* CELL 6586 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6586 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6490]),
			.N(gen[6491]),
			.NE(gen[6492]),

			.O(gen[6585]),
			.E(gen[6587]),

			.SO(gen[6680]),
			.S(gen[6681]),
			.SE(gen[6682]),

			.SELF(gen[6586]),
			.cell_state(gen[6586])
		); 

/******************* CELL 6587 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6587 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6491]),
			.N(gen[6492]),
			.NE(gen[6493]),

			.O(gen[6586]),
			.E(gen[6588]),

			.SO(gen[6681]),
			.S(gen[6682]),
			.SE(gen[6683]),

			.SELF(gen[6587]),
			.cell_state(gen[6587])
		); 

/******************* CELL 6588 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6588 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6492]),
			.N(gen[6493]),
			.NE(gen[6494]),

			.O(gen[6587]),
			.E(gen[6589]),

			.SO(gen[6682]),
			.S(gen[6683]),
			.SE(gen[6684]),

			.SELF(gen[6588]),
			.cell_state(gen[6588])
		); 

/******************* CELL 6589 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6589 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6493]),
			.N(gen[6494]),
			.NE(gen[6495]),

			.O(gen[6588]),
			.E(gen[6590]),

			.SO(gen[6683]),
			.S(gen[6684]),
			.SE(gen[6685]),

			.SELF(gen[6589]),
			.cell_state(gen[6589])
		); 

/******************* CELL 6590 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6590 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6494]),
			.N(gen[6495]),
			.NE(gen[6496]),

			.O(gen[6589]),
			.E(gen[6591]),

			.SO(gen[6684]),
			.S(gen[6685]),
			.SE(gen[6686]),

			.SELF(gen[6590]),
			.cell_state(gen[6590])
		); 

/******************* CELL 6591 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6591 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6495]),
			.N(gen[6496]),
			.NE(gen[6497]),

			.O(gen[6590]),
			.E(gen[6592]),

			.SO(gen[6685]),
			.S(gen[6686]),
			.SE(gen[6687]),

			.SELF(gen[6591]),
			.cell_state(gen[6591])
		); 

/******************* CELL 6592 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6592 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6496]),
			.N(gen[6497]),
			.NE(gen[6498]),

			.O(gen[6591]),
			.E(gen[6593]),

			.SO(gen[6686]),
			.S(gen[6687]),
			.SE(gen[6688]),

			.SELF(gen[6592]),
			.cell_state(gen[6592])
		); 

/******************* CELL 6593 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6593 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6497]),
			.N(gen[6498]),
			.NE(gen[6499]),

			.O(gen[6592]),
			.E(gen[6594]),

			.SO(gen[6687]),
			.S(gen[6688]),
			.SE(gen[6689]),

			.SELF(gen[6593]),
			.cell_state(gen[6593])
		); 

/******************* CELL 6594 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6594 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6498]),
			.N(gen[6499]),
			.NE(gen[6500]),

			.O(gen[6593]),
			.E(gen[6595]),

			.SO(gen[6688]),
			.S(gen[6689]),
			.SE(gen[6690]),

			.SELF(gen[6594]),
			.cell_state(gen[6594])
		); 

/******************* CELL 6595 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6595 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6499]),
			.N(gen[6500]),
			.NE(gen[6501]),

			.O(gen[6594]),
			.E(gen[6596]),

			.SO(gen[6689]),
			.S(gen[6690]),
			.SE(gen[6691]),

			.SELF(gen[6595]),
			.cell_state(gen[6595])
		); 

/******************* CELL 6596 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6596 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6500]),
			.N(gen[6501]),
			.NE(gen[6502]),

			.O(gen[6595]),
			.E(gen[6597]),

			.SO(gen[6690]),
			.S(gen[6691]),
			.SE(gen[6692]),

			.SELF(gen[6596]),
			.cell_state(gen[6596])
		); 

/******************* CELL 6597 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6597 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6501]),
			.N(gen[6502]),
			.NE(gen[6503]),

			.O(gen[6596]),
			.E(gen[6598]),

			.SO(gen[6691]),
			.S(gen[6692]),
			.SE(gen[6693]),

			.SELF(gen[6597]),
			.cell_state(gen[6597])
		); 

/******************* CELL 6598 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6598 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6502]),
			.N(gen[6503]),
			.NE(gen[6504]),

			.O(gen[6597]),
			.E(gen[6599]),

			.SO(gen[6692]),
			.S(gen[6693]),
			.SE(gen[6694]),

			.SELF(gen[6598]),
			.cell_state(gen[6598])
		); 

/******************* CELL 6599 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6599 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6503]),
			.N(gen[6504]),
			.NE(gen[6505]),

			.O(gen[6598]),
			.E(gen[6600]),

			.SO(gen[6693]),
			.S(gen[6694]),
			.SE(gen[6695]),

			.SELF(gen[6599]),
			.cell_state(gen[6599])
		); 

/******************* CELL 6600 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6600 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6504]),
			.N(gen[6505]),
			.NE(gen[6506]),

			.O(gen[6599]),
			.E(gen[6601]),

			.SO(gen[6694]),
			.S(gen[6695]),
			.SE(gen[6696]),

			.SELF(gen[6600]),
			.cell_state(gen[6600])
		); 

/******************* CELL 6601 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6601 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6505]),
			.N(gen[6506]),
			.NE(gen[6507]),

			.O(gen[6600]),
			.E(gen[6602]),

			.SO(gen[6695]),
			.S(gen[6696]),
			.SE(gen[6697]),

			.SELF(gen[6601]),
			.cell_state(gen[6601])
		); 

/******************* CELL 6602 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6602 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6506]),
			.N(gen[6507]),
			.NE(gen[6508]),

			.O(gen[6601]),
			.E(gen[6603]),

			.SO(gen[6696]),
			.S(gen[6697]),
			.SE(gen[6698]),

			.SELF(gen[6602]),
			.cell_state(gen[6602])
		); 

/******************* CELL 6603 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6603 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6507]),
			.N(gen[6508]),
			.NE(gen[6509]),

			.O(gen[6602]),
			.E(gen[6604]),

			.SO(gen[6697]),
			.S(gen[6698]),
			.SE(gen[6699]),

			.SELF(gen[6603]),
			.cell_state(gen[6603])
		); 

/******************* CELL 6604 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6604 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6508]),
			.N(gen[6509]),
			.NE(gen[6510]),

			.O(gen[6603]),
			.E(gen[6605]),

			.SO(gen[6698]),
			.S(gen[6699]),
			.SE(gen[6700]),

			.SELF(gen[6604]),
			.cell_state(gen[6604])
		); 

/******************* CELL 6605 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6605 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6509]),
			.N(gen[6510]),
			.NE(gen[6511]),

			.O(gen[6604]),
			.E(gen[6606]),

			.SO(gen[6699]),
			.S(gen[6700]),
			.SE(gen[6701]),

			.SELF(gen[6605]),
			.cell_state(gen[6605])
		); 

/******************* CELL 6606 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6606 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6510]),
			.N(gen[6511]),
			.NE(gen[6512]),

			.O(gen[6605]),
			.E(gen[6607]),

			.SO(gen[6700]),
			.S(gen[6701]),
			.SE(gen[6702]),

			.SELF(gen[6606]),
			.cell_state(gen[6606])
		); 

/******************* CELL 6607 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6607 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6511]),
			.N(gen[6512]),
			.NE(gen[6513]),

			.O(gen[6606]),
			.E(gen[6608]),

			.SO(gen[6701]),
			.S(gen[6702]),
			.SE(gen[6703]),

			.SELF(gen[6607]),
			.cell_state(gen[6607])
		); 

/******************* CELL 6608 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6608 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6512]),
			.N(gen[6513]),
			.NE(gen[6514]),

			.O(gen[6607]),
			.E(gen[6609]),

			.SO(gen[6702]),
			.S(gen[6703]),
			.SE(gen[6704]),

			.SELF(gen[6608]),
			.cell_state(gen[6608])
		); 

/******************* CELL 6609 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6609 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6513]),
			.N(gen[6514]),
			.NE(gen[6515]),

			.O(gen[6608]),
			.E(gen[6610]),

			.SO(gen[6703]),
			.S(gen[6704]),
			.SE(gen[6705]),

			.SELF(gen[6609]),
			.cell_state(gen[6609])
		); 

/******************* CELL 6610 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6610 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6514]),
			.N(gen[6515]),
			.NE(gen[6516]),

			.O(gen[6609]),
			.E(gen[6611]),

			.SO(gen[6704]),
			.S(gen[6705]),
			.SE(gen[6706]),

			.SELF(gen[6610]),
			.cell_state(gen[6610])
		); 

/******************* CELL 6611 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6611 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6515]),
			.N(gen[6516]),
			.NE(gen[6517]),

			.O(gen[6610]),
			.E(gen[6612]),

			.SO(gen[6705]),
			.S(gen[6706]),
			.SE(gen[6707]),

			.SELF(gen[6611]),
			.cell_state(gen[6611])
		); 

/******************* CELL 6612 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6612 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6516]),
			.N(gen[6517]),
			.NE(gen[6518]),

			.O(gen[6611]),
			.E(gen[6613]),

			.SO(gen[6706]),
			.S(gen[6707]),
			.SE(gen[6708]),

			.SELF(gen[6612]),
			.cell_state(gen[6612])
		); 

/******************* CELL 6613 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6613 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6517]),
			.N(gen[6518]),
			.NE(gen[6519]),

			.O(gen[6612]),
			.E(gen[6614]),

			.SO(gen[6707]),
			.S(gen[6708]),
			.SE(gen[6709]),

			.SELF(gen[6613]),
			.cell_state(gen[6613])
		); 

/******************* CELL 6614 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6614 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6518]),
			.N(gen[6519]),
			.NE(gen[6520]),

			.O(gen[6613]),
			.E(gen[6615]),

			.SO(gen[6708]),
			.S(gen[6709]),
			.SE(gen[6710]),

			.SELF(gen[6614]),
			.cell_state(gen[6614])
		); 

/******************* CELL 6615 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6615 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6519]),
			.N(gen[6520]),
			.NE(gen[6521]),

			.O(gen[6614]),
			.E(gen[6616]),

			.SO(gen[6709]),
			.S(gen[6710]),
			.SE(gen[6711]),

			.SELF(gen[6615]),
			.cell_state(gen[6615])
		); 

/******************* CELL 6616 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6616 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6520]),
			.N(gen[6521]),
			.NE(gen[6522]),

			.O(gen[6615]),
			.E(gen[6617]),

			.SO(gen[6710]),
			.S(gen[6711]),
			.SE(gen[6712]),

			.SELF(gen[6616]),
			.cell_state(gen[6616])
		); 

/******************* CELL 6617 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6617 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6521]),
			.N(gen[6522]),
			.NE(gen[6523]),

			.O(gen[6616]),
			.E(gen[6618]),

			.SO(gen[6711]),
			.S(gen[6712]),
			.SE(gen[6713]),

			.SELF(gen[6617]),
			.cell_state(gen[6617])
		); 

/******************* CELL 6618 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6618 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6522]),
			.N(gen[6523]),
			.NE(gen[6524]),

			.O(gen[6617]),
			.E(gen[6619]),

			.SO(gen[6712]),
			.S(gen[6713]),
			.SE(gen[6714]),

			.SELF(gen[6618]),
			.cell_state(gen[6618])
		); 

/******************* CELL 6619 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6619 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6523]),
			.N(gen[6524]),
			.NE(gen[6525]),

			.O(gen[6618]),
			.E(gen[6620]),

			.SO(gen[6713]),
			.S(gen[6714]),
			.SE(gen[6715]),

			.SELF(gen[6619]),
			.cell_state(gen[6619])
		); 

/******************* CELL 6620 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6620 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6524]),
			.N(gen[6525]),
			.NE(gen[6526]),

			.O(gen[6619]),
			.E(gen[6621]),

			.SO(gen[6714]),
			.S(gen[6715]),
			.SE(gen[6716]),

			.SELF(gen[6620]),
			.cell_state(gen[6620])
		); 

/******************* CELL 6621 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6621 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6525]),
			.N(gen[6526]),
			.NE(gen[6527]),

			.O(gen[6620]),
			.E(gen[6622]),

			.SO(gen[6715]),
			.S(gen[6716]),
			.SE(gen[6717]),

			.SELF(gen[6621]),
			.cell_state(gen[6621])
		); 

/******************* CELL 6622 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6622 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6526]),
			.N(gen[6527]),
			.NE(gen[6528]),

			.O(gen[6621]),
			.E(gen[6623]),

			.SO(gen[6716]),
			.S(gen[6717]),
			.SE(gen[6718]),

			.SELF(gen[6622]),
			.cell_state(gen[6622])
		); 

/******************* CELL 6623 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6623 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6527]),
			.N(gen[6528]),
			.NE(gen[6529]),

			.O(gen[6622]),
			.E(gen[6624]),

			.SO(gen[6717]),
			.S(gen[6718]),
			.SE(gen[6719]),

			.SELF(gen[6623]),
			.cell_state(gen[6623])
		); 

/******************* CELL 6624 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6624 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6528]),
			.N(gen[6529]),
			.NE(gen[6530]),

			.O(gen[6623]),
			.E(gen[6625]),

			.SO(gen[6718]),
			.S(gen[6719]),
			.SE(gen[6720]),

			.SELF(gen[6624]),
			.cell_state(gen[6624])
		); 

/******************* CELL 6625 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6625 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6529]),
			.N(gen[6530]),
			.NE(gen[6531]),

			.O(gen[6624]),
			.E(gen[6626]),

			.SO(gen[6719]),
			.S(gen[6720]),
			.SE(gen[6721]),

			.SELF(gen[6625]),
			.cell_state(gen[6625])
		); 

/******************* CELL 6626 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6626 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6530]),
			.N(gen[6531]),
			.NE(gen[6532]),

			.O(gen[6625]),
			.E(gen[6627]),

			.SO(gen[6720]),
			.S(gen[6721]),
			.SE(gen[6722]),

			.SELF(gen[6626]),
			.cell_state(gen[6626])
		); 

/******************* CELL 6627 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6627 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6531]),
			.N(gen[6532]),
			.NE(gen[6533]),

			.O(gen[6626]),
			.E(gen[6628]),

			.SO(gen[6721]),
			.S(gen[6722]),
			.SE(gen[6723]),

			.SELF(gen[6627]),
			.cell_state(gen[6627])
		); 

/******************* CELL 6628 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6628 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6532]),
			.N(gen[6533]),
			.NE(gen[6534]),

			.O(gen[6627]),
			.E(gen[6629]),

			.SO(gen[6722]),
			.S(gen[6723]),
			.SE(gen[6724]),

			.SELF(gen[6628]),
			.cell_state(gen[6628])
		); 

/******************* CELL 6629 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6629 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6533]),
			.N(gen[6534]),
			.NE(gen[6535]),

			.O(gen[6628]),
			.E(gen[6630]),

			.SO(gen[6723]),
			.S(gen[6724]),
			.SE(gen[6725]),

			.SELF(gen[6629]),
			.cell_state(gen[6629])
		); 

/******************* CELL 6630 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6630 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6534]),
			.N(gen[6535]),
			.NE(gen[6536]),

			.O(gen[6629]),
			.E(gen[6631]),

			.SO(gen[6724]),
			.S(gen[6725]),
			.SE(gen[6726]),

			.SELF(gen[6630]),
			.cell_state(gen[6630])
		); 

/******************* CELL 6631 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6631 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6535]),
			.N(gen[6536]),
			.NE(gen[6537]),

			.O(gen[6630]),
			.E(gen[6632]),

			.SO(gen[6725]),
			.S(gen[6726]),
			.SE(gen[6727]),

			.SELF(gen[6631]),
			.cell_state(gen[6631])
		); 

/******************* CELL 6632 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6632 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6536]),
			.N(gen[6537]),
			.NE(gen[6538]),

			.O(gen[6631]),
			.E(gen[6633]),

			.SO(gen[6726]),
			.S(gen[6727]),
			.SE(gen[6728]),

			.SELF(gen[6632]),
			.cell_state(gen[6632])
		); 

/******************* CELL 6633 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6633 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6537]),
			.N(gen[6538]),
			.NE(gen[6539]),

			.O(gen[6632]),
			.E(gen[6634]),

			.SO(gen[6727]),
			.S(gen[6728]),
			.SE(gen[6729]),

			.SELF(gen[6633]),
			.cell_state(gen[6633])
		); 

/******************* CELL 6634 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6634 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6538]),
			.N(gen[6539]),
			.NE(gen[6540]),

			.O(gen[6633]),
			.E(gen[6635]),

			.SO(gen[6728]),
			.S(gen[6729]),
			.SE(gen[6730]),

			.SELF(gen[6634]),
			.cell_state(gen[6634])
		); 

/******************* CELL 6635 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6635 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6539]),
			.N(gen[6540]),
			.NE(gen[6541]),

			.O(gen[6634]),
			.E(gen[6636]),

			.SO(gen[6729]),
			.S(gen[6730]),
			.SE(gen[6731]),

			.SELF(gen[6635]),
			.cell_state(gen[6635])
		); 

/******************* CELL 6636 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6636 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6540]),
			.N(gen[6541]),
			.NE(gen[6542]),

			.O(gen[6635]),
			.E(gen[6637]),

			.SO(gen[6730]),
			.S(gen[6731]),
			.SE(gen[6732]),

			.SELF(gen[6636]),
			.cell_state(gen[6636])
		); 

/******************* CELL 6637 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6637 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6541]),
			.N(gen[6542]),
			.NE(gen[6543]),

			.O(gen[6636]),
			.E(gen[6638]),

			.SO(gen[6731]),
			.S(gen[6732]),
			.SE(gen[6733]),

			.SELF(gen[6637]),
			.cell_state(gen[6637])
		); 

/******************* CELL 6638 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6638 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6542]),
			.N(gen[6543]),
			.NE(gen[6544]),

			.O(gen[6637]),
			.E(gen[6639]),

			.SO(gen[6732]),
			.S(gen[6733]),
			.SE(gen[6734]),

			.SELF(gen[6638]),
			.cell_state(gen[6638])
		); 

/******************* CELL 6639 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6639 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6543]),
			.N(gen[6544]),
			.NE(gen[6545]),

			.O(gen[6638]),
			.E(gen[6640]),

			.SO(gen[6733]),
			.S(gen[6734]),
			.SE(gen[6735]),

			.SELF(gen[6639]),
			.cell_state(gen[6639])
		); 

/******************* CELL 6640 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6640 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6544]),
			.N(gen[6545]),
			.NE(gen[6546]),

			.O(gen[6639]),
			.E(gen[6641]),

			.SO(gen[6734]),
			.S(gen[6735]),
			.SE(gen[6736]),

			.SELF(gen[6640]),
			.cell_state(gen[6640])
		); 

/******************* CELL 6641 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6641 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6545]),
			.N(gen[6546]),
			.NE(gen[6547]),

			.O(gen[6640]),
			.E(gen[6642]),

			.SO(gen[6735]),
			.S(gen[6736]),
			.SE(gen[6737]),

			.SELF(gen[6641]),
			.cell_state(gen[6641])
		); 

/******************* CELL 6642 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6642 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6546]),
			.N(gen[6547]),
			.NE(gen[6548]),

			.O(gen[6641]),
			.E(gen[6643]),

			.SO(gen[6736]),
			.S(gen[6737]),
			.SE(gen[6738]),

			.SELF(gen[6642]),
			.cell_state(gen[6642])
		); 

/******************* CELL 6643 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6643 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6547]),
			.N(gen[6548]),
			.NE(gen[6549]),

			.O(gen[6642]),
			.E(gen[6644]),

			.SO(gen[6737]),
			.S(gen[6738]),
			.SE(gen[6739]),

			.SELF(gen[6643]),
			.cell_state(gen[6643])
		); 

/******************* CELL 6644 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6644 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6548]),
			.N(gen[6549]),
			.NE(gen[6550]),

			.O(gen[6643]),
			.E(gen[6645]),

			.SO(gen[6738]),
			.S(gen[6739]),
			.SE(gen[6740]),

			.SELF(gen[6644]),
			.cell_state(gen[6644])
		); 

/******************* CELL 6645 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6645 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6549]),
			.N(gen[6550]),
			.NE(gen[6551]),

			.O(gen[6644]),
			.E(gen[6646]),

			.SO(gen[6739]),
			.S(gen[6740]),
			.SE(gen[6741]),

			.SELF(gen[6645]),
			.cell_state(gen[6645])
		); 

/******************* CELL 6646 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6646 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6550]),
			.N(gen[6551]),
			.NE(gen[6552]),

			.O(gen[6645]),
			.E(gen[6647]),

			.SO(gen[6740]),
			.S(gen[6741]),
			.SE(gen[6742]),

			.SELF(gen[6646]),
			.cell_state(gen[6646])
		); 

/******************* CELL 6647 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6647 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6551]),
			.N(gen[6552]),
			.NE(gen[6553]),

			.O(gen[6646]),
			.E(gen[6648]),

			.SO(gen[6741]),
			.S(gen[6742]),
			.SE(gen[6743]),

			.SELF(gen[6647]),
			.cell_state(gen[6647])
		); 

/******************* CELL 6648 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6648 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6552]),
			.N(gen[6553]),
			.NE(gen[6554]),

			.O(gen[6647]),
			.E(gen[6649]),

			.SO(gen[6742]),
			.S(gen[6743]),
			.SE(gen[6744]),

			.SELF(gen[6648]),
			.cell_state(gen[6648])
		); 

/******************* CELL 6649 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6649 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6553]),
			.N(gen[6554]),
			.NE(gen[6553]),

			.O(gen[6648]),
			.E(gen[6648]),

			.SO(gen[6743]),
			.S(gen[6744]),
			.SE(gen[6743]),

			.SELF(gen[6649]),
			.cell_state(gen[6649])
		); 

/******************* CELL 6650 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6650 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6556]),
			.N(gen[6555]),
			.NE(gen[6556]),

			.O(gen[6651]),
			.E(gen[6651]),

			.SO(gen[6746]),
			.S(gen[6745]),
			.SE(gen[6746]),

			.SELF(gen[6650]),
			.cell_state(gen[6650])
		); 

/******************* CELL 6651 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6651 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6555]),
			.N(gen[6556]),
			.NE(gen[6557]),

			.O(gen[6650]),
			.E(gen[6652]),

			.SO(gen[6745]),
			.S(gen[6746]),
			.SE(gen[6747]),

			.SELF(gen[6651]),
			.cell_state(gen[6651])
		); 

/******************* CELL 6652 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6652 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6556]),
			.N(gen[6557]),
			.NE(gen[6558]),

			.O(gen[6651]),
			.E(gen[6653]),

			.SO(gen[6746]),
			.S(gen[6747]),
			.SE(gen[6748]),

			.SELF(gen[6652]),
			.cell_state(gen[6652])
		); 

/******************* CELL 6653 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6653 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6557]),
			.N(gen[6558]),
			.NE(gen[6559]),

			.O(gen[6652]),
			.E(gen[6654]),

			.SO(gen[6747]),
			.S(gen[6748]),
			.SE(gen[6749]),

			.SELF(gen[6653]),
			.cell_state(gen[6653])
		); 

/******************* CELL 6654 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6654 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6558]),
			.N(gen[6559]),
			.NE(gen[6560]),

			.O(gen[6653]),
			.E(gen[6655]),

			.SO(gen[6748]),
			.S(gen[6749]),
			.SE(gen[6750]),

			.SELF(gen[6654]),
			.cell_state(gen[6654])
		); 

/******************* CELL 6655 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6655 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6559]),
			.N(gen[6560]),
			.NE(gen[6561]),

			.O(gen[6654]),
			.E(gen[6656]),

			.SO(gen[6749]),
			.S(gen[6750]),
			.SE(gen[6751]),

			.SELF(gen[6655]),
			.cell_state(gen[6655])
		); 

/******************* CELL 6656 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6656 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6560]),
			.N(gen[6561]),
			.NE(gen[6562]),

			.O(gen[6655]),
			.E(gen[6657]),

			.SO(gen[6750]),
			.S(gen[6751]),
			.SE(gen[6752]),

			.SELF(gen[6656]),
			.cell_state(gen[6656])
		); 

/******************* CELL 6657 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6657 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6561]),
			.N(gen[6562]),
			.NE(gen[6563]),

			.O(gen[6656]),
			.E(gen[6658]),

			.SO(gen[6751]),
			.S(gen[6752]),
			.SE(gen[6753]),

			.SELF(gen[6657]),
			.cell_state(gen[6657])
		); 

/******************* CELL 6658 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6658 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6562]),
			.N(gen[6563]),
			.NE(gen[6564]),

			.O(gen[6657]),
			.E(gen[6659]),

			.SO(gen[6752]),
			.S(gen[6753]),
			.SE(gen[6754]),

			.SELF(gen[6658]),
			.cell_state(gen[6658])
		); 

/******************* CELL 6659 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6659 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6563]),
			.N(gen[6564]),
			.NE(gen[6565]),

			.O(gen[6658]),
			.E(gen[6660]),

			.SO(gen[6753]),
			.S(gen[6754]),
			.SE(gen[6755]),

			.SELF(gen[6659]),
			.cell_state(gen[6659])
		); 

/******************* CELL 6660 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6660 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6564]),
			.N(gen[6565]),
			.NE(gen[6566]),

			.O(gen[6659]),
			.E(gen[6661]),

			.SO(gen[6754]),
			.S(gen[6755]),
			.SE(gen[6756]),

			.SELF(gen[6660]),
			.cell_state(gen[6660])
		); 

/******************* CELL 6661 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6661 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6565]),
			.N(gen[6566]),
			.NE(gen[6567]),

			.O(gen[6660]),
			.E(gen[6662]),

			.SO(gen[6755]),
			.S(gen[6756]),
			.SE(gen[6757]),

			.SELF(gen[6661]),
			.cell_state(gen[6661])
		); 

/******************* CELL 6662 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6662 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6566]),
			.N(gen[6567]),
			.NE(gen[6568]),

			.O(gen[6661]),
			.E(gen[6663]),

			.SO(gen[6756]),
			.S(gen[6757]),
			.SE(gen[6758]),

			.SELF(gen[6662]),
			.cell_state(gen[6662])
		); 

/******************* CELL 6663 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6663 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6567]),
			.N(gen[6568]),
			.NE(gen[6569]),

			.O(gen[6662]),
			.E(gen[6664]),

			.SO(gen[6757]),
			.S(gen[6758]),
			.SE(gen[6759]),

			.SELF(gen[6663]),
			.cell_state(gen[6663])
		); 

/******************* CELL 6664 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6664 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6568]),
			.N(gen[6569]),
			.NE(gen[6570]),

			.O(gen[6663]),
			.E(gen[6665]),

			.SO(gen[6758]),
			.S(gen[6759]),
			.SE(gen[6760]),

			.SELF(gen[6664]),
			.cell_state(gen[6664])
		); 

/******************* CELL 6665 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6665 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6569]),
			.N(gen[6570]),
			.NE(gen[6571]),

			.O(gen[6664]),
			.E(gen[6666]),

			.SO(gen[6759]),
			.S(gen[6760]),
			.SE(gen[6761]),

			.SELF(gen[6665]),
			.cell_state(gen[6665])
		); 

/******************* CELL 6666 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6666 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6570]),
			.N(gen[6571]),
			.NE(gen[6572]),

			.O(gen[6665]),
			.E(gen[6667]),

			.SO(gen[6760]),
			.S(gen[6761]),
			.SE(gen[6762]),

			.SELF(gen[6666]),
			.cell_state(gen[6666])
		); 

/******************* CELL 6667 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6667 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6571]),
			.N(gen[6572]),
			.NE(gen[6573]),

			.O(gen[6666]),
			.E(gen[6668]),

			.SO(gen[6761]),
			.S(gen[6762]),
			.SE(gen[6763]),

			.SELF(gen[6667]),
			.cell_state(gen[6667])
		); 

/******************* CELL 6668 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6668 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6572]),
			.N(gen[6573]),
			.NE(gen[6574]),

			.O(gen[6667]),
			.E(gen[6669]),

			.SO(gen[6762]),
			.S(gen[6763]),
			.SE(gen[6764]),

			.SELF(gen[6668]),
			.cell_state(gen[6668])
		); 

/******************* CELL 6669 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6669 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6573]),
			.N(gen[6574]),
			.NE(gen[6575]),

			.O(gen[6668]),
			.E(gen[6670]),

			.SO(gen[6763]),
			.S(gen[6764]),
			.SE(gen[6765]),

			.SELF(gen[6669]),
			.cell_state(gen[6669])
		); 

/******************* CELL 6670 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6670 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6574]),
			.N(gen[6575]),
			.NE(gen[6576]),

			.O(gen[6669]),
			.E(gen[6671]),

			.SO(gen[6764]),
			.S(gen[6765]),
			.SE(gen[6766]),

			.SELF(gen[6670]),
			.cell_state(gen[6670])
		); 

/******************* CELL 6671 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6671 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6575]),
			.N(gen[6576]),
			.NE(gen[6577]),

			.O(gen[6670]),
			.E(gen[6672]),

			.SO(gen[6765]),
			.S(gen[6766]),
			.SE(gen[6767]),

			.SELF(gen[6671]),
			.cell_state(gen[6671])
		); 

/******************* CELL 6672 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6672 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6576]),
			.N(gen[6577]),
			.NE(gen[6578]),

			.O(gen[6671]),
			.E(gen[6673]),

			.SO(gen[6766]),
			.S(gen[6767]),
			.SE(gen[6768]),

			.SELF(gen[6672]),
			.cell_state(gen[6672])
		); 

/******************* CELL 6673 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6673 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6577]),
			.N(gen[6578]),
			.NE(gen[6579]),

			.O(gen[6672]),
			.E(gen[6674]),

			.SO(gen[6767]),
			.S(gen[6768]),
			.SE(gen[6769]),

			.SELF(gen[6673]),
			.cell_state(gen[6673])
		); 

/******************* CELL 6674 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6674 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6578]),
			.N(gen[6579]),
			.NE(gen[6580]),

			.O(gen[6673]),
			.E(gen[6675]),

			.SO(gen[6768]),
			.S(gen[6769]),
			.SE(gen[6770]),

			.SELF(gen[6674]),
			.cell_state(gen[6674])
		); 

/******************* CELL 6675 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6675 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6579]),
			.N(gen[6580]),
			.NE(gen[6581]),

			.O(gen[6674]),
			.E(gen[6676]),

			.SO(gen[6769]),
			.S(gen[6770]),
			.SE(gen[6771]),

			.SELF(gen[6675]),
			.cell_state(gen[6675])
		); 

/******************* CELL 6676 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6676 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6580]),
			.N(gen[6581]),
			.NE(gen[6582]),

			.O(gen[6675]),
			.E(gen[6677]),

			.SO(gen[6770]),
			.S(gen[6771]),
			.SE(gen[6772]),

			.SELF(gen[6676]),
			.cell_state(gen[6676])
		); 

/******************* CELL 6677 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6677 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6581]),
			.N(gen[6582]),
			.NE(gen[6583]),

			.O(gen[6676]),
			.E(gen[6678]),

			.SO(gen[6771]),
			.S(gen[6772]),
			.SE(gen[6773]),

			.SELF(gen[6677]),
			.cell_state(gen[6677])
		); 

/******************* CELL 6678 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6678 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6582]),
			.N(gen[6583]),
			.NE(gen[6584]),

			.O(gen[6677]),
			.E(gen[6679]),

			.SO(gen[6772]),
			.S(gen[6773]),
			.SE(gen[6774]),

			.SELF(gen[6678]),
			.cell_state(gen[6678])
		); 

/******************* CELL 6679 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6679 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6583]),
			.N(gen[6584]),
			.NE(gen[6585]),

			.O(gen[6678]),
			.E(gen[6680]),

			.SO(gen[6773]),
			.S(gen[6774]),
			.SE(gen[6775]),

			.SELF(gen[6679]),
			.cell_state(gen[6679])
		); 

/******************* CELL 6680 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6680 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6584]),
			.N(gen[6585]),
			.NE(gen[6586]),

			.O(gen[6679]),
			.E(gen[6681]),

			.SO(gen[6774]),
			.S(gen[6775]),
			.SE(gen[6776]),

			.SELF(gen[6680]),
			.cell_state(gen[6680])
		); 

/******************* CELL 6681 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6681 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6585]),
			.N(gen[6586]),
			.NE(gen[6587]),

			.O(gen[6680]),
			.E(gen[6682]),

			.SO(gen[6775]),
			.S(gen[6776]),
			.SE(gen[6777]),

			.SELF(gen[6681]),
			.cell_state(gen[6681])
		); 

/******************* CELL 6682 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6682 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6586]),
			.N(gen[6587]),
			.NE(gen[6588]),

			.O(gen[6681]),
			.E(gen[6683]),

			.SO(gen[6776]),
			.S(gen[6777]),
			.SE(gen[6778]),

			.SELF(gen[6682]),
			.cell_state(gen[6682])
		); 

/******************* CELL 6683 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6683 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6587]),
			.N(gen[6588]),
			.NE(gen[6589]),

			.O(gen[6682]),
			.E(gen[6684]),

			.SO(gen[6777]),
			.S(gen[6778]),
			.SE(gen[6779]),

			.SELF(gen[6683]),
			.cell_state(gen[6683])
		); 

/******************* CELL 6684 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6684 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6588]),
			.N(gen[6589]),
			.NE(gen[6590]),

			.O(gen[6683]),
			.E(gen[6685]),

			.SO(gen[6778]),
			.S(gen[6779]),
			.SE(gen[6780]),

			.SELF(gen[6684]),
			.cell_state(gen[6684])
		); 

/******************* CELL 6685 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6685 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6589]),
			.N(gen[6590]),
			.NE(gen[6591]),

			.O(gen[6684]),
			.E(gen[6686]),

			.SO(gen[6779]),
			.S(gen[6780]),
			.SE(gen[6781]),

			.SELF(gen[6685]),
			.cell_state(gen[6685])
		); 

/******************* CELL 6686 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6686 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6590]),
			.N(gen[6591]),
			.NE(gen[6592]),

			.O(gen[6685]),
			.E(gen[6687]),

			.SO(gen[6780]),
			.S(gen[6781]),
			.SE(gen[6782]),

			.SELF(gen[6686]),
			.cell_state(gen[6686])
		); 

/******************* CELL 6687 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6687 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6591]),
			.N(gen[6592]),
			.NE(gen[6593]),

			.O(gen[6686]),
			.E(gen[6688]),

			.SO(gen[6781]),
			.S(gen[6782]),
			.SE(gen[6783]),

			.SELF(gen[6687]),
			.cell_state(gen[6687])
		); 

/******************* CELL 6688 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6688 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6592]),
			.N(gen[6593]),
			.NE(gen[6594]),

			.O(gen[6687]),
			.E(gen[6689]),

			.SO(gen[6782]),
			.S(gen[6783]),
			.SE(gen[6784]),

			.SELF(gen[6688]),
			.cell_state(gen[6688])
		); 

/******************* CELL 6689 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6689 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6593]),
			.N(gen[6594]),
			.NE(gen[6595]),

			.O(gen[6688]),
			.E(gen[6690]),

			.SO(gen[6783]),
			.S(gen[6784]),
			.SE(gen[6785]),

			.SELF(gen[6689]),
			.cell_state(gen[6689])
		); 

/******************* CELL 6690 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6690 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6594]),
			.N(gen[6595]),
			.NE(gen[6596]),

			.O(gen[6689]),
			.E(gen[6691]),

			.SO(gen[6784]),
			.S(gen[6785]),
			.SE(gen[6786]),

			.SELF(gen[6690]),
			.cell_state(gen[6690])
		); 

/******************* CELL 6691 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6691 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6595]),
			.N(gen[6596]),
			.NE(gen[6597]),

			.O(gen[6690]),
			.E(gen[6692]),

			.SO(gen[6785]),
			.S(gen[6786]),
			.SE(gen[6787]),

			.SELF(gen[6691]),
			.cell_state(gen[6691])
		); 

/******************* CELL 6692 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6692 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6596]),
			.N(gen[6597]),
			.NE(gen[6598]),

			.O(gen[6691]),
			.E(gen[6693]),

			.SO(gen[6786]),
			.S(gen[6787]),
			.SE(gen[6788]),

			.SELF(gen[6692]),
			.cell_state(gen[6692])
		); 

/******************* CELL 6693 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6693 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6597]),
			.N(gen[6598]),
			.NE(gen[6599]),

			.O(gen[6692]),
			.E(gen[6694]),

			.SO(gen[6787]),
			.S(gen[6788]),
			.SE(gen[6789]),

			.SELF(gen[6693]),
			.cell_state(gen[6693])
		); 

/******************* CELL 6694 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6694 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6598]),
			.N(gen[6599]),
			.NE(gen[6600]),

			.O(gen[6693]),
			.E(gen[6695]),

			.SO(gen[6788]),
			.S(gen[6789]),
			.SE(gen[6790]),

			.SELF(gen[6694]),
			.cell_state(gen[6694])
		); 

/******************* CELL 6695 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6695 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6599]),
			.N(gen[6600]),
			.NE(gen[6601]),

			.O(gen[6694]),
			.E(gen[6696]),

			.SO(gen[6789]),
			.S(gen[6790]),
			.SE(gen[6791]),

			.SELF(gen[6695]),
			.cell_state(gen[6695])
		); 

/******************* CELL 6696 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6696 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6600]),
			.N(gen[6601]),
			.NE(gen[6602]),

			.O(gen[6695]),
			.E(gen[6697]),

			.SO(gen[6790]),
			.S(gen[6791]),
			.SE(gen[6792]),

			.SELF(gen[6696]),
			.cell_state(gen[6696])
		); 

/******************* CELL 6697 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6697 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6601]),
			.N(gen[6602]),
			.NE(gen[6603]),

			.O(gen[6696]),
			.E(gen[6698]),

			.SO(gen[6791]),
			.S(gen[6792]),
			.SE(gen[6793]),

			.SELF(gen[6697]),
			.cell_state(gen[6697])
		); 

/******************* CELL 6698 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6698 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6602]),
			.N(gen[6603]),
			.NE(gen[6604]),

			.O(gen[6697]),
			.E(gen[6699]),

			.SO(gen[6792]),
			.S(gen[6793]),
			.SE(gen[6794]),

			.SELF(gen[6698]),
			.cell_state(gen[6698])
		); 

/******************* CELL 6699 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6699 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6603]),
			.N(gen[6604]),
			.NE(gen[6605]),

			.O(gen[6698]),
			.E(gen[6700]),

			.SO(gen[6793]),
			.S(gen[6794]),
			.SE(gen[6795]),

			.SELF(gen[6699]),
			.cell_state(gen[6699])
		); 

/******************* CELL 6700 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6700 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6604]),
			.N(gen[6605]),
			.NE(gen[6606]),

			.O(gen[6699]),
			.E(gen[6701]),

			.SO(gen[6794]),
			.S(gen[6795]),
			.SE(gen[6796]),

			.SELF(gen[6700]),
			.cell_state(gen[6700])
		); 

/******************* CELL 6701 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6701 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6605]),
			.N(gen[6606]),
			.NE(gen[6607]),

			.O(gen[6700]),
			.E(gen[6702]),

			.SO(gen[6795]),
			.S(gen[6796]),
			.SE(gen[6797]),

			.SELF(gen[6701]),
			.cell_state(gen[6701])
		); 

/******************* CELL 6702 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6702 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6606]),
			.N(gen[6607]),
			.NE(gen[6608]),

			.O(gen[6701]),
			.E(gen[6703]),

			.SO(gen[6796]),
			.S(gen[6797]),
			.SE(gen[6798]),

			.SELF(gen[6702]),
			.cell_state(gen[6702])
		); 

/******************* CELL 6703 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6703 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6607]),
			.N(gen[6608]),
			.NE(gen[6609]),

			.O(gen[6702]),
			.E(gen[6704]),

			.SO(gen[6797]),
			.S(gen[6798]),
			.SE(gen[6799]),

			.SELF(gen[6703]),
			.cell_state(gen[6703])
		); 

/******************* CELL 6704 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6704 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6608]),
			.N(gen[6609]),
			.NE(gen[6610]),

			.O(gen[6703]),
			.E(gen[6705]),

			.SO(gen[6798]),
			.S(gen[6799]),
			.SE(gen[6800]),

			.SELF(gen[6704]),
			.cell_state(gen[6704])
		); 

/******************* CELL 6705 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6705 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6609]),
			.N(gen[6610]),
			.NE(gen[6611]),

			.O(gen[6704]),
			.E(gen[6706]),

			.SO(gen[6799]),
			.S(gen[6800]),
			.SE(gen[6801]),

			.SELF(gen[6705]),
			.cell_state(gen[6705])
		); 

/******************* CELL 6706 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6706 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6610]),
			.N(gen[6611]),
			.NE(gen[6612]),

			.O(gen[6705]),
			.E(gen[6707]),

			.SO(gen[6800]),
			.S(gen[6801]),
			.SE(gen[6802]),

			.SELF(gen[6706]),
			.cell_state(gen[6706])
		); 

/******************* CELL 6707 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6707 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6611]),
			.N(gen[6612]),
			.NE(gen[6613]),

			.O(gen[6706]),
			.E(gen[6708]),

			.SO(gen[6801]),
			.S(gen[6802]),
			.SE(gen[6803]),

			.SELF(gen[6707]),
			.cell_state(gen[6707])
		); 

/******************* CELL 6708 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6708 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6612]),
			.N(gen[6613]),
			.NE(gen[6614]),

			.O(gen[6707]),
			.E(gen[6709]),

			.SO(gen[6802]),
			.S(gen[6803]),
			.SE(gen[6804]),

			.SELF(gen[6708]),
			.cell_state(gen[6708])
		); 

/******************* CELL 6709 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6709 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6613]),
			.N(gen[6614]),
			.NE(gen[6615]),

			.O(gen[6708]),
			.E(gen[6710]),

			.SO(gen[6803]),
			.S(gen[6804]),
			.SE(gen[6805]),

			.SELF(gen[6709]),
			.cell_state(gen[6709])
		); 

/******************* CELL 6710 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6710 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6614]),
			.N(gen[6615]),
			.NE(gen[6616]),

			.O(gen[6709]),
			.E(gen[6711]),

			.SO(gen[6804]),
			.S(gen[6805]),
			.SE(gen[6806]),

			.SELF(gen[6710]),
			.cell_state(gen[6710])
		); 

/******************* CELL 6711 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6711 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6615]),
			.N(gen[6616]),
			.NE(gen[6617]),

			.O(gen[6710]),
			.E(gen[6712]),

			.SO(gen[6805]),
			.S(gen[6806]),
			.SE(gen[6807]),

			.SELF(gen[6711]),
			.cell_state(gen[6711])
		); 

/******************* CELL 6712 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6712 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6616]),
			.N(gen[6617]),
			.NE(gen[6618]),

			.O(gen[6711]),
			.E(gen[6713]),

			.SO(gen[6806]),
			.S(gen[6807]),
			.SE(gen[6808]),

			.SELF(gen[6712]),
			.cell_state(gen[6712])
		); 

/******************* CELL 6713 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6713 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6617]),
			.N(gen[6618]),
			.NE(gen[6619]),

			.O(gen[6712]),
			.E(gen[6714]),

			.SO(gen[6807]),
			.S(gen[6808]),
			.SE(gen[6809]),

			.SELF(gen[6713]),
			.cell_state(gen[6713])
		); 

/******************* CELL 6714 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6714 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6618]),
			.N(gen[6619]),
			.NE(gen[6620]),

			.O(gen[6713]),
			.E(gen[6715]),

			.SO(gen[6808]),
			.S(gen[6809]),
			.SE(gen[6810]),

			.SELF(gen[6714]),
			.cell_state(gen[6714])
		); 

/******************* CELL 6715 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6715 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6619]),
			.N(gen[6620]),
			.NE(gen[6621]),

			.O(gen[6714]),
			.E(gen[6716]),

			.SO(gen[6809]),
			.S(gen[6810]),
			.SE(gen[6811]),

			.SELF(gen[6715]),
			.cell_state(gen[6715])
		); 

/******************* CELL 6716 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6716 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6620]),
			.N(gen[6621]),
			.NE(gen[6622]),

			.O(gen[6715]),
			.E(gen[6717]),

			.SO(gen[6810]),
			.S(gen[6811]),
			.SE(gen[6812]),

			.SELF(gen[6716]),
			.cell_state(gen[6716])
		); 

/******************* CELL 6717 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6717 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6621]),
			.N(gen[6622]),
			.NE(gen[6623]),

			.O(gen[6716]),
			.E(gen[6718]),

			.SO(gen[6811]),
			.S(gen[6812]),
			.SE(gen[6813]),

			.SELF(gen[6717]),
			.cell_state(gen[6717])
		); 

/******************* CELL 6718 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6718 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6622]),
			.N(gen[6623]),
			.NE(gen[6624]),

			.O(gen[6717]),
			.E(gen[6719]),

			.SO(gen[6812]),
			.S(gen[6813]),
			.SE(gen[6814]),

			.SELF(gen[6718]),
			.cell_state(gen[6718])
		); 

/******************* CELL 6719 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6719 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6623]),
			.N(gen[6624]),
			.NE(gen[6625]),

			.O(gen[6718]),
			.E(gen[6720]),

			.SO(gen[6813]),
			.S(gen[6814]),
			.SE(gen[6815]),

			.SELF(gen[6719]),
			.cell_state(gen[6719])
		); 

/******************* CELL 6720 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6720 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6624]),
			.N(gen[6625]),
			.NE(gen[6626]),

			.O(gen[6719]),
			.E(gen[6721]),

			.SO(gen[6814]),
			.S(gen[6815]),
			.SE(gen[6816]),

			.SELF(gen[6720]),
			.cell_state(gen[6720])
		); 

/******************* CELL 6721 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6721 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6625]),
			.N(gen[6626]),
			.NE(gen[6627]),

			.O(gen[6720]),
			.E(gen[6722]),

			.SO(gen[6815]),
			.S(gen[6816]),
			.SE(gen[6817]),

			.SELF(gen[6721]),
			.cell_state(gen[6721])
		); 

/******************* CELL 6722 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6722 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6626]),
			.N(gen[6627]),
			.NE(gen[6628]),

			.O(gen[6721]),
			.E(gen[6723]),

			.SO(gen[6816]),
			.S(gen[6817]),
			.SE(gen[6818]),

			.SELF(gen[6722]),
			.cell_state(gen[6722])
		); 

/******************* CELL 6723 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6723 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6627]),
			.N(gen[6628]),
			.NE(gen[6629]),

			.O(gen[6722]),
			.E(gen[6724]),

			.SO(gen[6817]),
			.S(gen[6818]),
			.SE(gen[6819]),

			.SELF(gen[6723]),
			.cell_state(gen[6723])
		); 

/******************* CELL 6724 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6724 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6628]),
			.N(gen[6629]),
			.NE(gen[6630]),

			.O(gen[6723]),
			.E(gen[6725]),

			.SO(gen[6818]),
			.S(gen[6819]),
			.SE(gen[6820]),

			.SELF(gen[6724]),
			.cell_state(gen[6724])
		); 

/******************* CELL 6725 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6725 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6629]),
			.N(gen[6630]),
			.NE(gen[6631]),

			.O(gen[6724]),
			.E(gen[6726]),

			.SO(gen[6819]),
			.S(gen[6820]),
			.SE(gen[6821]),

			.SELF(gen[6725]),
			.cell_state(gen[6725])
		); 

/******************* CELL 6726 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6726 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6630]),
			.N(gen[6631]),
			.NE(gen[6632]),

			.O(gen[6725]),
			.E(gen[6727]),

			.SO(gen[6820]),
			.S(gen[6821]),
			.SE(gen[6822]),

			.SELF(gen[6726]),
			.cell_state(gen[6726])
		); 

/******************* CELL 6727 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6727 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6631]),
			.N(gen[6632]),
			.NE(gen[6633]),

			.O(gen[6726]),
			.E(gen[6728]),

			.SO(gen[6821]),
			.S(gen[6822]),
			.SE(gen[6823]),

			.SELF(gen[6727]),
			.cell_state(gen[6727])
		); 

/******************* CELL 6728 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6728 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6632]),
			.N(gen[6633]),
			.NE(gen[6634]),

			.O(gen[6727]),
			.E(gen[6729]),

			.SO(gen[6822]),
			.S(gen[6823]),
			.SE(gen[6824]),

			.SELF(gen[6728]),
			.cell_state(gen[6728])
		); 

/******************* CELL 6729 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6729 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6633]),
			.N(gen[6634]),
			.NE(gen[6635]),

			.O(gen[6728]),
			.E(gen[6730]),

			.SO(gen[6823]),
			.S(gen[6824]),
			.SE(gen[6825]),

			.SELF(gen[6729]),
			.cell_state(gen[6729])
		); 

/******************* CELL 6730 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6730 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6634]),
			.N(gen[6635]),
			.NE(gen[6636]),

			.O(gen[6729]),
			.E(gen[6731]),

			.SO(gen[6824]),
			.S(gen[6825]),
			.SE(gen[6826]),

			.SELF(gen[6730]),
			.cell_state(gen[6730])
		); 

/******************* CELL 6731 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6731 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6635]),
			.N(gen[6636]),
			.NE(gen[6637]),

			.O(gen[6730]),
			.E(gen[6732]),

			.SO(gen[6825]),
			.S(gen[6826]),
			.SE(gen[6827]),

			.SELF(gen[6731]),
			.cell_state(gen[6731])
		); 

/******************* CELL 6732 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6732 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6636]),
			.N(gen[6637]),
			.NE(gen[6638]),

			.O(gen[6731]),
			.E(gen[6733]),

			.SO(gen[6826]),
			.S(gen[6827]),
			.SE(gen[6828]),

			.SELF(gen[6732]),
			.cell_state(gen[6732])
		); 

/******************* CELL 6733 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6733 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6637]),
			.N(gen[6638]),
			.NE(gen[6639]),

			.O(gen[6732]),
			.E(gen[6734]),

			.SO(gen[6827]),
			.S(gen[6828]),
			.SE(gen[6829]),

			.SELF(gen[6733]),
			.cell_state(gen[6733])
		); 

/******************* CELL 6734 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6734 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6638]),
			.N(gen[6639]),
			.NE(gen[6640]),

			.O(gen[6733]),
			.E(gen[6735]),

			.SO(gen[6828]),
			.S(gen[6829]),
			.SE(gen[6830]),

			.SELF(gen[6734]),
			.cell_state(gen[6734])
		); 

/******************* CELL 6735 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6735 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6639]),
			.N(gen[6640]),
			.NE(gen[6641]),

			.O(gen[6734]),
			.E(gen[6736]),

			.SO(gen[6829]),
			.S(gen[6830]),
			.SE(gen[6831]),

			.SELF(gen[6735]),
			.cell_state(gen[6735])
		); 

/******************* CELL 6736 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6736 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6640]),
			.N(gen[6641]),
			.NE(gen[6642]),

			.O(gen[6735]),
			.E(gen[6737]),

			.SO(gen[6830]),
			.S(gen[6831]),
			.SE(gen[6832]),

			.SELF(gen[6736]),
			.cell_state(gen[6736])
		); 

/******************* CELL 6737 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6737 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6641]),
			.N(gen[6642]),
			.NE(gen[6643]),

			.O(gen[6736]),
			.E(gen[6738]),

			.SO(gen[6831]),
			.S(gen[6832]),
			.SE(gen[6833]),

			.SELF(gen[6737]),
			.cell_state(gen[6737])
		); 

/******************* CELL 6738 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6738 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6642]),
			.N(gen[6643]),
			.NE(gen[6644]),

			.O(gen[6737]),
			.E(gen[6739]),

			.SO(gen[6832]),
			.S(gen[6833]),
			.SE(gen[6834]),

			.SELF(gen[6738]),
			.cell_state(gen[6738])
		); 

/******************* CELL 6739 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6739 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6643]),
			.N(gen[6644]),
			.NE(gen[6645]),

			.O(gen[6738]),
			.E(gen[6740]),

			.SO(gen[6833]),
			.S(gen[6834]),
			.SE(gen[6835]),

			.SELF(gen[6739]),
			.cell_state(gen[6739])
		); 

/******************* CELL 6740 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6740 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6644]),
			.N(gen[6645]),
			.NE(gen[6646]),

			.O(gen[6739]),
			.E(gen[6741]),

			.SO(gen[6834]),
			.S(gen[6835]),
			.SE(gen[6836]),

			.SELF(gen[6740]),
			.cell_state(gen[6740])
		); 

/******************* CELL 6741 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6741 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6645]),
			.N(gen[6646]),
			.NE(gen[6647]),

			.O(gen[6740]),
			.E(gen[6742]),

			.SO(gen[6835]),
			.S(gen[6836]),
			.SE(gen[6837]),

			.SELF(gen[6741]),
			.cell_state(gen[6741])
		); 

/******************* CELL 6742 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6742 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6646]),
			.N(gen[6647]),
			.NE(gen[6648]),

			.O(gen[6741]),
			.E(gen[6743]),

			.SO(gen[6836]),
			.S(gen[6837]),
			.SE(gen[6838]),

			.SELF(gen[6742]),
			.cell_state(gen[6742])
		); 

/******************* CELL 6743 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6743 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6647]),
			.N(gen[6648]),
			.NE(gen[6649]),

			.O(gen[6742]),
			.E(gen[6744]),

			.SO(gen[6837]),
			.S(gen[6838]),
			.SE(gen[6839]),

			.SELF(gen[6743]),
			.cell_state(gen[6743])
		); 

/******************* CELL 6744 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6744 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6648]),
			.N(gen[6649]),
			.NE(gen[6648]),

			.O(gen[6743]),
			.E(gen[6743]),

			.SO(gen[6838]),
			.S(gen[6839]),
			.SE(gen[6838]),

			.SELF(gen[6744]),
			.cell_state(gen[6744])
		); 

/******************* CELL 6745 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6745 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6651]),
			.N(gen[6650]),
			.NE(gen[6651]),

			.O(gen[6746]),
			.E(gen[6746]),

			.SO(gen[6841]),
			.S(gen[6840]),
			.SE(gen[6841]),

			.SELF(gen[6745]),
			.cell_state(gen[6745])
		); 

/******************* CELL 6746 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6746 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6650]),
			.N(gen[6651]),
			.NE(gen[6652]),

			.O(gen[6745]),
			.E(gen[6747]),

			.SO(gen[6840]),
			.S(gen[6841]),
			.SE(gen[6842]),

			.SELF(gen[6746]),
			.cell_state(gen[6746])
		); 

/******************* CELL 6747 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6747 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6651]),
			.N(gen[6652]),
			.NE(gen[6653]),

			.O(gen[6746]),
			.E(gen[6748]),

			.SO(gen[6841]),
			.S(gen[6842]),
			.SE(gen[6843]),

			.SELF(gen[6747]),
			.cell_state(gen[6747])
		); 

/******************* CELL 6748 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6748 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6652]),
			.N(gen[6653]),
			.NE(gen[6654]),

			.O(gen[6747]),
			.E(gen[6749]),

			.SO(gen[6842]),
			.S(gen[6843]),
			.SE(gen[6844]),

			.SELF(gen[6748]),
			.cell_state(gen[6748])
		); 

/******************* CELL 6749 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6749 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6653]),
			.N(gen[6654]),
			.NE(gen[6655]),

			.O(gen[6748]),
			.E(gen[6750]),

			.SO(gen[6843]),
			.S(gen[6844]),
			.SE(gen[6845]),

			.SELF(gen[6749]),
			.cell_state(gen[6749])
		); 

/******************* CELL 6750 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6750 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6654]),
			.N(gen[6655]),
			.NE(gen[6656]),

			.O(gen[6749]),
			.E(gen[6751]),

			.SO(gen[6844]),
			.S(gen[6845]),
			.SE(gen[6846]),

			.SELF(gen[6750]),
			.cell_state(gen[6750])
		); 

/******************* CELL 6751 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6751 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6655]),
			.N(gen[6656]),
			.NE(gen[6657]),

			.O(gen[6750]),
			.E(gen[6752]),

			.SO(gen[6845]),
			.S(gen[6846]),
			.SE(gen[6847]),

			.SELF(gen[6751]),
			.cell_state(gen[6751])
		); 

/******************* CELL 6752 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6752 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6656]),
			.N(gen[6657]),
			.NE(gen[6658]),

			.O(gen[6751]),
			.E(gen[6753]),

			.SO(gen[6846]),
			.S(gen[6847]),
			.SE(gen[6848]),

			.SELF(gen[6752]),
			.cell_state(gen[6752])
		); 

/******************* CELL 6753 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6753 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6657]),
			.N(gen[6658]),
			.NE(gen[6659]),

			.O(gen[6752]),
			.E(gen[6754]),

			.SO(gen[6847]),
			.S(gen[6848]),
			.SE(gen[6849]),

			.SELF(gen[6753]),
			.cell_state(gen[6753])
		); 

/******************* CELL 6754 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6754 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6658]),
			.N(gen[6659]),
			.NE(gen[6660]),

			.O(gen[6753]),
			.E(gen[6755]),

			.SO(gen[6848]),
			.S(gen[6849]),
			.SE(gen[6850]),

			.SELF(gen[6754]),
			.cell_state(gen[6754])
		); 

/******************* CELL 6755 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6755 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6659]),
			.N(gen[6660]),
			.NE(gen[6661]),

			.O(gen[6754]),
			.E(gen[6756]),

			.SO(gen[6849]),
			.S(gen[6850]),
			.SE(gen[6851]),

			.SELF(gen[6755]),
			.cell_state(gen[6755])
		); 

/******************* CELL 6756 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6756 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6660]),
			.N(gen[6661]),
			.NE(gen[6662]),

			.O(gen[6755]),
			.E(gen[6757]),

			.SO(gen[6850]),
			.S(gen[6851]),
			.SE(gen[6852]),

			.SELF(gen[6756]),
			.cell_state(gen[6756])
		); 

/******************* CELL 6757 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6757 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6661]),
			.N(gen[6662]),
			.NE(gen[6663]),

			.O(gen[6756]),
			.E(gen[6758]),

			.SO(gen[6851]),
			.S(gen[6852]),
			.SE(gen[6853]),

			.SELF(gen[6757]),
			.cell_state(gen[6757])
		); 

/******************* CELL 6758 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6758 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6662]),
			.N(gen[6663]),
			.NE(gen[6664]),

			.O(gen[6757]),
			.E(gen[6759]),

			.SO(gen[6852]),
			.S(gen[6853]),
			.SE(gen[6854]),

			.SELF(gen[6758]),
			.cell_state(gen[6758])
		); 

/******************* CELL 6759 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6759 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6663]),
			.N(gen[6664]),
			.NE(gen[6665]),

			.O(gen[6758]),
			.E(gen[6760]),

			.SO(gen[6853]),
			.S(gen[6854]),
			.SE(gen[6855]),

			.SELF(gen[6759]),
			.cell_state(gen[6759])
		); 

/******************* CELL 6760 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6760 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6664]),
			.N(gen[6665]),
			.NE(gen[6666]),

			.O(gen[6759]),
			.E(gen[6761]),

			.SO(gen[6854]),
			.S(gen[6855]),
			.SE(gen[6856]),

			.SELF(gen[6760]),
			.cell_state(gen[6760])
		); 

/******************* CELL 6761 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6761 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6665]),
			.N(gen[6666]),
			.NE(gen[6667]),

			.O(gen[6760]),
			.E(gen[6762]),

			.SO(gen[6855]),
			.S(gen[6856]),
			.SE(gen[6857]),

			.SELF(gen[6761]),
			.cell_state(gen[6761])
		); 

/******************* CELL 6762 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6762 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6666]),
			.N(gen[6667]),
			.NE(gen[6668]),

			.O(gen[6761]),
			.E(gen[6763]),

			.SO(gen[6856]),
			.S(gen[6857]),
			.SE(gen[6858]),

			.SELF(gen[6762]),
			.cell_state(gen[6762])
		); 

/******************* CELL 6763 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6763 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6667]),
			.N(gen[6668]),
			.NE(gen[6669]),

			.O(gen[6762]),
			.E(gen[6764]),

			.SO(gen[6857]),
			.S(gen[6858]),
			.SE(gen[6859]),

			.SELF(gen[6763]),
			.cell_state(gen[6763])
		); 

/******************* CELL 6764 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6764 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6668]),
			.N(gen[6669]),
			.NE(gen[6670]),

			.O(gen[6763]),
			.E(gen[6765]),

			.SO(gen[6858]),
			.S(gen[6859]),
			.SE(gen[6860]),

			.SELF(gen[6764]),
			.cell_state(gen[6764])
		); 

/******************* CELL 6765 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6765 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6669]),
			.N(gen[6670]),
			.NE(gen[6671]),

			.O(gen[6764]),
			.E(gen[6766]),

			.SO(gen[6859]),
			.S(gen[6860]),
			.SE(gen[6861]),

			.SELF(gen[6765]),
			.cell_state(gen[6765])
		); 

/******************* CELL 6766 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6766 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6670]),
			.N(gen[6671]),
			.NE(gen[6672]),

			.O(gen[6765]),
			.E(gen[6767]),

			.SO(gen[6860]),
			.S(gen[6861]),
			.SE(gen[6862]),

			.SELF(gen[6766]),
			.cell_state(gen[6766])
		); 

/******************* CELL 6767 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6767 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6671]),
			.N(gen[6672]),
			.NE(gen[6673]),

			.O(gen[6766]),
			.E(gen[6768]),

			.SO(gen[6861]),
			.S(gen[6862]),
			.SE(gen[6863]),

			.SELF(gen[6767]),
			.cell_state(gen[6767])
		); 

/******************* CELL 6768 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6768 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6672]),
			.N(gen[6673]),
			.NE(gen[6674]),

			.O(gen[6767]),
			.E(gen[6769]),

			.SO(gen[6862]),
			.S(gen[6863]),
			.SE(gen[6864]),

			.SELF(gen[6768]),
			.cell_state(gen[6768])
		); 

/******************* CELL 6769 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6769 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6673]),
			.N(gen[6674]),
			.NE(gen[6675]),

			.O(gen[6768]),
			.E(gen[6770]),

			.SO(gen[6863]),
			.S(gen[6864]),
			.SE(gen[6865]),

			.SELF(gen[6769]),
			.cell_state(gen[6769])
		); 

/******************* CELL 6770 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6770 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6674]),
			.N(gen[6675]),
			.NE(gen[6676]),

			.O(gen[6769]),
			.E(gen[6771]),

			.SO(gen[6864]),
			.S(gen[6865]),
			.SE(gen[6866]),

			.SELF(gen[6770]),
			.cell_state(gen[6770])
		); 

/******************* CELL 6771 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6771 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6675]),
			.N(gen[6676]),
			.NE(gen[6677]),

			.O(gen[6770]),
			.E(gen[6772]),

			.SO(gen[6865]),
			.S(gen[6866]),
			.SE(gen[6867]),

			.SELF(gen[6771]),
			.cell_state(gen[6771])
		); 

/******************* CELL 6772 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6772 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6676]),
			.N(gen[6677]),
			.NE(gen[6678]),

			.O(gen[6771]),
			.E(gen[6773]),

			.SO(gen[6866]),
			.S(gen[6867]),
			.SE(gen[6868]),

			.SELF(gen[6772]),
			.cell_state(gen[6772])
		); 

/******************* CELL 6773 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6773 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6677]),
			.N(gen[6678]),
			.NE(gen[6679]),

			.O(gen[6772]),
			.E(gen[6774]),

			.SO(gen[6867]),
			.S(gen[6868]),
			.SE(gen[6869]),

			.SELF(gen[6773]),
			.cell_state(gen[6773])
		); 

/******************* CELL 6774 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6774 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6678]),
			.N(gen[6679]),
			.NE(gen[6680]),

			.O(gen[6773]),
			.E(gen[6775]),

			.SO(gen[6868]),
			.S(gen[6869]),
			.SE(gen[6870]),

			.SELF(gen[6774]),
			.cell_state(gen[6774])
		); 

/******************* CELL 6775 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6775 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6679]),
			.N(gen[6680]),
			.NE(gen[6681]),

			.O(gen[6774]),
			.E(gen[6776]),

			.SO(gen[6869]),
			.S(gen[6870]),
			.SE(gen[6871]),

			.SELF(gen[6775]),
			.cell_state(gen[6775])
		); 

/******************* CELL 6776 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6776 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6680]),
			.N(gen[6681]),
			.NE(gen[6682]),

			.O(gen[6775]),
			.E(gen[6777]),

			.SO(gen[6870]),
			.S(gen[6871]),
			.SE(gen[6872]),

			.SELF(gen[6776]),
			.cell_state(gen[6776])
		); 

/******************* CELL 6777 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6777 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6681]),
			.N(gen[6682]),
			.NE(gen[6683]),

			.O(gen[6776]),
			.E(gen[6778]),

			.SO(gen[6871]),
			.S(gen[6872]),
			.SE(gen[6873]),

			.SELF(gen[6777]),
			.cell_state(gen[6777])
		); 

/******************* CELL 6778 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6778 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6682]),
			.N(gen[6683]),
			.NE(gen[6684]),

			.O(gen[6777]),
			.E(gen[6779]),

			.SO(gen[6872]),
			.S(gen[6873]),
			.SE(gen[6874]),

			.SELF(gen[6778]),
			.cell_state(gen[6778])
		); 

/******************* CELL 6779 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6779 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6683]),
			.N(gen[6684]),
			.NE(gen[6685]),

			.O(gen[6778]),
			.E(gen[6780]),

			.SO(gen[6873]),
			.S(gen[6874]),
			.SE(gen[6875]),

			.SELF(gen[6779]),
			.cell_state(gen[6779])
		); 

/******************* CELL 6780 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6780 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6684]),
			.N(gen[6685]),
			.NE(gen[6686]),

			.O(gen[6779]),
			.E(gen[6781]),

			.SO(gen[6874]),
			.S(gen[6875]),
			.SE(gen[6876]),

			.SELF(gen[6780]),
			.cell_state(gen[6780])
		); 

/******************* CELL 6781 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6781 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6685]),
			.N(gen[6686]),
			.NE(gen[6687]),

			.O(gen[6780]),
			.E(gen[6782]),

			.SO(gen[6875]),
			.S(gen[6876]),
			.SE(gen[6877]),

			.SELF(gen[6781]),
			.cell_state(gen[6781])
		); 

/******************* CELL 6782 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6782 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6686]),
			.N(gen[6687]),
			.NE(gen[6688]),

			.O(gen[6781]),
			.E(gen[6783]),

			.SO(gen[6876]),
			.S(gen[6877]),
			.SE(gen[6878]),

			.SELF(gen[6782]),
			.cell_state(gen[6782])
		); 

/******************* CELL 6783 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6783 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6687]),
			.N(gen[6688]),
			.NE(gen[6689]),

			.O(gen[6782]),
			.E(gen[6784]),

			.SO(gen[6877]),
			.S(gen[6878]),
			.SE(gen[6879]),

			.SELF(gen[6783]),
			.cell_state(gen[6783])
		); 

/******************* CELL 6784 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6784 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6688]),
			.N(gen[6689]),
			.NE(gen[6690]),

			.O(gen[6783]),
			.E(gen[6785]),

			.SO(gen[6878]),
			.S(gen[6879]),
			.SE(gen[6880]),

			.SELF(gen[6784]),
			.cell_state(gen[6784])
		); 

/******************* CELL 6785 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6785 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6689]),
			.N(gen[6690]),
			.NE(gen[6691]),

			.O(gen[6784]),
			.E(gen[6786]),

			.SO(gen[6879]),
			.S(gen[6880]),
			.SE(gen[6881]),

			.SELF(gen[6785]),
			.cell_state(gen[6785])
		); 

/******************* CELL 6786 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6786 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6690]),
			.N(gen[6691]),
			.NE(gen[6692]),

			.O(gen[6785]),
			.E(gen[6787]),

			.SO(gen[6880]),
			.S(gen[6881]),
			.SE(gen[6882]),

			.SELF(gen[6786]),
			.cell_state(gen[6786])
		); 

/******************* CELL 6787 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6787 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6691]),
			.N(gen[6692]),
			.NE(gen[6693]),

			.O(gen[6786]),
			.E(gen[6788]),

			.SO(gen[6881]),
			.S(gen[6882]),
			.SE(gen[6883]),

			.SELF(gen[6787]),
			.cell_state(gen[6787])
		); 

/******************* CELL 6788 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6788 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6692]),
			.N(gen[6693]),
			.NE(gen[6694]),

			.O(gen[6787]),
			.E(gen[6789]),

			.SO(gen[6882]),
			.S(gen[6883]),
			.SE(gen[6884]),

			.SELF(gen[6788]),
			.cell_state(gen[6788])
		); 

/******************* CELL 6789 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6789 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6693]),
			.N(gen[6694]),
			.NE(gen[6695]),

			.O(gen[6788]),
			.E(gen[6790]),

			.SO(gen[6883]),
			.S(gen[6884]),
			.SE(gen[6885]),

			.SELF(gen[6789]),
			.cell_state(gen[6789])
		); 

/******************* CELL 6790 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6790 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6694]),
			.N(gen[6695]),
			.NE(gen[6696]),

			.O(gen[6789]),
			.E(gen[6791]),

			.SO(gen[6884]),
			.S(gen[6885]),
			.SE(gen[6886]),

			.SELF(gen[6790]),
			.cell_state(gen[6790])
		); 

/******************* CELL 6791 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6791 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6695]),
			.N(gen[6696]),
			.NE(gen[6697]),

			.O(gen[6790]),
			.E(gen[6792]),

			.SO(gen[6885]),
			.S(gen[6886]),
			.SE(gen[6887]),

			.SELF(gen[6791]),
			.cell_state(gen[6791])
		); 

/******************* CELL 6792 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6792 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6696]),
			.N(gen[6697]),
			.NE(gen[6698]),

			.O(gen[6791]),
			.E(gen[6793]),

			.SO(gen[6886]),
			.S(gen[6887]),
			.SE(gen[6888]),

			.SELF(gen[6792]),
			.cell_state(gen[6792])
		); 

/******************* CELL 6793 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6793 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6697]),
			.N(gen[6698]),
			.NE(gen[6699]),

			.O(gen[6792]),
			.E(gen[6794]),

			.SO(gen[6887]),
			.S(gen[6888]),
			.SE(gen[6889]),

			.SELF(gen[6793]),
			.cell_state(gen[6793])
		); 

/******************* CELL 6794 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6794 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6698]),
			.N(gen[6699]),
			.NE(gen[6700]),

			.O(gen[6793]),
			.E(gen[6795]),

			.SO(gen[6888]),
			.S(gen[6889]),
			.SE(gen[6890]),

			.SELF(gen[6794]),
			.cell_state(gen[6794])
		); 

/******************* CELL 6795 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6795 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6699]),
			.N(gen[6700]),
			.NE(gen[6701]),

			.O(gen[6794]),
			.E(gen[6796]),

			.SO(gen[6889]),
			.S(gen[6890]),
			.SE(gen[6891]),

			.SELF(gen[6795]),
			.cell_state(gen[6795])
		); 

/******************* CELL 6796 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6796 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6700]),
			.N(gen[6701]),
			.NE(gen[6702]),

			.O(gen[6795]),
			.E(gen[6797]),

			.SO(gen[6890]),
			.S(gen[6891]),
			.SE(gen[6892]),

			.SELF(gen[6796]),
			.cell_state(gen[6796])
		); 

/******************* CELL 6797 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6797 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6701]),
			.N(gen[6702]),
			.NE(gen[6703]),

			.O(gen[6796]),
			.E(gen[6798]),

			.SO(gen[6891]),
			.S(gen[6892]),
			.SE(gen[6893]),

			.SELF(gen[6797]),
			.cell_state(gen[6797])
		); 

/******************* CELL 6798 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6798 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6702]),
			.N(gen[6703]),
			.NE(gen[6704]),

			.O(gen[6797]),
			.E(gen[6799]),

			.SO(gen[6892]),
			.S(gen[6893]),
			.SE(gen[6894]),

			.SELF(gen[6798]),
			.cell_state(gen[6798])
		); 

/******************* CELL 6799 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6799 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6703]),
			.N(gen[6704]),
			.NE(gen[6705]),

			.O(gen[6798]),
			.E(gen[6800]),

			.SO(gen[6893]),
			.S(gen[6894]),
			.SE(gen[6895]),

			.SELF(gen[6799]),
			.cell_state(gen[6799])
		); 

/******************* CELL 6800 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6800 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6704]),
			.N(gen[6705]),
			.NE(gen[6706]),

			.O(gen[6799]),
			.E(gen[6801]),

			.SO(gen[6894]),
			.S(gen[6895]),
			.SE(gen[6896]),

			.SELF(gen[6800]),
			.cell_state(gen[6800])
		); 

/******************* CELL 6801 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6801 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6705]),
			.N(gen[6706]),
			.NE(gen[6707]),

			.O(gen[6800]),
			.E(gen[6802]),

			.SO(gen[6895]),
			.S(gen[6896]),
			.SE(gen[6897]),

			.SELF(gen[6801]),
			.cell_state(gen[6801])
		); 

/******************* CELL 6802 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6802 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6706]),
			.N(gen[6707]),
			.NE(gen[6708]),

			.O(gen[6801]),
			.E(gen[6803]),

			.SO(gen[6896]),
			.S(gen[6897]),
			.SE(gen[6898]),

			.SELF(gen[6802]),
			.cell_state(gen[6802])
		); 

/******************* CELL 6803 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6803 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6707]),
			.N(gen[6708]),
			.NE(gen[6709]),

			.O(gen[6802]),
			.E(gen[6804]),

			.SO(gen[6897]),
			.S(gen[6898]),
			.SE(gen[6899]),

			.SELF(gen[6803]),
			.cell_state(gen[6803])
		); 

/******************* CELL 6804 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6804 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6708]),
			.N(gen[6709]),
			.NE(gen[6710]),

			.O(gen[6803]),
			.E(gen[6805]),

			.SO(gen[6898]),
			.S(gen[6899]),
			.SE(gen[6900]),

			.SELF(gen[6804]),
			.cell_state(gen[6804])
		); 

/******************* CELL 6805 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6805 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6709]),
			.N(gen[6710]),
			.NE(gen[6711]),

			.O(gen[6804]),
			.E(gen[6806]),

			.SO(gen[6899]),
			.S(gen[6900]),
			.SE(gen[6901]),

			.SELF(gen[6805]),
			.cell_state(gen[6805])
		); 

/******************* CELL 6806 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6806 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6710]),
			.N(gen[6711]),
			.NE(gen[6712]),

			.O(gen[6805]),
			.E(gen[6807]),

			.SO(gen[6900]),
			.S(gen[6901]),
			.SE(gen[6902]),

			.SELF(gen[6806]),
			.cell_state(gen[6806])
		); 

/******************* CELL 6807 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6807 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6711]),
			.N(gen[6712]),
			.NE(gen[6713]),

			.O(gen[6806]),
			.E(gen[6808]),

			.SO(gen[6901]),
			.S(gen[6902]),
			.SE(gen[6903]),

			.SELF(gen[6807]),
			.cell_state(gen[6807])
		); 

/******************* CELL 6808 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6808 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6712]),
			.N(gen[6713]),
			.NE(gen[6714]),

			.O(gen[6807]),
			.E(gen[6809]),

			.SO(gen[6902]),
			.S(gen[6903]),
			.SE(gen[6904]),

			.SELF(gen[6808]),
			.cell_state(gen[6808])
		); 

/******************* CELL 6809 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6809 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6713]),
			.N(gen[6714]),
			.NE(gen[6715]),

			.O(gen[6808]),
			.E(gen[6810]),

			.SO(gen[6903]),
			.S(gen[6904]),
			.SE(gen[6905]),

			.SELF(gen[6809]),
			.cell_state(gen[6809])
		); 

/******************* CELL 6810 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6810 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6714]),
			.N(gen[6715]),
			.NE(gen[6716]),

			.O(gen[6809]),
			.E(gen[6811]),

			.SO(gen[6904]),
			.S(gen[6905]),
			.SE(gen[6906]),

			.SELF(gen[6810]),
			.cell_state(gen[6810])
		); 

/******************* CELL 6811 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6811 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6715]),
			.N(gen[6716]),
			.NE(gen[6717]),

			.O(gen[6810]),
			.E(gen[6812]),

			.SO(gen[6905]),
			.S(gen[6906]),
			.SE(gen[6907]),

			.SELF(gen[6811]),
			.cell_state(gen[6811])
		); 

/******************* CELL 6812 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6812 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6716]),
			.N(gen[6717]),
			.NE(gen[6718]),

			.O(gen[6811]),
			.E(gen[6813]),

			.SO(gen[6906]),
			.S(gen[6907]),
			.SE(gen[6908]),

			.SELF(gen[6812]),
			.cell_state(gen[6812])
		); 

/******************* CELL 6813 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6813 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6717]),
			.N(gen[6718]),
			.NE(gen[6719]),

			.O(gen[6812]),
			.E(gen[6814]),

			.SO(gen[6907]),
			.S(gen[6908]),
			.SE(gen[6909]),

			.SELF(gen[6813]),
			.cell_state(gen[6813])
		); 

/******************* CELL 6814 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6814 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6718]),
			.N(gen[6719]),
			.NE(gen[6720]),

			.O(gen[6813]),
			.E(gen[6815]),

			.SO(gen[6908]),
			.S(gen[6909]),
			.SE(gen[6910]),

			.SELF(gen[6814]),
			.cell_state(gen[6814])
		); 

/******************* CELL 6815 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6815 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6719]),
			.N(gen[6720]),
			.NE(gen[6721]),

			.O(gen[6814]),
			.E(gen[6816]),

			.SO(gen[6909]),
			.S(gen[6910]),
			.SE(gen[6911]),

			.SELF(gen[6815]),
			.cell_state(gen[6815])
		); 

/******************* CELL 6816 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6816 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6720]),
			.N(gen[6721]),
			.NE(gen[6722]),

			.O(gen[6815]),
			.E(gen[6817]),

			.SO(gen[6910]),
			.S(gen[6911]),
			.SE(gen[6912]),

			.SELF(gen[6816]),
			.cell_state(gen[6816])
		); 

/******************* CELL 6817 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6817 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6721]),
			.N(gen[6722]),
			.NE(gen[6723]),

			.O(gen[6816]),
			.E(gen[6818]),

			.SO(gen[6911]),
			.S(gen[6912]),
			.SE(gen[6913]),

			.SELF(gen[6817]),
			.cell_state(gen[6817])
		); 

/******************* CELL 6818 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6818 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6722]),
			.N(gen[6723]),
			.NE(gen[6724]),

			.O(gen[6817]),
			.E(gen[6819]),

			.SO(gen[6912]),
			.S(gen[6913]),
			.SE(gen[6914]),

			.SELF(gen[6818]),
			.cell_state(gen[6818])
		); 

/******************* CELL 6819 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6819 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6723]),
			.N(gen[6724]),
			.NE(gen[6725]),

			.O(gen[6818]),
			.E(gen[6820]),

			.SO(gen[6913]),
			.S(gen[6914]),
			.SE(gen[6915]),

			.SELF(gen[6819]),
			.cell_state(gen[6819])
		); 

/******************* CELL 6820 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6820 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6724]),
			.N(gen[6725]),
			.NE(gen[6726]),

			.O(gen[6819]),
			.E(gen[6821]),

			.SO(gen[6914]),
			.S(gen[6915]),
			.SE(gen[6916]),

			.SELF(gen[6820]),
			.cell_state(gen[6820])
		); 

/******************* CELL 6821 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6821 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6725]),
			.N(gen[6726]),
			.NE(gen[6727]),

			.O(gen[6820]),
			.E(gen[6822]),

			.SO(gen[6915]),
			.S(gen[6916]),
			.SE(gen[6917]),

			.SELF(gen[6821]),
			.cell_state(gen[6821])
		); 

/******************* CELL 6822 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6822 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6726]),
			.N(gen[6727]),
			.NE(gen[6728]),

			.O(gen[6821]),
			.E(gen[6823]),

			.SO(gen[6916]),
			.S(gen[6917]),
			.SE(gen[6918]),

			.SELF(gen[6822]),
			.cell_state(gen[6822])
		); 

/******************* CELL 6823 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6823 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6727]),
			.N(gen[6728]),
			.NE(gen[6729]),

			.O(gen[6822]),
			.E(gen[6824]),

			.SO(gen[6917]),
			.S(gen[6918]),
			.SE(gen[6919]),

			.SELF(gen[6823]),
			.cell_state(gen[6823])
		); 

/******************* CELL 6824 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6824 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6728]),
			.N(gen[6729]),
			.NE(gen[6730]),

			.O(gen[6823]),
			.E(gen[6825]),

			.SO(gen[6918]),
			.S(gen[6919]),
			.SE(gen[6920]),

			.SELF(gen[6824]),
			.cell_state(gen[6824])
		); 

/******************* CELL 6825 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6825 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6729]),
			.N(gen[6730]),
			.NE(gen[6731]),

			.O(gen[6824]),
			.E(gen[6826]),

			.SO(gen[6919]),
			.S(gen[6920]),
			.SE(gen[6921]),

			.SELF(gen[6825]),
			.cell_state(gen[6825])
		); 

/******************* CELL 6826 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6826 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6730]),
			.N(gen[6731]),
			.NE(gen[6732]),

			.O(gen[6825]),
			.E(gen[6827]),

			.SO(gen[6920]),
			.S(gen[6921]),
			.SE(gen[6922]),

			.SELF(gen[6826]),
			.cell_state(gen[6826])
		); 

/******************* CELL 6827 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6827 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6731]),
			.N(gen[6732]),
			.NE(gen[6733]),

			.O(gen[6826]),
			.E(gen[6828]),

			.SO(gen[6921]),
			.S(gen[6922]),
			.SE(gen[6923]),

			.SELF(gen[6827]),
			.cell_state(gen[6827])
		); 

/******************* CELL 6828 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6828 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6732]),
			.N(gen[6733]),
			.NE(gen[6734]),

			.O(gen[6827]),
			.E(gen[6829]),

			.SO(gen[6922]),
			.S(gen[6923]),
			.SE(gen[6924]),

			.SELF(gen[6828]),
			.cell_state(gen[6828])
		); 

/******************* CELL 6829 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6829 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6733]),
			.N(gen[6734]),
			.NE(gen[6735]),

			.O(gen[6828]),
			.E(gen[6830]),

			.SO(gen[6923]),
			.S(gen[6924]),
			.SE(gen[6925]),

			.SELF(gen[6829]),
			.cell_state(gen[6829])
		); 

/******************* CELL 6830 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6830 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6734]),
			.N(gen[6735]),
			.NE(gen[6736]),

			.O(gen[6829]),
			.E(gen[6831]),

			.SO(gen[6924]),
			.S(gen[6925]),
			.SE(gen[6926]),

			.SELF(gen[6830]),
			.cell_state(gen[6830])
		); 

/******************* CELL 6831 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6831 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6735]),
			.N(gen[6736]),
			.NE(gen[6737]),

			.O(gen[6830]),
			.E(gen[6832]),

			.SO(gen[6925]),
			.S(gen[6926]),
			.SE(gen[6927]),

			.SELF(gen[6831]),
			.cell_state(gen[6831])
		); 

/******************* CELL 6832 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6832 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6736]),
			.N(gen[6737]),
			.NE(gen[6738]),

			.O(gen[6831]),
			.E(gen[6833]),

			.SO(gen[6926]),
			.S(gen[6927]),
			.SE(gen[6928]),

			.SELF(gen[6832]),
			.cell_state(gen[6832])
		); 

/******************* CELL 6833 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6833 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6737]),
			.N(gen[6738]),
			.NE(gen[6739]),

			.O(gen[6832]),
			.E(gen[6834]),

			.SO(gen[6927]),
			.S(gen[6928]),
			.SE(gen[6929]),

			.SELF(gen[6833]),
			.cell_state(gen[6833])
		); 

/******************* CELL 6834 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6834 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6738]),
			.N(gen[6739]),
			.NE(gen[6740]),

			.O(gen[6833]),
			.E(gen[6835]),

			.SO(gen[6928]),
			.S(gen[6929]),
			.SE(gen[6930]),

			.SELF(gen[6834]),
			.cell_state(gen[6834])
		); 

/******************* CELL 6835 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6835 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6739]),
			.N(gen[6740]),
			.NE(gen[6741]),

			.O(gen[6834]),
			.E(gen[6836]),

			.SO(gen[6929]),
			.S(gen[6930]),
			.SE(gen[6931]),

			.SELF(gen[6835]),
			.cell_state(gen[6835])
		); 

/******************* CELL 6836 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6836 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6740]),
			.N(gen[6741]),
			.NE(gen[6742]),

			.O(gen[6835]),
			.E(gen[6837]),

			.SO(gen[6930]),
			.S(gen[6931]),
			.SE(gen[6932]),

			.SELF(gen[6836]),
			.cell_state(gen[6836])
		); 

/******************* CELL 6837 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6837 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6741]),
			.N(gen[6742]),
			.NE(gen[6743]),

			.O(gen[6836]),
			.E(gen[6838]),

			.SO(gen[6931]),
			.S(gen[6932]),
			.SE(gen[6933]),

			.SELF(gen[6837]),
			.cell_state(gen[6837])
		); 

/******************* CELL 6838 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6838 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6742]),
			.N(gen[6743]),
			.NE(gen[6744]),

			.O(gen[6837]),
			.E(gen[6839]),

			.SO(gen[6932]),
			.S(gen[6933]),
			.SE(gen[6934]),

			.SELF(gen[6838]),
			.cell_state(gen[6838])
		); 

/******************* CELL 6839 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6839 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6743]),
			.N(gen[6744]),
			.NE(gen[6743]),

			.O(gen[6838]),
			.E(gen[6838]),

			.SO(gen[6933]),
			.S(gen[6934]),
			.SE(gen[6933]),

			.SELF(gen[6839]),
			.cell_state(gen[6839])
		); 

/******************* CELL 6840 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6840 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6746]),
			.N(gen[6745]),
			.NE(gen[6746]),

			.O(gen[6841]),
			.E(gen[6841]),

			.SO(gen[6936]),
			.S(gen[6935]),
			.SE(gen[6936]),

			.SELF(gen[6840]),
			.cell_state(gen[6840])
		); 

/******************* CELL 6841 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6841 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6745]),
			.N(gen[6746]),
			.NE(gen[6747]),

			.O(gen[6840]),
			.E(gen[6842]),

			.SO(gen[6935]),
			.S(gen[6936]),
			.SE(gen[6937]),

			.SELF(gen[6841]),
			.cell_state(gen[6841])
		); 

/******************* CELL 6842 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6842 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6746]),
			.N(gen[6747]),
			.NE(gen[6748]),

			.O(gen[6841]),
			.E(gen[6843]),

			.SO(gen[6936]),
			.S(gen[6937]),
			.SE(gen[6938]),

			.SELF(gen[6842]),
			.cell_state(gen[6842])
		); 

/******************* CELL 6843 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6843 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6747]),
			.N(gen[6748]),
			.NE(gen[6749]),

			.O(gen[6842]),
			.E(gen[6844]),

			.SO(gen[6937]),
			.S(gen[6938]),
			.SE(gen[6939]),

			.SELF(gen[6843]),
			.cell_state(gen[6843])
		); 

/******************* CELL 6844 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6844 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6748]),
			.N(gen[6749]),
			.NE(gen[6750]),

			.O(gen[6843]),
			.E(gen[6845]),

			.SO(gen[6938]),
			.S(gen[6939]),
			.SE(gen[6940]),

			.SELF(gen[6844]),
			.cell_state(gen[6844])
		); 

/******************* CELL 6845 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6845 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6749]),
			.N(gen[6750]),
			.NE(gen[6751]),

			.O(gen[6844]),
			.E(gen[6846]),

			.SO(gen[6939]),
			.S(gen[6940]),
			.SE(gen[6941]),

			.SELF(gen[6845]),
			.cell_state(gen[6845])
		); 

/******************* CELL 6846 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6846 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6750]),
			.N(gen[6751]),
			.NE(gen[6752]),

			.O(gen[6845]),
			.E(gen[6847]),

			.SO(gen[6940]),
			.S(gen[6941]),
			.SE(gen[6942]),

			.SELF(gen[6846]),
			.cell_state(gen[6846])
		); 

/******************* CELL 6847 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6847 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6751]),
			.N(gen[6752]),
			.NE(gen[6753]),

			.O(gen[6846]),
			.E(gen[6848]),

			.SO(gen[6941]),
			.S(gen[6942]),
			.SE(gen[6943]),

			.SELF(gen[6847]),
			.cell_state(gen[6847])
		); 

/******************* CELL 6848 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6848 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6752]),
			.N(gen[6753]),
			.NE(gen[6754]),

			.O(gen[6847]),
			.E(gen[6849]),

			.SO(gen[6942]),
			.S(gen[6943]),
			.SE(gen[6944]),

			.SELF(gen[6848]),
			.cell_state(gen[6848])
		); 

/******************* CELL 6849 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6849 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6753]),
			.N(gen[6754]),
			.NE(gen[6755]),

			.O(gen[6848]),
			.E(gen[6850]),

			.SO(gen[6943]),
			.S(gen[6944]),
			.SE(gen[6945]),

			.SELF(gen[6849]),
			.cell_state(gen[6849])
		); 

/******************* CELL 6850 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6850 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6754]),
			.N(gen[6755]),
			.NE(gen[6756]),

			.O(gen[6849]),
			.E(gen[6851]),

			.SO(gen[6944]),
			.S(gen[6945]),
			.SE(gen[6946]),

			.SELF(gen[6850]),
			.cell_state(gen[6850])
		); 

/******************* CELL 6851 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6851 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6755]),
			.N(gen[6756]),
			.NE(gen[6757]),

			.O(gen[6850]),
			.E(gen[6852]),

			.SO(gen[6945]),
			.S(gen[6946]),
			.SE(gen[6947]),

			.SELF(gen[6851]),
			.cell_state(gen[6851])
		); 

/******************* CELL 6852 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6852 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6756]),
			.N(gen[6757]),
			.NE(gen[6758]),

			.O(gen[6851]),
			.E(gen[6853]),

			.SO(gen[6946]),
			.S(gen[6947]),
			.SE(gen[6948]),

			.SELF(gen[6852]),
			.cell_state(gen[6852])
		); 

/******************* CELL 6853 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6853 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6757]),
			.N(gen[6758]),
			.NE(gen[6759]),

			.O(gen[6852]),
			.E(gen[6854]),

			.SO(gen[6947]),
			.S(gen[6948]),
			.SE(gen[6949]),

			.SELF(gen[6853]),
			.cell_state(gen[6853])
		); 

/******************* CELL 6854 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6854 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6758]),
			.N(gen[6759]),
			.NE(gen[6760]),

			.O(gen[6853]),
			.E(gen[6855]),

			.SO(gen[6948]),
			.S(gen[6949]),
			.SE(gen[6950]),

			.SELF(gen[6854]),
			.cell_state(gen[6854])
		); 

/******************* CELL 6855 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6855 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6759]),
			.N(gen[6760]),
			.NE(gen[6761]),

			.O(gen[6854]),
			.E(gen[6856]),

			.SO(gen[6949]),
			.S(gen[6950]),
			.SE(gen[6951]),

			.SELF(gen[6855]),
			.cell_state(gen[6855])
		); 

/******************* CELL 6856 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6856 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6760]),
			.N(gen[6761]),
			.NE(gen[6762]),

			.O(gen[6855]),
			.E(gen[6857]),

			.SO(gen[6950]),
			.S(gen[6951]),
			.SE(gen[6952]),

			.SELF(gen[6856]),
			.cell_state(gen[6856])
		); 

/******************* CELL 6857 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6857 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6761]),
			.N(gen[6762]),
			.NE(gen[6763]),

			.O(gen[6856]),
			.E(gen[6858]),

			.SO(gen[6951]),
			.S(gen[6952]),
			.SE(gen[6953]),

			.SELF(gen[6857]),
			.cell_state(gen[6857])
		); 

/******************* CELL 6858 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6858 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6762]),
			.N(gen[6763]),
			.NE(gen[6764]),

			.O(gen[6857]),
			.E(gen[6859]),

			.SO(gen[6952]),
			.S(gen[6953]),
			.SE(gen[6954]),

			.SELF(gen[6858]),
			.cell_state(gen[6858])
		); 

/******************* CELL 6859 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6859 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6763]),
			.N(gen[6764]),
			.NE(gen[6765]),

			.O(gen[6858]),
			.E(gen[6860]),

			.SO(gen[6953]),
			.S(gen[6954]),
			.SE(gen[6955]),

			.SELF(gen[6859]),
			.cell_state(gen[6859])
		); 

/******************* CELL 6860 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6860 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6764]),
			.N(gen[6765]),
			.NE(gen[6766]),

			.O(gen[6859]),
			.E(gen[6861]),

			.SO(gen[6954]),
			.S(gen[6955]),
			.SE(gen[6956]),

			.SELF(gen[6860]),
			.cell_state(gen[6860])
		); 

/******************* CELL 6861 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6861 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6765]),
			.N(gen[6766]),
			.NE(gen[6767]),

			.O(gen[6860]),
			.E(gen[6862]),

			.SO(gen[6955]),
			.S(gen[6956]),
			.SE(gen[6957]),

			.SELF(gen[6861]),
			.cell_state(gen[6861])
		); 

/******************* CELL 6862 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6862 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6766]),
			.N(gen[6767]),
			.NE(gen[6768]),

			.O(gen[6861]),
			.E(gen[6863]),

			.SO(gen[6956]),
			.S(gen[6957]),
			.SE(gen[6958]),

			.SELF(gen[6862]),
			.cell_state(gen[6862])
		); 

/******************* CELL 6863 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6863 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6767]),
			.N(gen[6768]),
			.NE(gen[6769]),

			.O(gen[6862]),
			.E(gen[6864]),

			.SO(gen[6957]),
			.S(gen[6958]),
			.SE(gen[6959]),

			.SELF(gen[6863]),
			.cell_state(gen[6863])
		); 

/******************* CELL 6864 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6864 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6768]),
			.N(gen[6769]),
			.NE(gen[6770]),

			.O(gen[6863]),
			.E(gen[6865]),

			.SO(gen[6958]),
			.S(gen[6959]),
			.SE(gen[6960]),

			.SELF(gen[6864]),
			.cell_state(gen[6864])
		); 

/******************* CELL 6865 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6865 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6769]),
			.N(gen[6770]),
			.NE(gen[6771]),

			.O(gen[6864]),
			.E(gen[6866]),

			.SO(gen[6959]),
			.S(gen[6960]),
			.SE(gen[6961]),

			.SELF(gen[6865]),
			.cell_state(gen[6865])
		); 

/******************* CELL 6866 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6866 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6770]),
			.N(gen[6771]),
			.NE(gen[6772]),

			.O(gen[6865]),
			.E(gen[6867]),

			.SO(gen[6960]),
			.S(gen[6961]),
			.SE(gen[6962]),

			.SELF(gen[6866]),
			.cell_state(gen[6866])
		); 

/******************* CELL 6867 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6867 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6771]),
			.N(gen[6772]),
			.NE(gen[6773]),

			.O(gen[6866]),
			.E(gen[6868]),

			.SO(gen[6961]),
			.S(gen[6962]),
			.SE(gen[6963]),

			.SELF(gen[6867]),
			.cell_state(gen[6867])
		); 

/******************* CELL 6868 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6868 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6772]),
			.N(gen[6773]),
			.NE(gen[6774]),

			.O(gen[6867]),
			.E(gen[6869]),

			.SO(gen[6962]),
			.S(gen[6963]),
			.SE(gen[6964]),

			.SELF(gen[6868]),
			.cell_state(gen[6868])
		); 

/******************* CELL 6869 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6869 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6773]),
			.N(gen[6774]),
			.NE(gen[6775]),

			.O(gen[6868]),
			.E(gen[6870]),

			.SO(gen[6963]),
			.S(gen[6964]),
			.SE(gen[6965]),

			.SELF(gen[6869]),
			.cell_state(gen[6869])
		); 

/******************* CELL 6870 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6870 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6774]),
			.N(gen[6775]),
			.NE(gen[6776]),

			.O(gen[6869]),
			.E(gen[6871]),

			.SO(gen[6964]),
			.S(gen[6965]),
			.SE(gen[6966]),

			.SELF(gen[6870]),
			.cell_state(gen[6870])
		); 

/******************* CELL 6871 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6871 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6775]),
			.N(gen[6776]),
			.NE(gen[6777]),

			.O(gen[6870]),
			.E(gen[6872]),

			.SO(gen[6965]),
			.S(gen[6966]),
			.SE(gen[6967]),

			.SELF(gen[6871]),
			.cell_state(gen[6871])
		); 

/******************* CELL 6872 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6872 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6776]),
			.N(gen[6777]),
			.NE(gen[6778]),

			.O(gen[6871]),
			.E(gen[6873]),

			.SO(gen[6966]),
			.S(gen[6967]),
			.SE(gen[6968]),

			.SELF(gen[6872]),
			.cell_state(gen[6872])
		); 

/******************* CELL 6873 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6873 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6777]),
			.N(gen[6778]),
			.NE(gen[6779]),

			.O(gen[6872]),
			.E(gen[6874]),

			.SO(gen[6967]),
			.S(gen[6968]),
			.SE(gen[6969]),

			.SELF(gen[6873]),
			.cell_state(gen[6873])
		); 

/******************* CELL 6874 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6874 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6778]),
			.N(gen[6779]),
			.NE(gen[6780]),

			.O(gen[6873]),
			.E(gen[6875]),

			.SO(gen[6968]),
			.S(gen[6969]),
			.SE(gen[6970]),

			.SELF(gen[6874]),
			.cell_state(gen[6874])
		); 

/******************* CELL 6875 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6875 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6779]),
			.N(gen[6780]),
			.NE(gen[6781]),

			.O(gen[6874]),
			.E(gen[6876]),

			.SO(gen[6969]),
			.S(gen[6970]),
			.SE(gen[6971]),

			.SELF(gen[6875]),
			.cell_state(gen[6875])
		); 

/******************* CELL 6876 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6876 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6780]),
			.N(gen[6781]),
			.NE(gen[6782]),

			.O(gen[6875]),
			.E(gen[6877]),

			.SO(gen[6970]),
			.S(gen[6971]),
			.SE(gen[6972]),

			.SELF(gen[6876]),
			.cell_state(gen[6876])
		); 

/******************* CELL 6877 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6877 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6781]),
			.N(gen[6782]),
			.NE(gen[6783]),

			.O(gen[6876]),
			.E(gen[6878]),

			.SO(gen[6971]),
			.S(gen[6972]),
			.SE(gen[6973]),

			.SELF(gen[6877]),
			.cell_state(gen[6877])
		); 

/******************* CELL 6878 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6878 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6782]),
			.N(gen[6783]),
			.NE(gen[6784]),

			.O(gen[6877]),
			.E(gen[6879]),

			.SO(gen[6972]),
			.S(gen[6973]),
			.SE(gen[6974]),

			.SELF(gen[6878]),
			.cell_state(gen[6878])
		); 

/******************* CELL 6879 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6879 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6783]),
			.N(gen[6784]),
			.NE(gen[6785]),

			.O(gen[6878]),
			.E(gen[6880]),

			.SO(gen[6973]),
			.S(gen[6974]),
			.SE(gen[6975]),

			.SELF(gen[6879]),
			.cell_state(gen[6879])
		); 

/******************* CELL 6880 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6880 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6784]),
			.N(gen[6785]),
			.NE(gen[6786]),

			.O(gen[6879]),
			.E(gen[6881]),

			.SO(gen[6974]),
			.S(gen[6975]),
			.SE(gen[6976]),

			.SELF(gen[6880]),
			.cell_state(gen[6880])
		); 

/******************* CELL 6881 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6881 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6785]),
			.N(gen[6786]),
			.NE(gen[6787]),

			.O(gen[6880]),
			.E(gen[6882]),

			.SO(gen[6975]),
			.S(gen[6976]),
			.SE(gen[6977]),

			.SELF(gen[6881]),
			.cell_state(gen[6881])
		); 

/******************* CELL 6882 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6882 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6786]),
			.N(gen[6787]),
			.NE(gen[6788]),

			.O(gen[6881]),
			.E(gen[6883]),

			.SO(gen[6976]),
			.S(gen[6977]),
			.SE(gen[6978]),

			.SELF(gen[6882]),
			.cell_state(gen[6882])
		); 

/******************* CELL 6883 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6883 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6787]),
			.N(gen[6788]),
			.NE(gen[6789]),

			.O(gen[6882]),
			.E(gen[6884]),

			.SO(gen[6977]),
			.S(gen[6978]),
			.SE(gen[6979]),

			.SELF(gen[6883]),
			.cell_state(gen[6883])
		); 

/******************* CELL 6884 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6884 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6788]),
			.N(gen[6789]),
			.NE(gen[6790]),

			.O(gen[6883]),
			.E(gen[6885]),

			.SO(gen[6978]),
			.S(gen[6979]),
			.SE(gen[6980]),

			.SELF(gen[6884]),
			.cell_state(gen[6884])
		); 

/******************* CELL 6885 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6885 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6789]),
			.N(gen[6790]),
			.NE(gen[6791]),

			.O(gen[6884]),
			.E(gen[6886]),

			.SO(gen[6979]),
			.S(gen[6980]),
			.SE(gen[6981]),

			.SELF(gen[6885]),
			.cell_state(gen[6885])
		); 

/******************* CELL 6886 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6886 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6790]),
			.N(gen[6791]),
			.NE(gen[6792]),

			.O(gen[6885]),
			.E(gen[6887]),

			.SO(gen[6980]),
			.S(gen[6981]),
			.SE(gen[6982]),

			.SELF(gen[6886]),
			.cell_state(gen[6886])
		); 

/******************* CELL 6887 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6887 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6791]),
			.N(gen[6792]),
			.NE(gen[6793]),

			.O(gen[6886]),
			.E(gen[6888]),

			.SO(gen[6981]),
			.S(gen[6982]),
			.SE(gen[6983]),

			.SELF(gen[6887]),
			.cell_state(gen[6887])
		); 

/******************* CELL 6888 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6888 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6792]),
			.N(gen[6793]),
			.NE(gen[6794]),

			.O(gen[6887]),
			.E(gen[6889]),

			.SO(gen[6982]),
			.S(gen[6983]),
			.SE(gen[6984]),

			.SELF(gen[6888]),
			.cell_state(gen[6888])
		); 

/******************* CELL 6889 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6889 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6793]),
			.N(gen[6794]),
			.NE(gen[6795]),

			.O(gen[6888]),
			.E(gen[6890]),

			.SO(gen[6983]),
			.S(gen[6984]),
			.SE(gen[6985]),

			.SELF(gen[6889]),
			.cell_state(gen[6889])
		); 

/******************* CELL 6890 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6890 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6794]),
			.N(gen[6795]),
			.NE(gen[6796]),

			.O(gen[6889]),
			.E(gen[6891]),

			.SO(gen[6984]),
			.S(gen[6985]),
			.SE(gen[6986]),

			.SELF(gen[6890]),
			.cell_state(gen[6890])
		); 

/******************* CELL 6891 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6891 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6795]),
			.N(gen[6796]),
			.NE(gen[6797]),

			.O(gen[6890]),
			.E(gen[6892]),

			.SO(gen[6985]),
			.S(gen[6986]),
			.SE(gen[6987]),

			.SELF(gen[6891]),
			.cell_state(gen[6891])
		); 

/******************* CELL 6892 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6892 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6796]),
			.N(gen[6797]),
			.NE(gen[6798]),

			.O(gen[6891]),
			.E(gen[6893]),

			.SO(gen[6986]),
			.S(gen[6987]),
			.SE(gen[6988]),

			.SELF(gen[6892]),
			.cell_state(gen[6892])
		); 

/******************* CELL 6893 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6893 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6797]),
			.N(gen[6798]),
			.NE(gen[6799]),

			.O(gen[6892]),
			.E(gen[6894]),

			.SO(gen[6987]),
			.S(gen[6988]),
			.SE(gen[6989]),

			.SELF(gen[6893]),
			.cell_state(gen[6893])
		); 

/******************* CELL 6894 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6894 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6798]),
			.N(gen[6799]),
			.NE(gen[6800]),

			.O(gen[6893]),
			.E(gen[6895]),

			.SO(gen[6988]),
			.S(gen[6989]),
			.SE(gen[6990]),

			.SELF(gen[6894]),
			.cell_state(gen[6894])
		); 

/******************* CELL 6895 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6895 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6799]),
			.N(gen[6800]),
			.NE(gen[6801]),

			.O(gen[6894]),
			.E(gen[6896]),

			.SO(gen[6989]),
			.S(gen[6990]),
			.SE(gen[6991]),

			.SELF(gen[6895]),
			.cell_state(gen[6895])
		); 

/******************* CELL 6896 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6896 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6800]),
			.N(gen[6801]),
			.NE(gen[6802]),

			.O(gen[6895]),
			.E(gen[6897]),

			.SO(gen[6990]),
			.S(gen[6991]),
			.SE(gen[6992]),

			.SELF(gen[6896]),
			.cell_state(gen[6896])
		); 

/******************* CELL 6897 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6897 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6801]),
			.N(gen[6802]),
			.NE(gen[6803]),

			.O(gen[6896]),
			.E(gen[6898]),

			.SO(gen[6991]),
			.S(gen[6992]),
			.SE(gen[6993]),

			.SELF(gen[6897]),
			.cell_state(gen[6897])
		); 

/******************* CELL 6898 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6898 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6802]),
			.N(gen[6803]),
			.NE(gen[6804]),

			.O(gen[6897]),
			.E(gen[6899]),

			.SO(gen[6992]),
			.S(gen[6993]),
			.SE(gen[6994]),

			.SELF(gen[6898]),
			.cell_state(gen[6898])
		); 

/******************* CELL 6899 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6899 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6803]),
			.N(gen[6804]),
			.NE(gen[6805]),

			.O(gen[6898]),
			.E(gen[6900]),

			.SO(gen[6993]),
			.S(gen[6994]),
			.SE(gen[6995]),

			.SELF(gen[6899]),
			.cell_state(gen[6899])
		); 

/******************* CELL 6900 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6900 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6804]),
			.N(gen[6805]),
			.NE(gen[6806]),

			.O(gen[6899]),
			.E(gen[6901]),

			.SO(gen[6994]),
			.S(gen[6995]),
			.SE(gen[6996]),

			.SELF(gen[6900]),
			.cell_state(gen[6900])
		); 

/******************* CELL 6901 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6901 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6805]),
			.N(gen[6806]),
			.NE(gen[6807]),

			.O(gen[6900]),
			.E(gen[6902]),

			.SO(gen[6995]),
			.S(gen[6996]),
			.SE(gen[6997]),

			.SELF(gen[6901]),
			.cell_state(gen[6901])
		); 

/******************* CELL 6902 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6902 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6806]),
			.N(gen[6807]),
			.NE(gen[6808]),

			.O(gen[6901]),
			.E(gen[6903]),

			.SO(gen[6996]),
			.S(gen[6997]),
			.SE(gen[6998]),

			.SELF(gen[6902]),
			.cell_state(gen[6902])
		); 

/******************* CELL 6903 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6903 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6807]),
			.N(gen[6808]),
			.NE(gen[6809]),

			.O(gen[6902]),
			.E(gen[6904]),

			.SO(gen[6997]),
			.S(gen[6998]),
			.SE(gen[6999]),

			.SELF(gen[6903]),
			.cell_state(gen[6903])
		); 

/******************* CELL 6904 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6904 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6808]),
			.N(gen[6809]),
			.NE(gen[6810]),

			.O(gen[6903]),
			.E(gen[6905]),

			.SO(gen[6998]),
			.S(gen[6999]),
			.SE(gen[7000]),

			.SELF(gen[6904]),
			.cell_state(gen[6904])
		); 

/******************* CELL 6905 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6905 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6809]),
			.N(gen[6810]),
			.NE(gen[6811]),

			.O(gen[6904]),
			.E(gen[6906]),

			.SO(gen[6999]),
			.S(gen[7000]),
			.SE(gen[7001]),

			.SELF(gen[6905]),
			.cell_state(gen[6905])
		); 

/******************* CELL 6906 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6906 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6810]),
			.N(gen[6811]),
			.NE(gen[6812]),

			.O(gen[6905]),
			.E(gen[6907]),

			.SO(gen[7000]),
			.S(gen[7001]),
			.SE(gen[7002]),

			.SELF(gen[6906]),
			.cell_state(gen[6906])
		); 

/******************* CELL 6907 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6907 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6811]),
			.N(gen[6812]),
			.NE(gen[6813]),

			.O(gen[6906]),
			.E(gen[6908]),

			.SO(gen[7001]),
			.S(gen[7002]),
			.SE(gen[7003]),

			.SELF(gen[6907]),
			.cell_state(gen[6907])
		); 

/******************* CELL 6908 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6908 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6812]),
			.N(gen[6813]),
			.NE(gen[6814]),

			.O(gen[6907]),
			.E(gen[6909]),

			.SO(gen[7002]),
			.S(gen[7003]),
			.SE(gen[7004]),

			.SELF(gen[6908]),
			.cell_state(gen[6908])
		); 

/******************* CELL 6909 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6909 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6813]),
			.N(gen[6814]),
			.NE(gen[6815]),

			.O(gen[6908]),
			.E(gen[6910]),

			.SO(gen[7003]),
			.S(gen[7004]),
			.SE(gen[7005]),

			.SELF(gen[6909]),
			.cell_state(gen[6909])
		); 

/******************* CELL 6910 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6910 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6814]),
			.N(gen[6815]),
			.NE(gen[6816]),

			.O(gen[6909]),
			.E(gen[6911]),

			.SO(gen[7004]),
			.S(gen[7005]),
			.SE(gen[7006]),

			.SELF(gen[6910]),
			.cell_state(gen[6910])
		); 

/******************* CELL 6911 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6911 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6815]),
			.N(gen[6816]),
			.NE(gen[6817]),

			.O(gen[6910]),
			.E(gen[6912]),

			.SO(gen[7005]),
			.S(gen[7006]),
			.SE(gen[7007]),

			.SELF(gen[6911]),
			.cell_state(gen[6911])
		); 

/******************* CELL 6912 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6912 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6816]),
			.N(gen[6817]),
			.NE(gen[6818]),

			.O(gen[6911]),
			.E(gen[6913]),

			.SO(gen[7006]),
			.S(gen[7007]),
			.SE(gen[7008]),

			.SELF(gen[6912]),
			.cell_state(gen[6912])
		); 

/******************* CELL 6913 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6913 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6817]),
			.N(gen[6818]),
			.NE(gen[6819]),

			.O(gen[6912]),
			.E(gen[6914]),

			.SO(gen[7007]),
			.S(gen[7008]),
			.SE(gen[7009]),

			.SELF(gen[6913]),
			.cell_state(gen[6913])
		); 

/******************* CELL 6914 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6914 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6818]),
			.N(gen[6819]),
			.NE(gen[6820]),

			.O(gen[6913]),
			.E(gen[6915]),

			.SO(gen[7008]),
			.S(gen[7009]),
			.SE(gen[7010]),

			.SELF(gen[6914]),
			.cell_state(gen[6914])
		); 

/******************* CELL 6915 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6915 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6819]),
			.N(gen[6820]),
			.NE(gen[6821]),

			.O(gen[6914]),
			.E(gen[6916]),

			.SO(gen[7009]),
			.S(gen[7010]),
			.SE(gen[7011]),

			.SELF(gen[6915]),
			.cell_state(gen[6915])
		); 

/******************* CELL 6916 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6916 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6820]),
			.N(gen[6821]),
			.NE(gen[6822]),

			.O(gen[6915]),
			.E(gen[6917]),

			.SO(gen[7010]),
			.S(gen[7011]),
			.SE(gen[7012]),

			.SELF(gen[6916]),
			.cell_state(gen[6916])
		); 

/******************* CELL 6917 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6917 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6821]),
			.N(gen[6822]),
			.NE(gen[6823]),

			.O(gen[6916]),
			.E(gen[6918]),

			.SO(gen[7011]),
			.S(gen[7012]),
			.SE(gen[7013]),

			.SELF(gen[6917]),
			.cell_state(gen[6917])
		); 

/******************* CELL 6918 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6918 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6822]),
			.N(gen[6823]),
			.NE(gen[6824]),

			.O(gen[6917]),
			.E(gen[6919]),

			.SO(gen[7012]),
			.S(gen[7013]),
			.SE(gen[7014]),

			.SELF(gen[6918]),
			.cell_state(gen[6918])
		); 

/******************* CELL 6919 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6919 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6823]),
			.N(gen[6824]),
			.NE(gen[6825]),

			.O(gen[6918]),
			.E(gen[6920]),

			.SO(gen[7013]),
			.S(gen[7014]),
			.SE(gen[7015]),

			.SELF(gen[6919]),
			.cell_state(gen[6919])
		); 

/******************* CELL 6920 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6920 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6824]),
			.N(gen[6825]),
			.NE(gen[6826]),

			.O(gen[6919]),
			.E(gen[6921]),

			.SO(gen[7014]),
			.S(gen[7015]),
			.SE(gen[7016]),

			.SELF(gen[6920]),
			.cell_state(gen[6920])
		); 

/******************* CELL 6921 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6921 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6825]),
			.N(gen[6826]),
			.NE(gen[6827]),

			.O(gen[6920]),
			.E(gen[6922]),

			.SO(gen[7015]),
			.S(gen[7016]),
			.SE(gen[7017]),

			.SELF(gen[6921]),
			.cell_state(gen[6921])
		); 

/******************* CELL 6922 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6922 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6826]),
			.N(gen[6827]),
			.NE(gen[6828]),

			.O(gen[6921]),
			.E(gen[6923]),

			.SO(gen[7016]),
			.S(gen[7017]),
			.SE(gen[7018]),

			.SELF(gen[6922]),
			.cell_state(gen[6922])
		); 

/******************* CELL 6923 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6923 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6827]),
			.N(gen[6828]),
			.NE(gen[6829]),

			.O(gen[6922]),
			.E(gen[6924]),

			.SO(gen[7017]),
			.S(gen[7018]),
			.SE(gen[7019]),

			.SELF(gen[6923]),
			.cell_state(gen[6923])
		); 

/******************* CELL 6924 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6924 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6828]),
			.N(gen[6829]),
			.NE(gen[6830]),

			.O(gen[6923]),
			.E(gen[6925]),

			.SO(gen[7018]),
			.S(gen[7019]),
			.SE(gen[7020]),

			.SELF(gen[6924]),
			.cell_state(gen[6924])
		); 

/******************* CELL 6925 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6925 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6829]),
			.N(gen[6830]),
			.NE(gen[6831]),

			.O(gen[6924]),
			.E(gen[6926]),

			.SO(gen[7019]),
			.S(gen[7020]),
			.SE(gen[7021]),

			.SELF(gen[6925]),
			.cell_state(gen[6925])
		); 

/******************* CELL 6926 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6926 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6830]),
			.N(gen[6831]),
			.NE(gen[6832]),

			.O(gen[6925]),
			.E(gen[6927]),

			.SO(gen[7020]),
			.S(gen[7021]),
			.SE(gen[7022]),

			.SELF(gen[6926]),
			.cell_state(gen[6926])
		); 

/******************* CELL 6927 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6927 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6831]),
			.N(gen[6832]),
			.NE(gen[6833]),

			.O(gen[6926]),
			.E(gen[6928]),

			.SO(gen[7021]),
			.S(gen[7022]),
			.SE(gen[7023]),

			.SELF(gen[6927]),
			.cell_state(gen[6927])
		); 

/******************* CELL 6928 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6928 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6832]),
			.N(gen[6833]),
			.NE(gen[6834]),

			.O(gen[6927]),
			.E(gen[6929]),

			.SO(gen[7022]),
			.S(gen[7023]),
			.SE(gen[7024]),

			.SELF(gen[6928]),
			.cell_state(gen[6928])
		); 

/******************* CELL 6929 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6929 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6833]),
			.N(gen[6834]),
			.NE(gen[6835]),

			.O(gen[6928]),
			.E(gen[6930]),

			.SO(gen[7023]),
			.S(gen[7024]),
			.SE(gen[7025]),

			.SELF(gen[6929]),
			.cell_state(gen[6929])
		); 

/******************* CELL 6930 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6930 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6834]),
			.N(gen[6835]),
			.NE(gen[6836]),

			.O(gen[6929]),
			.E(gen[6931]),

			.SO(gen[7024]),
			.S(gen[7025]),
			.SE(gen[7026]),

			.SELF(gen[6930]),
			.cell_state(gen[6930])
		); 

/******************* CELL 6931 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6931 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6835]),
			.N(gen[6836]),
			.NE(gen[6837]),

			.O(gen[6930]),
			.E(gen[6932]),

			.SO(gen[7025]),
			.S(gen[7026]),
			.SE(gen[7027]),

			.SELF(gen[6931]),
			.cell_state(gen[6931])
		); 

/******************* CELL 6932 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6932 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6836]),
			.N(gen[6837]),
			.NE(gen[6838]),

			.O(gen[6931]),
			.E(gen[6933]),

			.SO(gen[7026]),
			.S(gen[7027]),
			.SE(gen[7028]),

			.SELF(gen[6932]),
			.cell_state(gen[6932])
		); 

/******************* CELL 6933 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6933 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6837]),
			.N(gen[6838]),
			.NE(gen[6839]),

			.O(gen[6932]),
			.E(gen[6934]),

			.SO(gen[7027]),
			.S(gen[7028]),
			.SE(gen[7029]),

			.SELF(gen[6933]),
			.cell_state(gen[6933])
		); 

/******************* CELL 6934 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6934 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6838]),
			.N(gen[6839]),
			.NE(gen[6838]),

			.O(gen[6933]),
			.E(gen[6933]),

			.SO(gen[7028]),
			.S(gen[7029]),
			.SE(gen[7028]),

			.SELF(gen[6934]),
			.cell_state(gen[6934])
		); 

/******************* CELL 6935 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6935 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6841]),
			.N(gen[6840]),
			.NE(gen[6841]),

			.O(gen[6936]),
			.E(gen[6936]),

			.SO(gen[7031]),
			.S(gen[7030]),
			.SE(gen[7031]),

			.SELF(gen[6935]),
			.cell_state(gen[6935])
		); 

/******************* CELL 6936 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6936 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6840]),
			.N(gen[6841]),
			.NE(gen[6842]),

			.O(gen[6935]),
			.E(gen[6937]),

			.SO(gen[7030]),
			.S(gen[7031]),
			.SE(gen[7032]),

			.SELF(gen[6936]),
			.cell_state(gen[6936])
		); 

/******************* CELL 6937 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6937 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6841]),
			.N(gen[6842]),
			.NE(gen[6843]),

			.O(gen[6936]),
			.E(gen[6938]),

			.SO(gen[7031]),
			.S(gen[7032]),
			.SE(gen[7033]),

			.SELF(gen[6937]),
			.cell_state(gen[6937])
		); 

/******************* CELL 6938 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6938 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6842]),
			.N(gen[6843]),
			.NE(gen[6844]),

			.O(gen[6937]),
			.E(gen[6939]),

			.SO(gen[7032]),
			.S(gen[7033]),
			.SE(gen[7034]),

			.SELF(gen[6938]),
			.cell_state(gen[6938])
		); 

/******************* CELL 6939 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6939 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6843]),
			.N(gen[6844]),
			.NE(gen[6845]),

			.O(gen[6938]),
			.E(gen[6940]),

			.SO(gen[7033]),
			.S(gen[7034]),
			.SE(gen[7035]),

			.SELF(gen[6939]),
			.cell_state(gen[6939])
		); 

/******************* CELL 6940 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6940 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6844]),
			.N(gen[6845]),
			.NE(gen[6846]),

			.O(gen[6939]),
			.E(gen[6941]),

			.SO(gen[7034]),
			.S(gen[7035]),
			.SE(gen[7036]),

			.SELF(gen[6940]),
			.cell_state(gen[6940])
		); 

/******************* CELL 6941 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6941 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6845]),
			.N(gen[6846]),
			.NE(gen[6847]),

			.O(gen[6940]),
			.E(gen[6942]),

			.SO(gen[7035]),
			.S(gen[7036]),
			.SE(gen[7037]),

			.SELF(gen[6941]),
			.cell_state(gen[6941])
		); 

/******************* CELL 6942 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6942 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6846]),
			.N(gen[6847]),
			.NE(gen[6848]),

			.O(gen[6941]),
			.E(gen[6943]),

			.SO(gen[7036]),
			.S(gen[7037]),
			.SE(gen[7038]),

			.SELF(gen[6942]),
			.cell_state(gen[6942])
		); 

/******************* CELL 6943 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6943 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6847]),
			.N(gen[6848]),
			.NE(gen[6849]),

			.O(gen[6942]),
			.E(gen[6944]),

			.SO(gen[7037]),
			.S(gen[7038]),
			.SE(gen[7039]),

			.SELF(gen[6943]),
			.cell_state(gen[6943])
		); 

/******************* CELL 6944 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6944 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6848]),
			.N(gen[6849]),
			.NE(gen[6850]),

			.O(gen[6943]),
			.E(gen[6945]),

			.SO(gen[7038]),
			.S(gen[7039]),
			.SE(gen[7040]),

			.SELF(gen[6944]),
			.cell_state(gen[6944])
		); 

/******************* CELL 6945 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6945 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6849]),
			.N(gen[6850]),
			.NE(gen[6851]),

			.O(gen[6944]),
			.E(gen[6946]),

			.SO(gen[7039]),
			.S(gen[7040]),
			.SE(gen[7041]),

			.SELF(gen[6945]),
			.cell_state(gen[6945])
		); 

/******************* CELL 6946 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6946 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6850]),
			.N(gen[6851]),
			.NE(gen[6852]),

			.O(gen[6945]),
			.E(gen[6947]),

			.SO(gen[7040]),
			.S(gen[7041]),
			.SE(gen[7042]),

			.SELF(gen[6946]),
			.cell_state(gen[6946])
		); 

/******************* CELL 6947 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6947 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6851]),
			.N(gen[6852]),
			.NE(gen[6853]),

			.O(gen[6946]),
			.E(gen[6948]),

			.SO(gen[7041]),
			.S(gen[7042]),
			.SE(gen[7043]),

			.SELF(gen[6947]),
			.cell_state(gen[6947])
		); 

/******************* CELL 6948 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6948 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6852]),
			.N(gen[6853]),
			.NE(gen[6854]),

			.O(gen[6947]),
			.E(gen[6949]),

			.SO(gen[7042]),
			.S(gen[7043]),
			.SE(gen[7044]),

			.SELF(gen[6948]),
			.cell_state(gen[6948])
		); 

/******************* CELL 6949 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6949 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6853]),
			.N(gen[6854]),
			.NE(gen[6855]),

			.O(gen[6948]),
			.E(gen[6950]),

			.SO(gen[7043]),
			.S(gen[7044]),
			.SE(gen[7045]),

			.SELF(gen[6949]),
			.cell_state(gen[6949])
		); 

/******************* CELL 6950 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6950 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6854]),
			.N(gen[6855]),
			.NE(gen[6856]),

			.O(gen[6949]),
			.E(gen[6951]),

			.SO(gen[7044]),
			.S(gen[7045]),
			.SE(gen[7046]),

			.SELF(gen[6950]),
			.cell_state(gen[6950])
		); 

/******************* CELL 6951 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6951 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6855]),
			.N(gen[6856]),
			.NE(gen[6857]),

			.O(gen[6950]),
			.E(gen[6952]),

			.SO(gen[7045]),
			.S(gen[7046]),
			.SE(gen[7047]),

			.SELF(gen[6951]),
			.cell_state(gen[6951])
		); 

/******************* CELL 6952 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6952 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6856]),
			.N(gen[6857]),
			.NE(gen[6858]),

			.O(gen[6951]),
			.E(gen[6953]),

			.SO(gen[7046]),
			.S(gen[7047]),
			.SE(gen[7048]),

			.SELF(gen[6952]),
			.cell_state(gen[6952])
		); 

/******************* CELL 6953 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6953 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6857]),
			.N(gen[6858]),
			.NE(gen[6859]),

			.O(gen[6952]),
			.E(gen[6954]),

			.SO(gen[7047]),
			.S(gen[7048]),
			.SE(gen[7049]),

			.SELF(gen[6953]),
			.cell_state(gen[6953])
		); 

/******************* CELL 6954 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6954 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6858]),
			.N(gen[6859]),
			.NE(gen[6860]),

			.O(gen[6953]),
			.E(gen[6955]),

			.SO(gen[7048]),
			.S(gen[7049]),
			.SE(gen[7050]),

			.SELF(gen[6954]),
			.cell_state(gen[6954])
		); 

/******************* CELL 6955 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6955 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6859]),
			.N(gen[6860]),
			.NE(gen[6861]),

			.O(gen[6954]),
			.E(gen[6956]),

			.SO(gen[7049]),
			.S(gen[7050]),
			.SE(gen[7051]),

			.SELF(gen[6955]),
			.cell_state(gen[6955])
		); 

/******************* CELL 6956 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6956 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6860]),
			.N(gen[6861]),
			.NE(gen[6862]),

			.O(gen[6955]),
			.E(gen[6957]),

			.SO(gen[7050]),
			.S(gen[7051]),
			.SE(gen[7052]),

			.SELF(gen[6956]),
			.cell_state(gen[6956])
		); 

/******************* CELL 6957 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6957 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6861]),
			.N(gen[6862]),
			.NE(gen[6863]),

			.O(gen[6956]),
			.E(gen[6958]),

			.SO(gen[7051]),
			.S(gen[7052]),
			.SE(gen[7053]),

			.SELF(gen[6957]),
			.cell_state(gen[6957])
		); 

/******************* CELL 6958 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6958 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6862]),
			.N(gen[6863]),
			.NE(gen[6864]),

			.O(gen[6957]),
			.E(gen[6959]),

			.SO(gen[7052]),
			.S(gen[7053]),
			.SE(gen[7054]),

			.SELF(gen[6958]),
			.cell_state(gen[6958])
		); 

/******************* CELL 6959 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6959 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6863]),
			.N(gen[6864]),
			.NE(gen[6865]),

			.O(gen[6958]),
			.E(gen[6960]),

			.SO(gen[7053]),
			.S(gen[7054]),
			.SE(gen[7055]),

			.SELF(gen[6959]),
			.cell_state(gen[6959])
		); 

/******************* CELL 6960 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6960 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6864]),
			.N(gen[6865]),
			.NE(gen[6866]),

			.O(gen[6959]),
			.E(gen[6961]),

			.SO(gen[7054]),
			.S(gen[7055]),
			.SE(gen[7056]),

			.SELF(gen[6960]),
			.cell_state(gen[6960])
		); 

/******************* CELL 6961 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6961 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6865]),
			.N(gen[6866]),
			.NE(gen[6867]),

			.O(gen[6960]),
			.E(gen[6962]),

			.SO(gen[7055]),
			.S(gen[7056]),
			.SE(gen[7057]),

			.SELF(gen[6961]),
			.cell_state(gen[6961])
		); 

/******************* CELL 6962 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6962 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6866]),
			.N(gen[6867]),
			.NE(gen[6868]),

			.O(gen[6961]),
			.E(gen[6963]),

			.SO(gen[7056]),
			.S(gen[7057]),
			.SE(gen[7058]),

			.SELF(gen[6962]),
			.cell_state(gen[6962])
		); 

/******************* CELL 6963 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6963 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6867]),
			.N(gen[6868]),
			.NE(gen[6869]),

			.O(gen[6962]),
			.E(gen[6964]),

			.SO(gen[7057]),
			.S(gen[7058]),
			.SE(gen[7059]),

			.SELF(gen[6963]),
			.cell_state(gen[6963])
		); 

/******************* CELL 6964 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6964 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6868]),
			.N(gen[6869]),
			.NE(gen[6870]),

			.O(gen[6963]),
			.E(gen[6965]),

			.SO(gen[7058]),
			.S(gen[7059]),
			.SE(gen[7060]),

			.SELF(gen[6964]),
			.cell_state(gen[6964])
		); 

/******************* CELL 6965 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6965 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6869]),
			.N(gen[6870]),
			.NE(gen[6871]),

			.O(gen[6964]),
			.E(gen[6966]),

			.SO(gen[7059]),
			.S(gen[7060]),
			.SE(gen[7061]),

			.SELF(gen[6965]),
			.cell_state(gen[6965])
		); 

/******************* CELL 6966 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6966 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6870]),
			.N(gen[6871]),
			.NE(gen[6872]),

			.O(gen[6965]),
			.E(gen[6967]),

			.SO(gen[7060]),
			.S(gen[7061]),
			.SE(gen[7062]),

			.SELF(gen[6966]),
			.cell_state(gen[6966])
		); 

/******************* CELL 6967 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6967 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6871]),
			.N(gen[6872]),
			.NE(gen[6873]),

			.O(gen[6966]),
			.E(gen[6968]),

			.SO(gen[7061]),
			.S(gen[7062]),
			.SE(gen[7063]),

			.SELF(gen[6967]),
			.cell_state(gen[6967])
		); 

/******************* CELL 6968 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6968 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6872]),
			.N(gen[6873]),
			.NE(gen[6874]),

			.O(gen[6967]),
			.E(gen[6969]),

			.SO(gen[7062]),
			.S(gen[7063]),
			.SE(gen[7064]),

			.SELF(gen[6968]),
			.cell_state(gen[6968])
		); 

/******************* CELL 6969 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6969 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6873]),
			.N(gen[6874]),
			.NE(gen[6875]),

			.O(gen[6968]),
			.E(gen[6970]),

			.SO(gen[7063]),
			.S(gen[7064]),
			.SE(gen[7065]),

			.SELF(gen[6969]),
			.cell_state(gen[6969])
		); 

/******************* CELL 6970 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6970 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6874]),
			.N(gen[6875]),
			.NE(gen[6876]),

			.O(gen[6969]),
			.E(gen[6971]),

			.SO(gen[7064]),
			.S(gen[7065]),
			.SE(gen[7066]),

			.SELF(gen[6970]),
			.cell_state(gen[6970])
		); 

/******************* CELL 6971 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6971 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6875]),
			.N(gen[6876]),
			.NE(gen[6877]),

			.O(gen[6970]),
			.E(gen[6972]),

			.SO(gen[7065]),
			.S(gen[7066]),
			.SE(gen[7067]),

			.SELF(gen[6971]),
			.cell_state(gen[6971])
		); 

/******************* CELL 6972 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6972 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6876]),
			.N(gen[6877]),
			.NE(gen[6878]),

			.O(gen[6971]),
			.E(gen[6973]),

			.SO(gen[7066]),
			.S(gen[7067]),
			.SE(gen[7068]),

			.SELF(gen[6972]),
			.cell_state(gen[6972])
		); 

/******************* CELL 6973 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6973 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6877]),
			.N(gen[6878]),
			.NE(gen[6879]),

			.O(gen[6972]),
			.E(gen[6974]),

			.SO(gen[7067]),
			.S(gen[7068]),
			.SE(gen[7069]),

			.SELF(gen[6973]),
			.cell_state(gen[6973])
		); 

/******************* CELL 6974 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6974 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6878]),
			.N(gen[6879]),
			.NE(gen[6880]),

			.O(gen[6973]),
			.E(gen[6975]),

			.SO(gen[7068]),
			.S(gen[7069]),
			.SE(gen[7070]),

			.SELF(gen[6974]),
			.cell_state(gen[6974])
		); 

/******************* CELL 6975 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6975 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6879]),
			.N(gen[6880]),
			.NE(gen[6881]),

			.O(gen[6974]),
			.E(gen[6976]),

			.SO(gen[7069]),
			.S(gen[7070]),
			.SE(gen[7071]),

			.SELF(gen[6975]),
			.cell_state(gen[6975])
		); 

/******************* CELL 6976 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6976 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6880]),
			.N(gen[6881]),
			.NE(gen[6882]),

			.O(gen[6975]),
			.E(gen[6977]),

			.SO(gen[7070]),
			.S(gen[7071]),
			.SE(gen[7072]),

			.SELF(gen[6976]),
			.cell_state(gen[6976])
		); 

/******************* CELL 6977 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6977 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6881]),
			.N(gen[6882]),
			.NE(gen[6883]),

			.O(gen[6976]),
			.E(gen[6978]),

			.SO(gen[7071]),
			.S(gen[7072]),
			.SE(gen[7073]),

			.SELF(gen[6977]),
			.cell_state(gen[6977])
		); 

/******************* CELL 6978 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6978 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6882]),
			.N(gen[6883]),
			.NE(gen[6884]),

			.O(gen[6977]),
			.E(gen[6979]),

			.SO(gen[7072]),
			.S(gen[7073]),
			.SE(gen[7074]),

			.SELF(gen[6978]),
			.cell_state(gen[6978])
		); 

/******************* CELL 6979 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6979 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6883]),
			.N(gen[6884]),
			.NE(gen[6885]),

			.O(gen[6978]),
			.E(gen[6980]),

			.SO(gen[7073]),
			.S(gen[7074]),
			.SE(gen[7075]),

			.SELF(gen[6979]),
			.cell_state(gen[6979])
		); 

/******************* CELL 6980 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6980 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6884]),
			.N(gen[6885]),
			.NE(gen[6886]),

			.O(gen[6979]),
			.E(gen[6981]),

			.SO(gen[7074]),
			.S(gen[7075]),
			.SE(gen[7076]),

			.SELF(gen[6980]),
			.cell_state(gen[6980])
		); 

/******************* CELL 6981 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6981 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6885]),
			.N(gen[6886]),
			.NE(gen[6887]),

			.O(gen[6980]),
			.E(gen[6982]),

			.SO(gen[7075]),
			.S(gen[7076]),
			.SE(gen[7077]),

			.SELF(gen[6981]),
			.cell_state(gen[6981])
		); 

/******************* CELL 6982 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6982 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6886]),
			.N(gen[6887]),
			.NE(gen[6888]),

			.O(gen[6981]),
			.E(gen[6983]),

			.SO(gen[7076]),
			.S(gen[7077]),
			.SE(gen[7078]),

			.SELF(gen[6982]),
			.cell_state(gen[6982])
		); 

/******************* CELL 6983 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6983 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6887]),
			.N(gen[6888]),
			.NE(gen[6889]),

			.O(gen[6982]),
			.E(gen[6984]),

			.SO(gen[7077]),
			.S(gen[7078]),
			.SE(gen[7079]),

			.SELF(gen[6983]),
			.cell_state(gen[6983])
		); 

/******************* CELL 6984 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6984 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6888]),
			.N(gen[6889]),
			.NE(gen[6890]),

			.O(gen[6983]),
			.E(gen[6985]),

			.SO(gen[7078]),
			.S(gen[7079]),
			.SE(gen[7080]),

			.SELF(gen[6984]),
			.cell_state(gen[6984])
		); 

/******************* CELL 6985 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6985 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6889]),
			.N(gen[6890]),
			.NE(gen[6891]),

			.O(gen[6984]),
			.E(gen[6986]),

			.SO(gen[7079]),
			.S(gen[7080]),
			.SE(gen[7081]),

			.SELF(gen[6985]),
			.cell_state(gen[6985])
		); 

/******************* CELL 6986 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6986 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6890]),
			.N(gen[6891]),
			.NE(gen[6892]),

			.O(gen[6985]),
			.E(gen[6987]),

			.SO(gen[7080]),
			.S(gen[7081]),
			.SE(gen[7082]),

			.SELF(gen[6986]),
			.cell_state(gen[6986])
		); 

/******************* CELL 6987 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6987 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6891]),
			.N(gen[6892]),
			.NE(gen[6893]),

			.O(gen[6986]),
			.E(gen[6988]),

			.SO(gen[7081]),
			.S(gen[7082]),
			.SE(gen[7083]),

			.SELF(gen[6987]),
			.cell_state(gen[6987])
		); 

/******************* CELL 6988 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6988 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6892]),
			.N(gen[6893]),
			.NE(gen[6894]),

			.O(gen[6987]),
			.E(gen[6989]),

			.SO(gen[7082]),
			.S(gen[7083]),
			.SE(gen[7084]),

			.SELF(gen[6988]),
			.cell_state(gen[6988])
		); 

/******************* CELL 6989 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6989 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6893]),
			.N(gen[6894]),
			.NE(gen[6895]),

			.O(gen[6988]),
			.E(gen[6990]),

			.SO(gen[7083]),
			.S(gen[7084]),
			.SE(gen[7085]),

			.SELF(gen[6989]),
			.cell_state(gen[6989])
		); 

/******************* CELL 6990 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6990 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6894]),
			.N(gen[6895]),
			.NE(gen[6896]),

			.O(gen[6989]),
			.E(gen[6991]),

			.SO(gen[7084]),
			.S(gen[7085]),
			.SE(gen[7086]),

			.SELF(gen[6990]),
			.cell_state(gen[6990])
		); 

/******************* CELL 6991 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6991 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6895]),
			.N(gen[6896]),
			.NE(gen[6897]),

			.O(gen[6990]),
			.E(gen[6992]),

			.SO(gen[7085]),
			.S(gen[7086]),
			.SE(gen[7087]),

			.SELF(gen[6991]),
			.cell_state(gen[6991])
		); 

/******************* CELL 6992 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6992 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6896]),
			.N(gen[6897]),
			.NE(gen[6898]),

			.O(gen[6991]),
			.E(gen[6993]),

			.SO(gen[7086]),
			.S(gen[7087]),
			.SE(gen[7088]),

			.SELF(gen[6992]),
			.cell_state(gen[6992])
		); 

/******************* CELL 6993 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6993 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6897]),
			.N(gen[6898]),
			.NE(gen[6899]),

			.O(gen[6992]),
			.E(gen[6994]),

			.SO(gen[7087]),
			.S(gen[7088]),
			.SE(gen[7089]),

			.SELF(gen[6993]),
			.cell_state(gen[6993])
		); 

/******************* CELL 6994 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6994 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6898]),
			.N(gen[6899]),
			.NE(gen[6900]),

			.O(gen[6993]),
			.E(gen[6995]),

			.SO(gen[7088]),
			.S(gen[7089]),
			.SE(gen[7090]),

			.SELF(gen[6994]),
			.cell_state(gen[6994])
		); 

/******************* CELL 6995 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6995 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6899]),
			.N(gen[6900]),
			.NE(gen[6901]),

			.O(gen[6994]),
			.E(gen[6996]),

			.SO(gen[7089]),
			.S(gen[7090]),
			.SE(gen[7091]),

			.SELF(gen[6995]),
			.cell_state(gen[6995])
		); 

/******************* CELL 6996 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6996 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6900]),
			.N(gen[6901]),
			.NE(gen[6902]),

			.O(gen[6995]),
			.E(gen[6997]),

			.SO(gen[7090]),
			.S(gen[7091]),
			.SE(gen[7092]),

			.SELF(gen[6996]),
			.cell_state(gen[6996])
		); 

/******************* CELL 6997 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6997 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6901]),
			.N(gen[6902]),
			.NE(gen[6903]),

			.O(gen[6996]),
			.E(gen[6998]),

			.SO(gen[7091]),
			.S(gen[7092]),
			.SE(gen[7093]),

			.SELF(gen[6997]),
			.cell_state(gen[6997])
		); 

/******************* CELL 6998 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6998 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6902]),
			.N(gen[6903]),
			.NE(gen[6904]),

			.O(gen[6997]),
			.E(gen[6999]),

			.SO(gen[7092]),
			.S(gen[7093]),
			.SE(gen[7094]),

			.SELF(gen[6998]),
			.cell_state(gen[6998])
		); 

/******************* CELL 6999 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell6999 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6903]),
			.N(gen[6904]),
			.NE(gen[6905]),

			.O(gen[6998]),
			.E(gen[7000]),

			.SO(gen[7093]),
			.S(gen[7094]),
			.SE(gen[7095]),

			.SELF(gen[6999]),
			.cell_state(gen[6999])
		); 

/******************* CELL 7000 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7000 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6904]),
			.N(gen[6905]),
			.NE(gen[6906]),

			.O(gen[6999]),
			.E(gen[7001]),

			.SO(gen[7094]),
			.S(gen[7095]),
			.SE(gen[7096]),

			.SELF(gen[7000]),
			.cell_state(gen[7000])
		); 

/******************* CELL 7001 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7001 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6905]),
			.N(gen[6906]),
			.NE(gen[6907]),

			.O(gen[7000]),
			.E(gen[7002]),

			.SO(gen[7095]),
			.S(gen[7096]),
			.SE(gen[7097]),

			.SELF(gen[7001]),
			.cell_state(gen[7001])
		); 

/******************* CELL 7002 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7002 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6906]),
			.N(gen[6907]),
			.NE(gen[6908]),

			.O(gen[7001]),
			.E(gen[7003]),

			.SO(gen[7096]),
			.S(gen[7097]),
			.SE(gen[7098]),

			.SELF(gen[7002]),
			.cell_state(gen[7002])
		); 

/******************* CELL 7003 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7003 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6907]),
			.N(gen[6908]),
			.NE(gen[6909]),

			.O(gen[7002]),
			.E(gen[7004]),

			.SO(gen[7097]),
			.S(gen[7098]),
			.SE(gen[7099]),

			.SELF(gen[7003]),
			.cell_state(gen[7003])
		); 

/******************* CELL 7004 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7004 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6908]),
			.N(gen[6909]),
			.NE(gen[6910]),

			.O(gen[7003]),
			.E(gen[7005]),

			.SO(gen[7098]),
			.S(gen[7099]),
			.SE(gen[7100]),

			.SELF(gen[7004]),
			.cell_state(gen[7004])
		); 

/******************* CELL 7005 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7005 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6909]),
			.N(gen[6910]),
			.NE(gen[6911]),

			.O(gen[7004]),
			.E(gen[7006]),

			.SO(gen[7099]),
			.S(gen[7100]),
			.SE(gen[7101]),

			.SELF(gen[7005]),
			.cell_state(gen[7005])
		); 

/******************* CELL 7006 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7006 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6910]),
			.N(gen[6911]),
			.NE(gen[6912]),

			.O(gen[7005]),
			.E(gen[7007]),

			.SO(gen[7100]),
			.S(gen[7101]),
			.SE(gen[7102]),

			.SELF(gen[7006]),
			.cell_state(gen[7006])
		); 

/******************* CELL 7007 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7007 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6911]),
			.N(gen[6912]),
			.NE(gen[6913]),

			.O(gen[7006]),
			.E(gen[7008]),

			.SO(gen[7101]),
			.S(gen[7102]),
			.SE(gen[7103]),

			.SELF(gen[7007]),
			.cell_state(gen[7007])
		); 

/******************* CELL 7008 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7008 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6912]),
			.N(gen[6913]),
			.NE(gen[6914]),

			.O(gen[7007]),
			.E(gen[7009]),

			.SO(gen[7102]),
			.S(gen[7103]),
			.SE(gen[7104]),

			.SELF(gen[7008]),
			.cell_state(gen[7008])
		); 

/******************* CELL 7009 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7009 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6913]),
			.N(gen[6914]),
			.NE(gen[6915]),

			.O(gen[7008]),
			.E(gen[7010]),

			.SO(gen[7103]),
			.S(gen[7104]),
			.SE(gen[7105]),

			.SELF(gen[7009]),
			.cell_state(gen[7009])
		); 

/******************* CELL 7010 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7010 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6914]),
			.N(gen[6915]),
			.NE(gen[6916]),

			.O(gen[7009]),
			.E(gen[7011]),

			.SO(gen[7104]),
			.S(gen[7105]),
			.SE(gen[7106]),

			.SELF(gen[7010]),
			.cell_state(gen[7010])
		); 

/******************* CELL 7011 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7011 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6915]),
			.N(gen[6916]),
			.NE(gen[6917]),

			.O(gen[7010]),
			.E(gen[7012]),

			.SO(gen[7105]),
			.S(gen[7106]),
			.SE(gen[7107]),

			.SELF(gen[7011]),
			.cell_state(gen[7011])
		); 

/******************* CELL 7012 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7012 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6916]),
			.N(gen[6917]),
			.NE(gen[6918]),

			.O(gen[7011]),
			.E(gen[7013]),

			.SO(gen[7106]),
			.S(gen[7107]),
			.SE(gen[7108]),

			.SELF(gen[7012]),
			.cell_state(gen[7012])
		); 

/******************* CELL 7013 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7013 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6917]),
			.N(gen[6918]),
			.NE(gen[6919]),

			.O(gen[7012]),
			.E(gen[7014]),

			.SO(gen[7107]),
			.S(gen[7108]),
			.SE(gen[7109]),

			.SELF(gen[7013]),
			.cell_state(gen[7013])
		); 

/******************* CELL 7014 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7014 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6918]),
			.N(gen[6919]),
			.NE(gen[6920]),

			.O(gen[7013]),
			.E(gen[7015]),

			.SO(gen[7108]),
			.S(gen[7109]),
			.SE(gen[7110]),

			.SELF(gen[7014]),
			.cell_state(gen[7014])
		); 

/******************* CELL 7015 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7015 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6919]),
			.N(gen[6920]),
			.NE(gen[6921]),

			.O(gen[7014]),
			.E(gen[7016]),

			.SO(gen[7109]),
			.S(gen[7110]),
			.SE(gen[7111]),

			.SELF(gen[7015]),
			.cell_state(gen[7015])
		); 

/******************* CELL 7016 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7016 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6920]),
			.N(gen[6921]),
			.NE(gen[6922]),

			.O(gen[7015]),
			.E(gen[7017]),

			.SO(gen[7110]),
			.S(gen[7111]),
			.SE(gen[7112]),

			.SELF(gen[7016]),
			.cell_state(gen[7016])
		); 

/******************* CELL 7017 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7017 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6921]),
			.N(gen[6922]),
			.NE(gen[6923]),

			.O(gen[7016]),
			.E(gen[7018]),

			.SO(gen[7111]),
			.S(gen[7112]),
			.SE(gen[7113]),

			.SELF(gen[7017]),
			.cell_state(gen[7017])
		); 

/******************* CELL 7018 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7018 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6922]),
			.N(gen[6923]),
			.NE(gen[6924]),

			.O(gen[7017]),
			.E(gen[7019]),

			.SO(gen[7112]),
			.S(gen[7113]),
			.SE(gen[7114]),

			.SELF(gen[7018]),
			.cell_state(gen[7018])
		); 

/******************* CELL 7019 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7019 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6923]),
			.N(gen[6924]),
			.NE(gen[6925]),

			.O(gen[7018]),
			.E(gen[7020]),

			.SO(gen[7113]),
			.S(gen[7114]),
			.SE(gen[7115]),

			.SELF(gen[7019]),
			.cell_state(gen[7019])
		); 

/******************* CELL 7020 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7020 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6924]),
			.N(gen[6925]),
			.NE(gen[6926]),

			.O(gen[7019]),
			.E(gen[7021]),

			.SO(gen[7114]),
			.S(gen[7115]),
			.SE(gen[7116]),

			.SELF(gen[7020]),
			.cell_state(gen[7020])
		); 

/******************* CELL 7021 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7021 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6925]),
			.N(gen[6926]),
			.NE(gen[6927]),

			.O(gen[7020]),
			.E(gen[7022]),

			.SO(gen[7115]),
			.S(gen[7116]),
			.SE(gen[7117]),

			.SELF(gen[7021]),
			.cell_state(gen[7021])
		); 

/******************* CELL 7022 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7022 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6926]),
			.N(gen[6927]),
			.NE(gen[6928]),

			.O(gen[7021]),
			.E(gen[7023]),

			.SO(gen[7116]),
			.S(gen[7117]),
			.SE(gen[7118]),

			.SELF(gen[7022]),
			.cell_state(gen[7022])
		); 

/******************* CELL 7023 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7023 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6927]),
			.N(gen[6928]),
			.NE(gen[6929]),

			.O(gen[7022]),
			.E(gen[7024]),

			.SO(gen[7117]),
			.S(gen[7118]),
			.SE(gen[7119]),

			.SELF(gen[7023]),
			.cell_state(gen[7023])
		); 

/******************* CELL 7024 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7024 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6928]),
			.N(gen[6929]),
			.NE(gen[6930]),

			.O(gen[7023]),
			.E(gen[7025]),

			.SO(gen[7118]),
			.S(gen[7119]),
			.SE(gen[7120]),

			.SELF(gen[7024]),
			.cell_state(gen[7024])
		); 

/******************* CELL 7025 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7025 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6929]),
			.N(gen[6930]),
			.NE(gen[6931]),

			.O(gen[7024]),
			.E(gen[7026]),

			.SO(gen[7119]),
			.S(gen[7120]),
			.SE(gen[7121]),

			.SELF(gen[7025]),
			.cell_state(gen[7025])
		); 

/******************* CELL 7026 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7026 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6930]),
			.N(gen[6931]),
			.NE(gen[6932]),

			.O(gen[7025]),
			.E(gen[7027]),

			.SO(gen[7120]),
			.S(gen[7121]),
			.SE(gen[7122]),

			.SELF(gen[7026]),
			.cell_state(gen[7026])
		); 

/******************* CELL 7027 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7027 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6931]),
			.N(gen[6932]),
			.NE(gen[6933]),

			.O(gen[7026]),
			.E(gen[7028]),

			.SO(gen[7121]),
			.S(gen[7122]),
			.SE(gen[7123]),

			.SELF(gen[7027]),
			.cell_state(gen[7027])
		); 

/******************* CELL 7028 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7028 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6932]),
			.N(gen[6933]),
			.NE(gen[6934]),

			.O(gen[7027]),
			.E(gen[7029]),

			.SO(gen[7122]),
			.S(gen[7123]),
			.SE(gen[7124]),

			.SELF(gen[7028]),
			.cell_state(gen[7028])
		); 

/******************* CELL 7029 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7029 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6933]),
			.N(gen[6934]),
			.NE(gen[6933]),

			.O(gen[7028]),
			.E(gen[7028]),

			.SO(gen[7123]),
			.S(gen[7124]),
			.SE(gen[7123]),

			.SELF(gen[7029]),
			.cell_state(gen[7029])
		); 

/******************* CELL 7030 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7030 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6936]),
			.N(gen[6935]),
			.NE(gen[6936]),

			.O(gen[7031]),
			.E(gen[7031]),

			.SO(gen[7126]),
			.S(gen[7125]),
			.SE(gen[7126]),

			.SELF(gen[7030]),
			.cell_state(gen[7030])
		); 

/******************* CELL 7031 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7031 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6935]),
			.N(gen[6936]),
			.NE(gen[6937]),

			.O(gen[7030]),
			.E(gen[7032]),

			.SO(gen[7125]),
			.S(gen[7126]),
			.SE(gen[7127]),

			.SELF(gen[7031]),
			.cell_state(gen[7031])
		); 

/******************* CELL 7032 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7032 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6936]),
			.N(gen[6937]),
			.NE(gen[6938]),

			.O(gen[7031]),
			.E(gen[7033]),

			.SO(gen[7126]),
			.S(gen[7127]),
			.SE(gen[7128]),

			.SELF(gen[7032]),
			.cell_state(gen[7032])
		); 

/******************* CELL 7033 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7033 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6937]),
			.N(gen[6938]),
			.NE(gen[6939]),

			.O(gen[7032]),
			.E(gen[7034]),

			.SO(gen[7127]),
			.S(gen[7128]),
			.SE(gen[7129]),

			.SELF(gen[7033]),
			.cell_state(gen[7033])
		); 

/******************* CELL 7034 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7034 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6938]),
			.N(gen[6939]),
			.NE(gen[6940]),

			.O(gen[7033]),
			.E(gen[7035]),

			.SO(gen[7128]),
			.S(gen[7129]),
			.SE(gen[7130]),

			.SELF(gen[7034]),
			.cell_state(gen[7034])
		); 

/******************* CELL 7035 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7035 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6939]),
			.N(gen[6940]),
			.NE(gen[6941]),

			.O(gen[7034]),
			.E(gen[7036]),

			.SO(gen[7129]),
			.S(gen[7130]),
			.SE(gen[7131]),

			.SELF(gen[7035]),
			.cell_state(gen[7035])
		); 

/******************* CELL 7036 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7036 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6940]),
			.N(gen[6941]),
			.NE(gen[6942]),

			.O(gen[7035]),
			.E(gen[7037]),

			.SO(gen[7130]),
			.S(gen[7131]),
			.SE(gen[7132]),

			.SELF(gen[7036]),
			.cell_state(gen[7036])
		); 

/******************* CELL 7037 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7037 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6941]),
			.N(gen[6942]),
			.NE(gen[6943]),

			.O(gen[7036]),
			.E(gen[7038]),

			.SO(gen[7131]),
			.S(gen[7132]),
			.SE(gen[7133]),

			.SELF(gen[7037]),
			.cell_state(gen[7037])
		); 

/******************* CELL 7038 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7038 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6942]),
			.N(gen[6943]),
			.NE(gen[6944]),

			.O(gen[7037]),
			.E(gen[7039]),

			.SO(gen[7132]),
			.S(gen[7133]),
			.SE(gen[7134]),

			.SELF(gen[7038]),
			.cell_state(gen[7038])
		); 

/******************* CELL 7039 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7039 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6943]),
			.N(gen[6944]),
			.NE(gen[6945]),

			.O(gen[7038]),
			.E(gen[7040]),

			.SO(gen[7133]),
			.S(gen[7134]),
			.SE(gen[7135]),

			.SELF(gen[7039]),
			.cell_state(gen[7039])
		); 

/******************* CELL 7040 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7040 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6944]),
			.N(gen[6945]),
			.NE(gen[6946]),

			.O(gen[7039]),
			.E(gen[7041]),

			.SO(gen[7134]),
			.S(gen[7135]),
			.SE(gen[7136]),

			.SELF(gen[7040]),
			.cell_state(gen[7040])
		); 

/******************* CELL 7041 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7041 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6945]),
			.N(gen[6946]),
			.NE(gen[6947]),

			.O(gen[7040]),
			.E(gen[7042]),

			.SO(gen[7135]),
			.S(gen[7136]),
			.SE(gen[7137]),

			.SELF(gen[7041]),
			.cell_state(gen[7041])
		); 

/******************* CELL 7042 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7042 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6946]),
			.N(gen[6947]),
			.NE(gen[6948]),

			.O(gen[7041]),
			.E(gen[7043]),

			.SO(gen[7136]),
			.S(gen[7137]),
			.SE(gen[7138]),

			.SELF(gen[7042]),
			.cell_state(gen[7042])
		); 

/******************* CELL 7043 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7043 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6947]),
			.N(gen[6948]),
			.NE(gen[6949]),

			.O(gen[7042]),
			.E(gen[7044]),

			.SO(gen[7137]),
			.S(gen[7138]),
			.SE(gen[7139]),

			.SELF(gen[7043]),
			.cell_state(gen[7043])
		); 

/******************* CELL 7044 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7044 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6948]),
			.N(gen[6949]),
			.NE(gen[6950]),

			.O(gen[7043]),
			.E(gen[7045]),

			.SO(gen[7138]),
			.S(gen[7139]),
			.SE(gen[7140]),

			.SELF(gen[7044]),
			.cell_state(gen[7044])
		); 

/******************* CELL 7045 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7045 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6949]),
			.N(gen[6950]),
			.NE(gen[6951]),

			.O(gen[7044]),
			.E(gen[7046]),

			.SO(gen[7139]),
			.S(gen[7140]),
			.SE(gen[7141]),

			.SELF(gen[7045]),
			.cell_state(gen[7045])
		); 

/******************* CELL 7046 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7046 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6950]),
			.N(gen[6951]),
			.NE(gen[6952]),

			.O(gen[7045]),
			.E(gen[7047]),

			.SO(gen[7140]),
			.S(gen[7141]),
			.SE(gen[7142]),

			.SELF(gen[7046]),
			.cell_state(gen[7046])
		); 

/******************* CELL 7047 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7047 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6951]),
			.N(gen[6952]),
			.NE(gen[6953]),

			.O(gen[7046]),
			.E(gen[7048]),

			.SO(gen[7141]),
			.S(gen[7142]),
			.SE(gen[7143]),

			.SELF(gen[7047]),
			.cell_state(gen[7047])
		); 

/******************* CELL 7048 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7048 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6952]),
			.N(gen[6953]),
			.NE(gen[6954]),

			.O(gen[7047]),
			.E(gen[7049]),

			.SO(gen[7142]),
			.S(gen[7143]),
			.SE(gen[7144]),

			.SELF(gen[7048]),
			.cell_state(gen[7048])
		); 

/******************* CELL 7049 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7049 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6953]),
			.N(gen[6954]),
			.NE(gen[6955]),

			.O(gen[7048]),
			.E(gen[7050]),

			.SO(gen[7143]),
			.S(gen[7144]),
			.SE(gen[7145]),

			.SELF(gen[7049]),
			.cell_state(gen[7049])
		); 

/******************* CELL 7050 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7050 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6954]),
			.N(gen[6955]),
			.NE(gen[6956]),

			.O(gen[7049]),
			.E(gen[7051]),

			.SO(gen[7144]),
			.S(gen[7145]),
			.SE(gen[7146]),

			.SELF(gen[7050]),
			.cell_state(gen[7050])
		); 

/******************* CELL 7051 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7051 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6955]),
			.N(gen[6956]),
			.NE(gen[6957]),

			.O(gen[7050]),
			.E(gen[7052]),

			.SO(gen[7145]),
			.S(gen[7146]),
			.SE(gen[7147]),

			.SELF(gen[7051]),
			.cell_state(gen[7051])
		); 

/******************* CELL 7052 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7052 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6956]),
			.N(gen[6957]),
			.NE(gen[6958]),

			.O(gen[7051]),
			.E(gen[7053]),

			.SO(gen[7146]),
			.S(gen[7147]),
			.SE(gen[7148]),

			.SELF(gen[7052]),
			.cell_state(gen[7052])
		); 

/******************* CELL 7053 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7053 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6957]),
			.N(gen[6958]),
			.NE(gen[6959]),

			.O(gen[7052]),
			.E(gen[7054]),

			.SO(gen[7147]),
			.S(gen[7148]),
			.SE(gen[7149]),

			.SELF(gen[7053]),
			.cell_state(gen[7053])
		); 

/******************* CELL 7054 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7054 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6958]),
			.N(gen[6959]),
			.NE(gen[6960]),

			.O(gen[7053]),
			.E(gen[7055]),

			.SO(gen[7148]),
			.S(gen[7149]),
			.SE(gen[7150]),

			.SELF(gen[7054]),
			.cell_state(gen[7054])
		); 

/******************* CELL 7055 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7055 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6959]),
			.N(gen[6960]),
			.NE(gen[6961]),

			.O(gen[7054]),
			.E(gen[7056]),

			.SO(gen[7149]),
			.S(gen[7150]),
			.SE(gen[7151]),

			.SELF(gen[7055]),
			.cell_state(gen[7055])
		); 

/******************* CELL 7056 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7056 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6960]),
			.N(gen[6961]),
			.NE(gen[6962]),

			.O(gen[7055]),
			.E(gen[7057]),

			.SO(gen[7150]),
			.S(gen[7151]),
			.SE(gen[7152]),

			.SELF(gen[7056]),
			.cell_state(gen[7056])
		); 

/******************* CELL 7057 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7057 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6961]),
			.N(gen[6962]),
			.NE(gen[6963]),

			.O(gen[7056]),
			.E(gen[7058]),

			.SO(gen[7151]),
			.S(gen[7152]),
			.SE(gen[7153]),

			.SELF(gen[7057]),
			.cell_state(gen[7057])
		); 

/******************* CELL 7058 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7058 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6962]),
			.N(gen[6963]),
			.NE(gen[6964]),

			.O(gen[7057]),
			.E(gen[7059]),

			.SO(gen[7152]),
			.S(gen[7153]),
			.SE(gen[7154]),

			.SELF(gen[7058]),
			.cell_state(gen[7058])
		); 

/******************* CELL 7059 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7059 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6963]),
			.N(gen[6964]),
			.NE(gen[6965]),

			.O(gen[7058]),
			.E(gen[7060]),

			.SO(gen[7153]),
			.S(gen[7154]),
			.SE(gen[7155]),

			.SELF(gen[7059]),
			.cell_state(gen[7059])
		); 

/******************* CELL 7060 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7060 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6964]),
			.N(gen[6965]),
			.NE(gen[6966]),

			.O(gen[7059]),
			.E(gen[7061]),

			.SO(gen[7154]),
			.S(gen[7155]),
			.SE(gen[7156]),

			.SELF(gen[7060]),
			.cell_state(gen[7060])
		); 

/******************* CELL 7061 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7061 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6965]),
			.N(gen[6966]),
			.NE(gen[6967]),

			.O(gen[7060]),
			.E(gen[7062]),

			.SO(gen[7155]),
			.S(gen[7156]),
			.SE(gen[7157]),

			.SELF(gen[7061]),
			.cell_state(gen[7061])
		); 

/******************* CELL 7062 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7062 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6966]),
			.N(gen[6967]),
			.NE(gen[6968]),

			.O(gen[7061]),
			.E(gen[7063]),

			.SO(gen[7156]),
			.S(gen[7157]),
			.SE(gen[7158]),

			.SELF(gen[7062]),
			.cell_state(gen[7062])
		); 

/******************* CELL 7063 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7063 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6967]),
			.N(gen[6968]),
			.NE(gen[6969]),

			.O(gen[7062]),
			.E(gen[7064]),

			.SO(gen[7157]),
			.S(gen[7158]),
			.SE(gen[7159]),

			.SELF(gen[7063]),
			.cell_state(gen[7063])
		); 

/******************* CELL 7064 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7064 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6968]),
			.N(gen[6969]),
			.NE(gen[6970]),

			.O(gen[7063]),
			.E(gen[7065]),

			.SO(gen[7158]),
			.S(gen[7159]),
			.SE(gen[7160]),

			.SELF(gen[7064]),
			.cell_state(gen[7064])
		); 

/******************* CELL 7065 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7065 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6969]),
			.N(gen[6970]),
			.NE(gen[6971]),

			.O(gen[7064]),
			.E(gen[7066]),

			.SO(gen[7159]),
			.S(gen[7160]),
			.SE(gen[7161]),

			.SELF(gen[7065]),
			.cell_state(gen[7065])
		); 

/******************* CELL 7066 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7066 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6970]),
			.N(gen[6971]),
			.NE(gen[6972]),

			.O(gen[7065]),
			.E(gen[7067]),

			.SO(gen[7160]),
			.S(gen[7161]),
			.SE(gen[7162]),

			.SELF(gen[7066]),
			.cell_state(gen[7066])
		); 

/******************* CELL 7067 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7067 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6971]),
			.N(gen[6972]),
			.NE(gen[6973]),

			.O(gen[7066]),
			.E(gen[7068]),

			.SO(gen[7161]),
			.S(gen[7162]),
			.SE(gen[7163]),

			.SELF(gen[7067]),
			.cell_state(gen[7067])
		); 

/******************* CELL 7068 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7068 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6972]),
			.N(gen[6973]),
			.NE(gen[6974]),

			.O(gen[7067]),
			.E(gen[7069]),

			.SO(gen[7162]),
			.S(gen[7163]),
			.SE(gen[7164]),

			.SELF(gen[7068]),
			.cell_state(gen[7068])
		); 

/******************* CELL 7069 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7069 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6973]),
			.N(gen[6974]),
			.NE(gen[6975]),

			.O(gen[7068]),
			.E(gen[7070]),

			.SO(gen[7163]),
			.S(gen[7164]),
			.SE(gen[7165]),

			.SELF(gen[7069]),
			.cell_state(gen[7069])
		); 

/******************* CELL 7070 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7070 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6974]),
			.N(gen[6975]),
			.NE(gen[6976]),

			.O(gen[7069]),
			.E(gen[7071]),

			.SO(gen[7164]),
			.S(gen[7165]),
			.SE(gen[7166]),

			.SELF(gen[7070]),
			.cell_state(gen[7070])
		); 

/******************* CELL 7071 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7071 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6975]),
			.N(gen[6976]),
			.NE(gen[6977]),

			.O(gen[7070]),
			.E(gen[7072]),

			.SO(gen[7165]),
			.S(gen[7166]),
			.SE(gen[7167]),

			.SELF(gen[7071]),
			.cell_state(gen[7071])
		); 

/******************* CELL 7072 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7072 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6976]),
			.N(gen[6977]),
			.NE(gen[6978]),

			.O(gen[7071]),
			.E(gen[7073]),

			.SO(gen[7166]),
			.S(gen[7167]),
			.SE(gen[7168]),

			.SELF(gen[7072]),
			.cell_state(gen[7072])
		); 

/******************* CELL 7073 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7073 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6977]),
			.N(gen[6978]),
			.NE(gen[6979]),

			.O(gen[7072]),
			.E(gen[7074]),

			.SO(gen[7167]),
			.S(gen[7168]),
			.SE(gen[7169]),

			.SELF(gen[7073]),
			.cell_state(gen[7073])
		); 

/******************* CELL 7074 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7074 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6978]),
			.N(gen[6979]),
			.NE(gen[6980]),

			.O(gen[7073]),
			.E(gen[7075]),

			.SO(gen[7168]),
			.S(gen[7169]),
			.SE(gen[7170]),

			.SELF(gen[7074]),
			.cell_state(gen[7074])
		); 

/******************* CELL 7075 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7075 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6979]),
			.N(gen[6980]),
			.NE(gen[6981]),

			.O(gen[7074]),
			.E(gen[7076]),

			.SO(gen[7169]),
			.S(gen[7170]),
			.SE(gen[7171]),

			.SELF(gen[7075]),
			.cell_state(gen[7075])
		); 

/******************* CELL 7076 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7076 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6980]),
			.N(gen[6981]),
			.NE(gen[6982]),

			.O(gen[7075]),
			.E(gen[7077]),

			.SO(gen[7170]),
			.S(gen[7171]),
			.SE(gen[7172]),

			.SELF(gen[7076]),
			.cell_state(gen[7076])
		); 

/******************* CELL 7077 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7077 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6981]),
			.N(gen[6982]),
			.NE(gen[6983]),

			.O(gen[7076]),
			.E(gen[7078]),

			.SO(gen[7171]),
			.S(gen[7172]),
			.SE(gen[7173]),

			.SELF(gen[7077]),
			.cell_state(gen[7077])
		); 

/******************* CELL 7078 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7078 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6982]),
			.N(gen[6983]),
			.NE(gen[6984]),

			.O(gen[7077]),
			.E(gen[7079]),

			.SO(gen[7172]),
			.S(gen[7173]),
			.SE(gen[7174]),

			.SELF(gen[7078]),
			.cell_state(gen[7078])
		); 

/******************* CELL 7079 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7079 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6983]),
			.N(gen[6984]),
			.NE(gen[6985]),

			.O(gen[7078]),
			.E(gen[7080]),

			.SO(gen[7173]),
			.S(gen[7174]),
			.SE(gen[7175]),

			.SELF(gen[7079]),
			.cell_state(gen[7079])
		); 

/******************* CELL 7080 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7080 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6984]),
			.N(gen[6985]),
			.NE(gen[6986]),

			.O(gen[7079]),
			.E(gen[7081]),

			.SO(gen[7174]),
			.S(gen[7175]),
			.SE(gen[7176]),

			.SELF(gen[7080]),
			.cell_state(gen[7080])
		); 

/******************* CELL 7081 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7081 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6985]),
			.N(gen[6986]),
			.NE(gen[6987]),

			.O(gen[7080]),
			.E(gen[7082]),

			.SO(gen[7175]),
			.S(gen[7176]),
			.SE(gen[7177]),

			.SELF(gen[7081]),
			.cell_state(gen[7081])
		); 

/******************* CELL 7082 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7082 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6986]),
			.N(gen[6987]),
			.NE(gen[6988]),

			.O(gen[7081]),
			.E(gen[7083]),

			.SO(gen[7176]),
			.S(gen[7177]),
			.SE(gen[7178]),

			.SELF(gen[7082]),
			.cell_state(gen[7082])
		); 

/******************* CELL 7083 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7083 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6987]),
			.N(gen[6988]),
			.NE(gen[6989]),

			.O(gen[7082]),
			.E(gen[7084]),

			.SO(gen[7177]),
			.S(gen[7178]),
			.SE(gen[7179]),

			.SELF(gen[7083]),
			.cell_state(gen[7083])
		); 

/******************* CELL 7084 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7084 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6988]),
			.N(gen[6989]),
			.NE(gen[6990]),

			.O(gen[7083]),
			.E(gen[7085]),

			.SO(gen[7178]),
			.S(gen[7179]),
			.SE(gen[7180]),

			.SELF(gen[7084]),
			.cell_state(gen[7084])
		); 

/******************* CELL 7085 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7085 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6989]),
			.N(gen[6990]),
			.NE(gen[6991]),

			.O(gen[7084]),
			.E(gen[7086]),

			.SO(gen[7179]),
			.S(gen[7180]),
			.SE(gen[7181]),

			.SELF(gen[7085]),
			.cell_state(gen[7085])
		); 

/******************* CELL 7086 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7086 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6990]),
			.N(gen[6991]),
			.NE(gen[6992]),

			.O(gen[7085]),
			.E(gen[7087]),

			.SO(gen[7180]),
			.S(gen[7181]),
			.SE(gen[7182]),

			.SELF(gen[7086]),
			.cell_state(gen[7086])
		); 

/******************* CELL 7087 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7087 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6991]),
			.N(gen[6992]),
			.NE(gen[6993]),

			.O(gen[7086]),
			.E(gen[7088]),

			.SO(gen[7181]),
			.S(gen[7182]),
			.SE(gen[7183]),

			.SELF(gen[7087]),
			.cell_state(gen[7087])
		); 

/******************* CELL 7088 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7088 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6992]),
			.N(gen[6993]),
			.NE(gen[6994]),

			.O(gen[7087]),
			.E(gen[7089]),

			.SO(gen[7182]),
			.S(gen[7183]),
			.SE(gen[7184]),

			.SELF(gen[7088]),
			.cell_state(gen[7088])
		); 

/******************* CELL 7089 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7089 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6993]),
			.N(gen[6994]),
			.NE(gen[6995]),

			.O(gen[7088]),
			.E(gen[7090]),

			.SO(gen[7183]),
			.S(gen[7184]),
			.SE(gen[7185]),

			.SELF(gen[7089]),
			.cell_state(gen[7089])
		); 

/******************* CELL 7090 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7090 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6994]),
			.N(gen[6995]),
			.NE(gen[6996]),

			.O(gen[7089]),
			.E(gen[7091]),

			.SO(gen[7184]),
			.S(gen[7185]),
			.SE(gen[7186]),

			.SELF(gen[7090]),
			.cell_state(gen[7090])
		); 

/******************* CELL 7091 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7091 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6995]),
			.N(gen[6996]),
			.NE(gen[6997]),

			.O(gen[7090]),
			.E(gen[7092]),

			.SO(gen[7185]),
			.S(gen[7186]),
			.SE(gen[7187]),

			.SELF(gen[7091]),
			.cell_state(gen[7091])
		); 

/******************* CELL 7092 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7092 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6996]),
			.N(gen[6997]),
			.NE(gen[6998]),

			.O(gen[7091]),
			.E(gen[7093]),

			.SO(gen[7186]),
			.S(gen[7187]),
			.SE(gen[7188]),

			.SELF(gen[7092]),
			.cell_state(gen[7092])
		); 

/******************* CELL 7093 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7093 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6997]),
			.N(gen[6998]),
			.NE(gen[6999]),

			.O(gen[7092]),
			.E(gen[7094]),

			.SO(gen[7187]),
			.S(gen[7188]),
			.SE(gen[7189]),

			.SELF(gen[7093]),
			.cell_state(gen[7093])
		); 

/******************* CELL 7094 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7094 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6998]),
			.N(gen[6999]),
			.NE(gen[7000]),

			.O(gen[7093]),
			.E(gen[7095]),

			.SO(gen[7188]),
			.S(gen[7189]),
			.SE(gen[7190]),

			.SELF(gen[7094]),
			.cell_state(gen[7094])
		); 

/******************* CELL 7095 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7095 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6999]),
			.N(gen[7000]),
			.NE(gen[7001]),

			.O(gen[7094]),
			.E(gen[7096]),

			.SO(gen[7189]),
			.S(gen[7190]),
			.SE(gen[7191]),

			.SELF(gen[7095]),
			.cell_state(gen[7095])
		); 

/******************* CELL 7096 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7096 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7000]),
			.N(gen[7001]),
			.NE(gen[7002]),

			.O(gen[7095]),
			.E(gen[7097]),

			.SO(gen[7190]),
			.S(gen[7191]),
			.SE(gen[7192]),

			.SELF(gen[7096]),
			.cell_state(gen[7096])
		); 

/******************* CELL 7097 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7097 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7001]),
			.N(gen[7002]),
			.NE(gen[7003]),

			.O(gen[7096]),
			.E(gen[7098]),

			.SO(gen[7191]),
			.S(gen[7192]),
			.SE(gen[7193]),

			.SELF(gen[7097]),
			.cell_state(gen[7097])
		); 

/******************* CELL 7098 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7098 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7002]),
			.N(gen[7003]),
			.NE(gen[7004]),

			.O(gen[7097]),
			.E(gen[7099]),

			.SO(gen[7192]),
			.S(gen[7193]),
			.SE(gen[7194]),

			.SELF(gen[7098]),
			.cell_state(gen[7098])
		); 

/******************* CELL 7099 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7099 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7003]),
			.N(gen[7004]),
			.NE(gen[7005]),

			.O(gen[7098]),
			.E(gen[7100]),

			.SO(gen[7193]),
			.S(gen[7194]),
			.SE(gen[7195]),

			.SELF(gen[7099]),
			.cell_state(gen[7099])
		); 

/******************* CELL 7100 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7100 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7004]),
			.N(gen[7005]),
			.NE(gen[7006]),

			.O(gen[7099]),
			.E(gen[7101]),

			.SO(gen[7194]),
			.S(gen[7195]),
			.SE(gen[7196]),

			.SELF(gen[7100]),
			.cell_state(gen[7100])
		); 

/******************* CELL 7101 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7101 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7005]),
			.N(gen[7006]),
			.NE(gen[7007]),

			.O(gen[7100]),
			.E(gen[7102]),

			.SO(gen[7195]),
			.S(gen[7196]),
			.SE(gen[7197]),

			.SELF(gen[7101]),
			.cell_state(gen[7101])
		); 

/******************* CELL 7102 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7102 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7006]),
			.N(gen[7007]),
			.NE(gen[7008]),

			.O(gen[7101]),
			.E(gen[7103]),

			.SO(gen[7196]),
			.S(gen[7197]),
			.SE(gen[7198]),

			.SELF(gen[7102]),
			.cell_state(gen[7102])
		); 

/******************* CELL 7103 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7103 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7007]),
			.N(gen[7008]),
			.NE(gen[7009]),

			.O(gen[7102]),
			.E(gen[7104]),

			.SO(gen[7197]),
			.S(gen[7198]),
			.SE(gen[7199]),

			.SELF(gen[7103]),
			.cell_state(gen[7103])
		); 

/******************* CELL 7104 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7104 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7008]),
			.N(gen[7009]),
			.NE(gen[7010]),

			.O(gen[7103]),
			.E(gen[7105]),

			.SO(gen[7198]),
			.S(gen[7199]),
			.SE(gen[7200]),

			.SELF(gen[7104]),
			.cell_state(gen[7104])
		); 

/******************* CELL 7105 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7105 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7009]),
			.N(gen[7010]),
			.NE(gen[7011]),

			.O(gen[7104]),
			.E(gen[7106]),

			.SO(gen[7199]),
			.S(gen[7200]),
			.SE(gen[7201]),

			.SELF(gen[7105]),
			.cell_state(gen[7105])
		); 

/******************* CELL 7106 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7106 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7010]),
			.N(gen[7011]),
			.NE(gen[7012]),

			.O(gen[7105]),
			.E(gen[7107]),

			.SO(gen[7200]),
			.S(gen[7201]),
			.SE(gen[7202]),

			.SELF(gen[7106]),
			.cell_state(gen[7106])
		); 

/******************* CELL 7107 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7107 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7011]),
			.N(gen[7012]),
			.NE(gen[7013]),

			.O(gen[7106]),
			.E(gen[7108]),

			.SO(gen[7201]),
			.S(gen[7202]),
			.SE(gen[7203]),

			.SELF(gen[7107]),
			.cell_state(gen[7107])
		); 

/******************* CELL 7108 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7108 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7012]),
			.N(gen[7013]),
			.NE(gen[7014]),

			.O(gen[7107]),
			.E(gen[7109]),

			.SO(gen[7202]),
			.S(gen[7203]),
			.SE(gen[7204]),

			.SELF(gen[7108]),
			.cell_state(gen[7108])
		); 

/******************* CELL 7109 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7109 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7013]),
			.N(gen[7014]),
			.NE(gen[7015]),

			.O(gen[7108]),
			.E(gen[7110]),

			.SO(gen[7203]),
			.S(gen[7204]),
			.SE(gen[7205]),

			.SELF(gen[7109]),
			.cell_state(gen[7109])
		); 

/******************* CELL 7110 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7110 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7014]),
			.N(gen[7015]),
			.NE(gen[7016]),

			.O(gen[7109]),
			.E(gen[7111]),

			.SO(gen[7204]),
			.S(gen[7205]),
			.SE(gen[7206]),

			.SELF(gen[7110]),
			.cell_state(gen[7110])
		); 

/******************* CELL 7111 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7111 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7015]),
			.N(gen[7016]),
			.NE(gen[7017]),

			.O(gen[7110]),
			.E(gen[7112]),

			.SO(gen[7205]),
			.S(gen[7206]),
			.SE(gen[7207]),

			.SELF(gen[7111]),
			.cell_state(gen[7111])
		); 

/******************* CELL 7112 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7112 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7016]),
			.N(gen[7017]),
			.NE(gen[7018]),

			.O(gen[7111]),
			.E(gen[7113]),

			.SO(gen[7206]),
			.S(gen[7207]),
			.SE(gen[7208]),

			.SELF(gen[7112]),
			.cell_state(gen[7112])
		); 

/******************* CELL 7113 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7113 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7017]),
			.N(gen[7018]),
			.NE(gen[7019]),

			.O(gen[7112]),
			.E(gen[7114]),

			.SO(gen[7207]),
			.S(gen[7208]),
			.SE(gen[7209]),

			.SELF(gen[7113]),
			.cell_state(gen[7113])
		); 

/******************* CELL 7114 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7114 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7018]),
			.N(gen[7019]),
			.NE(gen[7020]),

			.O(gen[7113]),
			.E(gen[7115]),

			.SO(gen[7208]),
			.S(gen[7209]),
			.SE(gen[7210]),

			.SELF(gen[7114]),
			.cell_state(gen[7114])
		); 

/******************* CELL 7115 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7115 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7019]),
			.N(gen[7020]),
			.NE(gen[7021]),

			.O(gen[7114]),
			.E(gen[7116]),

			.SO(gen[7209]),
			.S(gen[7210]),
			.SE(gen[7211]),

			.SELF(gen[7115]),
			.cell_state(gen[7115])
		); 

/******************* CELL 7116 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7116 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7020]),
			.N(gen[7021]),
			.NE(gen[7022]),

			.O(gen[7115]),
			.E(gen[7117]),

			.SO(gen[7210]),
			.S(gen[7211]),
			.SE(gen[7212]),

			.SELF(gen[7116]),
			.cell_state(gen[7116])
		); 

/******************* CELL 7117 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7117 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7021]),
			.N(gen[7022]),
			.NE(gen[7023]),

			.O(gen[7116]),
			.E(gen[7118]),

			.SO(gen[7211]),
			.S(gen[7212]),
			.SE(gen[7213]),

			.SELF(gen[7117]),
			.cell_state(gen[7117])
		); 

/******************* CELL 7118 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7118 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7022]),
			.N(gen[7023]),
			.NE(gen[7024]),

			.O(gen[7117]),
			.E(gen[7119]),

			.SO(gen[7212]),
			.S(gen[7213]),
			.SE(gen[7214]),

			.SELF(gen[7118]),
			.cell_state(gen[7118])
		); 

/******************* CELL 7119 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7119 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7023]),
			.N(gen[7024]),
			.NE(gen[7025]),

			.O(gen[7118]),
			.E(gen[7120]),

			.SO(gen[7213]),
			.S(gen[7214]),
			.SE(gen[7215]),

			.SELF(gen[7119]),
			.cell_state(gen[7119])
		); 

/******************* CELL 7120 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7120 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7024]),
			.N(gen[7025]),
			.NE(gen[7026]),

			.O(gen[7119]),
			.E(gen[7121]),

			.SO(gen[7214]),
			.S(gen[7215]),
			.SE(gen[7216]),

			.SELF(gen[7120]),
			.cell_state(gen[7120])
		); 

/******************* CELL 7121 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7121 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7025]),
			.N(gen[7026]),
			.NE(gen[7027]),

			.O(gen[7120]),
			.E(gen[7122]),

			.SO(gen[7215]),
			.S(gen[7216]),
			.SE(gen[7217]),

			.SELF(gen[7121]),
			.cell_state(gen[7121])
		); 

/******************* CELL 7122 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7122 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7026]),
			.N(gen[7027]),
			.NE(gen[7028]),

			.O(gen[7121]),
			.E(gen[7123]),

			.SO(gen[7216]),
			.S(gen[7217]),
			.SE(gen[7218]),

			.SELF(gen[7122]),
			.cell_state(gen[7122])
		); 

/******************* CELL 7123 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7123 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7027]),
			.N(gen[7028]),
			.NE(gen[7029]),

			.O(gen[7122]),
			.E(gen[7124]),

			.SO(gen[7217]),
			.S(gen[7218]),
			.SE(gen[7219]),

			.SELF(gen[7123]),
			.cell_state(gen[7123])
		); 

/******************* CELL 7124 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7124 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7028]),
			.N(gen[7029]),
			.NE(gen[7028]),

			.O(gen[7123]),
			.E(gen[7123]),

			.SO(gen[7218]),
			.S(gen[7219]),
			.SE(gen[7218]),

			.SELF(gen[7124]),
			.cell_state(gen[7124])
		); 

/******************* CELL 7125 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7125 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7031]),
			.N(gen[7030]),
			.NE(gen[7031]),

			.O(gen[7126]),
			.E(gen[7126]),

			.SO(gen[7221]),
			.S(gen[7220]),
			.SE(gen[7221]),

			.SELF(gen[7125]),
			.cell_state(gen[7125])
		); 

/******************* CELL 7126 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7126 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7030]),
			.N(gen[7031]),
			.NE(gen[7032]),

			.O(gen[7125]),
			.E(gen[7127]),

			.SO(gen[7220]),
			.S(gen[7221]),
			.SE(gen[7222]),

			.SELF(gen[7126]),
			.cell_state(gen[7126])
		); 

/******************* CELL 7127 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7127 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7031]),
			.N(gen[7032]),
			.NE(gen[7033]),

			.O(gen[7126]),
			.E(gen[7128]),

			.SO(gen[7221]),
			.S(gen[7222]),
			.SE(gen[7223]),

			.SELF(gen[7127]),
			.cell_state(gen[7127])
		); 

/******************* CELL 7128 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7128 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7032]),
			.N(gen[7033]),
			.NE(gen[7034]),

			.O(gen[7127]),
			.E(gen[7129]),

			.SO(gen[7222]),
			.S(gen[7223]),
			.SE(gen[7224]),

			.SELF(gen[7128]),
			.cell_state(gen[7128])
		); 

/******************* CELL 7129 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7129 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7033]),
			.N(gen[7034]),
			.NE(gen[7035]),

			.O(gen[7128]),
			.E(gen[7130]),

			.SO(gen[7223]),
			.S(gen[7224]),
			.SE(gen[7225]),

			.SELF(gen[7129]),
			.cell_state(gen[7129])
		); 

/******************* CELL 7130 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7130 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7034]),
			.N(gen[7035]),
			.NE(gen[7036]),

			.O(gen[7129]),
			.E(gen[7131]),

			.SO(gen[7224]),
			.S(gen[7225]),
			.SE(gen[7226]),

			.SELF(gen[7130]),
			.cell_state(gen[7130])
		); 

/******************* CELL 7131 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7131 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7035]),
			.N(gen[7036]),
			.NE(gen[7037]),

			.O(gen[7130]),
			.E(gen[7132]),

			.SO(gen[7225]),
			.S(gen[7226]),
			.SE(gen[7227]),

			.SELF(gen[7131]),
			.cell_state(gen[7131])
		); 

/******************* CELL 7132 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7132 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7036]),
			.N(gen[7037]),
			.NE(gen[7038]),

			.O(gen[7131]),
			.E(gen[7133]),

			.SO(gen[7226]),
			.S(gen[7227]),
			.SE(gen[7228]),

			.SELF(gen[7132]),
			.cell_state(gen[7132])
		); 

/******************* CELL 7133 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7133 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7037]),
			.N(gen[7038]),
			.NE(gen[7039]),

			.O(gen[7132]),
			.E(gen[7134]),

			.SO(gen[7227]),
			.S(gen[7228]),
			.SE(gen[7229]),

			.SELF(gen[7133]),
			.cell_state(gen[7133])
		); 

/******************* CELL 7134 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7134 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7038]),
			.N(gen[7039]),
			.NE(gen[7040]),

			.O(gen[7133]),
			.E(gen[7135]),

			.SO(gen[7228]),
			.S(gen[7229]),
			.SE(gen[7230]),

			.SELF(gen[7134]),
			.cell_state(gen[7134])
		); 

/******************* CELL 7135 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7135 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7039]),
			.N(gen[7040]),
			.NE(gen[7041]),

			.O(gen[7134]),
			.E(gen[7136]),

			.SO(gen[7229]),
			.S(gen[7230]),
			.SE(gen[7231]),

			.SELF(gen[7135]),
			.cell_state(gen[7135])
		); 

/******************* CELL 7136 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7136 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7040]),
			.N(gen[7041]),
			.NE(gen[7042]),

			.O(gen[7135]),
			.E(gen[7137]),

			.SO(gen[7230]),
			.S(gen[7231]),
			.SE(gen[7232]),

			.SELF(gen[7136]),
			.cell_state(gen[7136])
		); 

/******************* CELL 7137 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7137 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7041]),
			.N(gen[7042]),
			.NE(gen[7043]),

			.O(gen[7136]),
			.E(gen[7138]),

			.SO(gen[7231]),
			.S(gen[7232]),
			.SE(gen[7233]),

			.SELF(gen[7137]),
			.cell_state(gen[7137])
		); 

/******************* CELL 7138 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7138 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7042]),
			.N(gen[7043]),
			.NE(gen[7044]),

			.O(gen[7137]),
			.E(gen[7139]),

			.SO(gen[7232]),
			.S(gen[7233]),
			.SE(gen[7234]),

			.SELF(gen[7138]),
			.cell_state(gen[7138])
		); 

/******************* CELL 7139 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7139 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7043]),
			.N(gen[7044]),
			.NE(gen[7045]),

			.O(gen[7138]),
			.E(gen[7140]),

			.SO(gen[7233]),
			.S(gen[7234]),
			.SE(gen[7235]),

			.SELF(gen[7139]),
			.cell_state(gen[7139])
		); 

/******************* CELL 7140 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7140 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7044]),
			.N(gen[7045]),
			.NE(gen[7046]),

			.O(gen[7139]),
			.E(gen[7141]),

			.SO(gen[7234]),
			.S(gen[7235]),
			.SE(gen[7236]),

			.SELF(gen[7140]),
			.cell_state(gen[7140])
		); 

/******************* CELL 7141 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7141 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7045]),
			.N(gen[7046]),
			.NE(gen[7047]),

			.O(gen[7140]),
			.E(gen[7142]),

			.SO(gen[7235]),
			.S(gen[7236]),
			.SE(gen[7237]),

			.SELF(gen[7141]),
			.cell_state(gen[7141])
		); 

/******************* CELL 7142 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7142 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7046]),
			.N(gen[7047]),
			.NE(gen[7048]),

			.O(gen[7141]),
			.E(gen[7143]),

			.SO(gen[7236]),
			.S(gen[7237]),
			.SE(gen[7238]),

			.SELF(gen[7142]),
			.cell_state(gen[7142])
		); 

/******************* CELL 7143 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7143 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7047]),
			.N(gen[7048]),
			.NE(gen[7049]),

			.O(gen[7142]),
			.E(gen[7144]),

			.SO(gen[7237]),
			.S(gen[7238]),
			.SE(gen[7239]),

			.SELF(gen[7143]),
			.cell_state(gen[7143])
		); 

/******************* CELL 7144 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7144 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7048]),
			.N(gen[7049]),
			.NE(gen[7050]),

			.O(gen[7143]),
			.E(gen[7145]),

			.SO(gen[7238]),
			.S(gen[7239]),
			.SE(gen[7240]),

			.SELF(gen[7144]),
			.cell_state(gen[7144])
		); 

/******************* CELL 7145 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7145 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7049]),
			.N(gen[7050]),
			.NE(gen[7051]),

			.O(gen[7144]),
			.E(gen[7146]),

			.SO(gen[7239]),
			.S(gen[7240]),
			.SE(gen[7241]),

			.SELF(gen[7145]),
			.cell_state(gen[7145])
		); 

/******************* CELL 7146 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7146 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7050]),
			.N(gen[7051]),
			.NE(gen[7052]),

			.O(gen[7145]),
			.E(gen[7147]),

			.SO(gen[7240]),
			.S(gen[7241]),
			.SE(gen[7242]),

			.SELF(gen[7146]),
			.cell_state(gen[7146])
		); 

/******************* CELL 7147 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7147 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7051]),
			.N(gen[7052]),
			.NE(gen[7053]),

			.O(gen[7146]),
			.E(gen[7148]),

			.SO(gen[7241]),
			.S(gen[7242]),
			.SE(gen[7243]),

			.SELF(gen[7147]),
			.cell_state(gen[7147])
		); 

/******************* CELL 7148 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7148 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7052]),
			.N(gen[7053]),
			.NE(gen[7054]),

			.O(gen[7147]),
			.E(gen[7149]),

			.SO(gen[7242]),
			.S(gen[7243]),
			.SE(gen[7244]),

			.SELF(gen[7148]),
			.cell_state(gen[7148])
		); 

/******************* CELL 7149 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7149 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7053]),
			.N(gen[7054]),
			.NE(gen[7055]),

			.O(gen[7148]),
			.E(gen[7150]),

			.SO(gen[7243]),
			.S(gen[7244]),
			.SE(gen[7245]),

			.SELF(gen[7149]),
			.cell_state(gen[7149])
		); 

/******************* CELL 7150 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7150 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7054]),
			.N(gen[7055]),
			.NE(gen[7056]),

			.O(gen[7149]),
			.E(gen[7151]),

			.SO(gen[7244]),
			.S(gen[7245]),
			.SE(gen[7246]),

			.SELF(gen[7150]),
			.cell_state(gen[7150])
		); 

/******************* CELL 7151 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7151 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7055]),
			.N(gen[7056]),
			.NE(gen[7057]),

			.O(gen[7150]),
			.E(gen[7152]),

			.SO(gen[7245]),
			.S(gen[7246]),
			.SE(gen[7247]),

			.SELF(gen[7151]),
			.cell_state(gen[7151])
		); 

/******************* CELL 7152 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7152 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7056]),
			.N(gen[7057]),
			.NE(gen[7058]),

			.O(gen[7151]),
			.E(gen[7153]),

			.SO(gen[7246]),
			.S(gen[7247]),
			.SE(gen[7248]),

			.SELF(gen[7152]),
			.cell_state(gen[7152])
		); 

/******************* CELL 7153 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7153 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7057]),
			.N(gen[7058]),
			.NE(gen[7059]),

			.O(gen[7152]),
			.E(gen[7154]),

			.SO(gen[7247]),
			.S(gen[7248]),
			.SE(gen[7249]),

			.SELF(gen[7153]),
			.cell_state(gen[7153])
		); 

/******************* CELL 7154 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7154 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7058]),
			.N(gen[7059]),
			.NE(gen[7060]),

			.O(gen[7153]),
			.E(gen[7155]),

			.SO(gen[7248]),
			.S(gen[7249]),
			.SE(gen[7250]),

			.SELF(gen[7154]),
			.cell_state(gen[7154])
		); 

/******************* CELL 7155 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7155 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7059]),
			.N(gen[7060]),
			.NE(gen[7061]),

			.O(gen[7154]),
			.E(gen[7156]),

			.SO(gen[7249]),
			.S(gen[7250]),
			.SE(gen[7251]),

			.SELF(gen[7155]),
			.cell_state(gen[7155])
		); 

/******************* CELL 7156 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7156 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7060]),
			.N(gen[7061]),
			.NE(gen[7062]),

			.O(gen[7155]),
			.E(gen[7157]),

			.SO(gen[7250]),
			.S(gen[7251]),
			.SE(gen[7252]),

			.SELF(gen[7156]),
			.cell_state(gen[7156])
		); 

/******************* CELL 7157 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7157 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7061]),
			.N(gen[7062]),
			.NE(gen[7063]),

			.O(gen[7156]),
			.E(gen[7158]),

			.SO(gen[7251]),
			.S(gen[7252]),
			.SE(gen[7253]),

			.SELF(gen[7157]),
			.cell_state(gen[7157])
		); 

/******************* CELL 7158 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7158 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7062]),
			.N(gen[7063]),
			.NE(gen[7064]),

			.O(gen[7157]),
			.E(gen[7159]),

			.SO(gen[7252]),
			.S(gen[7253]),
			.SE(gen[7254]),

			.SELF(gen[7158]),
			.cell_state(gen[7158])
		); 

/******************* CELL 7159 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7159 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7063]),
			.N(gen[7064]),
			.NE(gen[7065]),

			.O(gen[7158]),
			.E(gen[7160]),

			.SO(gen[7253]),
			.S(gen[7254]),
			.SE(gen[7255]),

			.SELF(gen[7159]),
			.cell_state(gen[7159])
		); 

/******************* CELL 7160 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7160 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7064]),
			.N(gen[7065]),
			.NE(gen[7066]),

			.O(gen[7159]),
			.E(gen[7161]),

			.SO(gen[7254]),
			.S(gen[7255]),
			.SE(gen[7256]),

			.SELF(gen[7160]),
			.cell_state(gen[7160])
		); 

/******************* CELL 7161 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7161 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7065]),
			.N(gen[7066]),
			.NE(gen[7067]),

			.O(gen[7160]),
			.E(gen[7162]),

			.SO(gen[7255]),
			.S(gen[7256]),
			.SE(gen[7257]),

			.SELF(gen[7161]),
			.cell_state(gen[7161])
		); 

/******************* CELL 7162 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7162 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7066]),
			.N(gen[7067]),
			.NE(gen[7068]),

			.O(gen[7161]),
			.E(gen[7163]),

			.SO(gen[7256]),
			.S(gen[7257]),
			.SE(gen[7258]),

			.SELF(gen[7162]),
			.cell_state(gen[7162])
		); 

/******************* CELL 7163 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7163 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7067]),
			.N(gen[7068]),
			.NE(gen[7069]),

			.O(gen[7162]),
			.E(gen[7164]),

			.SO(gen[7257]),
			.S(gen[7258]),
			.SE(gen[7259]),

			.SELF(gen[7163]),
			.cell_state(gen[7163])
		); 

/******************* CELL 7164 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7164 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7068]),
			.N(gen[7069]),
			.NE(gen[7070]),

			.O(gen[7163]),
			.E(gen[7165]),

			.SO(gen[7258]),
			.S(gen[7259]),
			.SE(gen[7260]),

			.SELF(gen[7164]),
			.cell_state(gen[7164])
		); 

/******************* CELL 7165 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7165 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7069]),
			.N(gen[7070]),
			.NE(gen[7071]),

			.O(gen[7164]),
			.E(gen[7166]),

			.SO(gen[7259]),
			.S(gen[7260]),
			.SE(gen[7261]),

			.SELF(gen[7165]),
			.cell_state(gen[7165])
		); 

/******************* CELL 7166 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7166 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7070]),
			.N(gen[7071]),
			.NE(gen[7072]),

			.O(gen[7165]),
			.E(gen[7167]),

			.SO(gen[7260]),
			.S(gen[7261]),
			.SE(gen[7262]),

			.SELF(gen[7166]),
			.cell_state(gen[7166])
		); 

/******************* CELL 7167 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7167 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7071]),
			.N(gen[7072]),
			.NE(gen[7073]),

			.O(gen[7166]),
			.E(gen[7168]),

			.SO(gen[7261]),
			.S(gen[7262]),
			.SE(gen[7263]),

			.SELF(gen[7167]),
			.cell_state(gen[7167])
		); 

/******************* CELL 7168 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7168 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7072]),
			.N(gen[7073]),
			.NE(gen[7074]),

			.O(gen[7167]),
			.E(gen[7169]),

			.SO(gen[7262]),
			.S(gen[7263]),
			.SE(gen[7264]),

			.SELF(gen[7168]),
			.cell_state(gen[7168])
		); 

/******************* CELL 7169 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7169 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7073]),
			.N(gen[7074]),
			.NE(gen[7075]),

			.O(gen[7168]),
			.E(gen[7170]),

			.SO(gen[7263]),
			.S(gen[7264]),
			.SE(gen[7265]),

			.SELF(gen[7169]),
			.cell_state(gen[7169])
		); 

/******************* CELL 7170 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7170 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7074]),
			.N(gen[7075]),
			.NE(gen[7076]),

			.O(gen[7169]),
			.E(gen[7171]),

			.SO(gen[7264]),
			.S(gen[7265]),
			.SE(gen[7266]),

			.SELF(gen[7170]),
			.cell_state(gen[7170])
		); 

/******************* CELL 7171 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7171 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7075]),
			.N(gen[7076]),
			.NE(gen[7077]),

			.O(gen[7170]),
			.E(gen[7172]),

			.SO(gen[7265]),
			.S(gen[7266]),
			.SE(gen[7267]),

			.SELF(gen[7171]),
			.cell_state(gen[7171])
		); 

/******************* CELL 7172 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7172 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7076]),
			.N(gen[7077]),
			.NE(gen[7078]),

			.O(gen[7171]),
			.E(gen[7173]),

			.SO(gen[7266]),
			.S(gen[7267]),
			.SE(gen[7268]),

			.SELF(gen[7172]),
			.cell_state(gen[7172])
		); 

/******************* CELL 7173 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7173 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7077]),
			.N(gen[7078]),
			.NE(gen[7079]),

			.O(gen[7172]),
			.E(gen[7174]),

			.SO(gen[7267]),
			.S(gen[7268]),
			.SE(gen[7269]),

			.SELF(gen[7173]),
			.cell_state(gen[7173])
		); 

/******************* CELL 7174 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7174 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7078]),
			.N(gen[7079]),
			.NE(gen[7080]),

			.O(gen[7173]),
			.E(gen[7175]),

			.SO(gen[7268]),
			.S(gen[7269]),
			.SE(gen[7270]),

			.SELF(gen[7174]),
			.cell_state(gen[7174])
		); 

/******************* CELL 7175 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7175 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7079]),
			.N(gen[7080]),
			.NE(gen[7081]),

			.O(gen[7174]),
			.E(gen[7176]),

			.SO(gen[7269]),
			.S(gen[7270]),
			.SE(gen[7271]),

			.SELF(gen[7175]),
			.cell_state(gen[7175])
		); 

/******************* CELL 7176 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7176 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7080]),
			.N(gen[7081]),
			.NE(gen[7082]),

			.O(gen[7175]),
			.E(gen[7177]),

			.SO(gen[7270]),
			.S(gen[7271]),
			.SE(gen[7272]),

			.SELF(gen[7176]),
			.cell_state(gen[7176])
		); 

/******************* CELL 7177 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7177 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7081]),
			.N(gen[7082]),
			.NE(gen[7083]),

			.O(gen[7176]),
			.E(gen[7178]),

			.SO(gen[7271]),
			.S(gen[7272]),
			.SE(gen[7273]),

			.SELF(gen[7177]),
			.cell_state(gen[7177])
		); 

/******************* CELL 7178 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7178 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7082]),
			.N(gen[7083]),
			.NE(gen[7084]),

			.O(gen[7177]),
			.E(gen[7179]),

			.SO(gen[7272]),
			.S(gen[7273]),
			.SE(gen[7274]),

			.SELF(gen[7178]),
			.cell_state(gen[7178])
		); 

/******************* CELL 7179 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7179 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7083]),
			.N(gen[7084]),
			.NE(gen[7085]),

			.O(gen[7178]),
			.E(gen[7180]),

			.SO(gen[7273]),
			.S(gen[7274]),
			.SE(gen[7275]),

			.SELF(gen[7179]),
			.cell_state(gen[7179])
		); 

/******************* CELL 7180 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7180 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7084]),
			.N(gen[7085]),
			.NE(gen[7086]),

			.O(gen[7179]),
			.E(gen[7181]),

			.SO(gen[7274]),
			.S(gen[7275]),
			.SE(gen[7276]),

			.SELF(gen[7180]),
			.cell_state(gen[7180])
		); 

/******************* CELL 7181 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7181 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7085]),
			.N(gen[7086]),
			.NE(gen[7087]),

			.O(gen[7180]),
			.E(gen[7182]),

			.SO(gen[7275]),
			.S(gen[7276]),
			.SE(gen[7277]),

			.SELF(gen[7181]),
			.cell_state(gen[7181])
		); 

/******************* CELL 7182 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7182 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7086]),
			.N(gen[7087]),
			.NE(gen[7088]),

			.O(gen[7181]),
			.E(gen[7183]),

			.SO(gen[7276]),
			.S(gen[7277]),
			.SE(gen[7278]),

			.SELF(gen[7182]),
			.cell_state(gen[7182])
		); 

/******************* CELL 7183 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7183 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7087]),
			.N(gen[7088]),
			.NE(gen[7089]),

			.O(gen[7182]),
			.E(gen[7184]),

			.SO(gen[7277]),
			.S(gen[7278]),
			.SE(gen[7279]),

			.SELF(gen[7183]),
			.cell_state(gen[7183])
		); 

/******************* CELL 7184 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7184 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7088]),
			.N(gen[7089]),
			.NE(gen[7090]),

			.O(gen[7183]),
			.E(gen[7185]),

			.SO(gen[7278]),
			.S(gen[7279]),
			.SE(gen[7280]),

			.SELF(gen[7184]),
			.cell_state(gen[7184])
		); 

/******************* CELL 7185 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7185 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7089]),
			.N(gen[7090]),
			.NE(gen[7091]),

			.O(gen[7184]),
			.E(gen[7186]),

			.SO(gen[7279]),
			.S(gen[7280]),
			.SE(gen[7281]),

			.SELF(gen[7185]),
			.cell_state(gen[7185])
		); 

/******************* CELL 7186 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7186 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7090]),
			.N(gen[7091]),
			.NE(gen[7092]),

			.O(gen[7185]),
			.E(gen[7187]),

			.SO(gen[7280]),
			.S(gen[7281]),
			.SE(gen[7282]),

			.SELF(gen[7186]),
			.cell_state(gen[7186])
		); 

/******************* CELL 7187 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7187 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7091]),
			.N(gen[7092]),
			.NE(gen[7093]),

			.O(gen[7186]),
			.E(gen[7188]),

			.SO(gen[7281]),
			.S(gen[7282]),
			.SE(gen[7283]),

			.SELF(gen[7187]),
			.cell_state(gen[7187])
		); 

/******************* CELL 7188 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7188 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7092]),
			.N(gen[7093]),
			.NE(gen[7094]),

			.O(gen[7187]),
			.E(gen[7189]),

			.SO(gen[7282]),
			.S(gen[7283]),
			.SE(gen[7284]),

			.SELF(gen[7188]),
			.cell_state(gen[7188])
		); 

/******************* CELL 7189 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7189 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7093]),
			.N(gen[7094]),
			.NE(gen[7095]),

			.O(gen[7188]),
			.E(gen[7190]),

			.SO(gen[7283]),
			.S(gen[7284]),
			.SE(gen[7285]),

			.SELF(gen[7189]),
			.cell_state(gen[7189])
		); 

/******************* CELL 7190 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7190 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7094]),
			.N(gen[7095]),
			.NE(gen[7096]),

			.O(gen[7189]),
			.E(gen[7191]),

			.SO(gen[7284]),
			.S(gen[7285]),
			.SE(gen[7286]),

			.SELF(gen[7190]),
			.cell_state(gen[7190])
		); 

/******************* CELL 7191 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7191 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7095]),
			.N(gen[7096]),
			.NE(gen[7097]),

			.O(gen[7190]),
			.E(gen[7192]),

			.SO(gen[7285]),
			.S(gen[7286]),
			.SE(gen[7287]),

			.SELF(gen[7191]),
			.cell_state(gen[7191])
		); 

/******************* CELL 7192 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7192 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7096]),
			.N(gen[7097]),
			.NE(gen[7098]),

			.O(gen[7191]),
			.E(gen[7193]),

			.SO(gen[7286]),
			.S(gen[7287]),
			.SE(gen[7288]),

			.SELF(gen[7192]),
			.cell_state(gen[7192])
		); 

/******************* CELL 7193 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7193 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7097]),
			.N(gen[7098]),
			.NE(gen[7099]),

			.O(gen[7192]),
			.E(gen[7194]),

			.SO(gen[7287]),
			.S(gen[7288]),
			.SE(gen[7289]),

			.SELF(gen[7193]),
			.cell_state(gen[7193])
		); 

/******************* CELL 7194 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7194 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7098]),
			.N(gen[7099]),
			.NE(gen[7100]),

			.O(gen[7193]),
			.E(gen[7195]),

			.SO(gen[7288]),
			.S(gen[7289]),
			.SE(gen[7290]),

			.SELF(gen[7194]),
			.cell_state(gen[7194])
		); 

/******************* CELL 7195 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7195 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7099]),
			.N(gen[7100]),
			.NE(gen[7101]),

			.O(gen[7194]),
			.E(gen[7196]),

			.SO(gen[7289]),
			.S(gen[7290]),
			.SE(gen[7291]),

			.SELF(gen[7195]),
			.cell_state(gen[7195])
		); 

/******************* CELL 7196 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7196 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7100]),
			.N(gen[7101]),
			.NE(gen[7102]),

			.O(gen[7195]),
			.E(gen[7197]),

			.SO(gen[7290]),
			.S(gen[7291]),
			.SE(gen[7292]),

			.SELF(gen[7196]),
			.cell_state(gen[7196])
		); 

/******************* CELL 7197 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7197 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7101]),
			.N(gen[7102]),
			.NE(gen[7103]),

			.O(gen[7196]),
			.E(gen[7198]),

			.SO(gen[7291]),
			.S(gen[7292]),
			.SE(gen[7293]),

			.SELF(gen[7197]),
			.cell_state(gen[7197])
		); 

/******************* CELL 7198 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7198 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7102]),
			.N(gen[7103]),
			.NE(gen[7104]),

			.O(gen[7197]),
			.E(gen[7199]),

			.SO(gen[7292]),
			.S(gen[7293]),
			.SE(gen[7294]),

			.SELF(gen[7198]),
			.cell_state(gen[7198])
		); 

/******************* CELL 7199 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7199 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7103]),
			.N(gen[7104]),
			.NE(gen[7105]),

			.O(gen[7198]),
			.E(gen[7200]),

			.SO(gen[7293]),
			.S(gen[7294]),
			.SE(gen[7295]),

			.SELF(gen[7199]),
			.cell_state(gen[7199])
		); 

/******************* CELL 7200 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7200 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7104]),
			.N(gen[7105]),
			.NE(gen[7106]),

			.O(gen[7199]),
			.E(gen[7201]),

			.SO(gen[7294]),
			.S(gen[7295]),
			.SE(gen[7296]),

			.SELF(gen[7200]),
			.cell_state(gen[7200])
		); 

/******************* CELL 7201 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7201 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7105]),
			.N(gen[7106]),
			.NE(gen[7107]),

			.O(gen[7200]),
			.E(gen[7202]),

			.SO(gen[7295]),
			.S(gen[7296]),
			.SE(gen[7297]),

			.SELF(gen[7201]),
			.cell_state(gen[7201])
		); 

/******************* CELL 7202 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7202 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7106]),
			.N(gen[7107]),
			.NE(gen[7108]),

			.O(gen[7201]),
			.E(gen[7203]),

			.SO(gen[7296]),
			.S(gen[7297]),
			.SE(gen[7298]),

			.SELF(gen[7202]),
			.cell_state(gen[7202])
		); 

/******************* CELL 7203 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7203 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7107]),
			.N(gen[7108]),
			.NE(gen[7109]),

			.O(gen[7202]),
			.E(gen[7204]),

			.SO(gen[7297]),
			.S(gen[7298]),
			.SE(gen[7299]),

			.SELF(gen[7203]),
			.cell_state(gen[7203])
		); 

/******************* CELL 7204 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7204 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7108]),
			.N(gen[7109]),
			.NE(gen[7110]),

			.O(gen[7203]),
			.E(gen[7205]),

			.SO(gen[7298]),
			.S(gen[7299]),
			.SE(gen[7300]),

			.SELF(gen[7204]),
			.cell_state(gen[7204])
		); 

/******************* CELL 7205 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7205 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7109]),
			.N(gen[7110]),
			.NE(gen[7111]),

			.O(gen[7204]),
			.E(gen[7206]),

			.SO(gen[7299]),
			.S(gen[7300]),
			.SE(gen[7301]),

			.SELF(gen[7205]),
			.cell_state(gen[7205])
		); 

/******************* CELL 7206 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7206 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7110]),
			.N(gen[7111]),
			.NE(gen[7112]),

			.O(gen[7205]),
			.E(gen[7207]),

			.SO(gen[7300]),
			.S(gen[7301]),
			.SE(gen[7302]),

			.SELF(gen[7206]),
			.cell_state(gen[7206])
		); 

/******************* CELL 7207 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7207 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7111]),
			.N(gen[7112]),
			.NE(gen[7113]),

			.O(gen[7206]),
			.E(gen[7208]),

			.SO(gen[7301]),
			.S(gen[7302]),
			.SE(gen[7303]),

			.SELF(gen[7207]),
			.cell_state(gen[7207])
		); 

/******************* CELL 7208 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7208 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7112]),
			.N(gen[7113]),
			.NE(gen[7114]),

			.O(gen[7207]),
			.E(gen[7209]),

			.SO(gen[7302]),
			.S(gen[7303]),
			.SE(gen[7304]),

			.SELF(gen[7208]),
			.cell_state(gen[7208])
		); 

/******************* CELL 7209 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7209 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7113]),
			.N(gen[7114]),
			.NE(gen[7115]),

			.O(gen[7208]),
			.E(gen[7210]),

			.SO(gen[7303]),
			.S(gen[7304]),
			.SE(gen[7305]),

			.SELF(gen[7209]),
			.cell_state(gen[7209])
		); 

/******************* CELL 7210 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7210 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7114]),
			.N(gen[7115]),
			.NE(gen[7116]),

			.O(gen[7209]),
			.E(gen[7211]),

			.SO(gen[7304]),
			.S(gen[7305]),
			.SE(gen[7306]),

			.SELF(gen[7210]),
			.cell_state(gen[7210])
		); 

/******************* CELL 7211 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7211 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7115]),
			.N(gen[7116]),
			.NE(gen[7117]),

			.O(gen[7210]),
			.E(gen[7212]),

			.SO(gen[7305]),
			.S(gen[7306]),
			.SE(gen[7307]),

			.SELF(gen[7211]),
			.cell_state(gen[7211])
		); 

/******************* CELL 7212 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7212 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7116]),
			.N(gen[7117]),
			.NE(gen[7118]),

			.O(gen[7211]),
			.E(gen[7213]),

			.SO(gen[7306]),
			.S(gen[7307]),
			.SE(gen[7308]),

			.SELF(gen[7212]),
			.cell_state(gen[7212])
		); 

/******************* CELL 7213 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7213 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7117]),
			.N(gen[7118]),
			.NE(gen[7119]),

			.O(gen[7212]),
			.E(gen[7214]),

			.SO(gen[7307]),
			.S(gen[7308]),
			.SE(gen[7309]),

			.SELF(gen[7213]),
			.cell_state(gen[7213])
		); 

/******************* CELL 7214 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7214 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7118]),
			.N(gen[7119]),
			.NE(gen[7120]),

			.O(gen[7213]),
			.E(gen[7215]),

			.SO(gen[7308]),
			.S(gen[7309]),
			.SE(gen[7310]),

			.SELF(gen[7214]),
			.cell_state(gen[7214])
		); 

/******************* CELL 7215 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7215 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7119]),
			.N(gen[7120]),
			.NE(gen[7121]),

			.O(gen[7214]),
			.E(gen[7216]),

			.SO(gen[7309]),
			.S(gen[7310]),
			.SE(gen[7311]),

			.SELF(gen[7215]),
			.cell_state(gen[7215])
		); 

/******************* CELL 7216 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7216 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7120]),
			.N(gen[7121]),
			.NE(gen[7122]),

			.O(gen[7215]),
			.E(gen[7217]),

			.SO(gen[7310]),
			.S(gen[7311]),
			.SE(gen[7312]),

			.SELF(gen[7216]),
			.cell_state(gen[7216])
		); 

/******************* CELL 7217 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7217 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7121]),
			.N(gen[7122]),
			.NE(gen[7123]),

			.O(gen[7216]),
			.E(gen[7218]),

			.SO(gen[7311]),
			.S(gen[7312]),
			.SE(gen[7313]),

			.SELF(gen[7217]),
			.cell_state(gen[7217])
		); 

/******************* CELL 7218 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7218 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7122]),
			.N(gen[7123]),
			.NE(gen[7124]),

			.O(gen[7217]),
			.E(gen[7219]),

			.SO(gen[7312]),
			.S(gen[7313]),
			.SE(gen[7314]),

			.SELF(gen[7218]),
			.cell_state(gen[7218])
		); 

/******************* CELL 7219 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7219 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7123]),
			.N(gen[7124]),
			.NE(gen[7123]),

			.O(gen[7218]),
			.E(gen[7218]),

			.SO(gen[7313]),
			.S(gen[7314]),
			.SE(gen[7313]),

			.SELF(gen[7219]),
			.cell_state(gen[7219])
		); 

/******************* CELL 7220 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7220 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7126]),
			.N(gen[7125]),
			.NE(gen[7126]),

			.O(gen[7221]),
			.E(gen[7221]),

			.SO(gen[7316]),
			.S(gen[7315]),
			.SE(gen[7316]),

			.SELF(gen[7220]),
			.cell_state(gen[7220])
		); 

/******************* CELL 7221 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7221 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7125]),
			.N(gen[7126]),
			.NE(gen[7127]),

			.O(gen[7220]),
			.E(gen[7222]),

			.SO(gen[7315]),
			.S(gen[7316]),
			.SE(gen[7317]),

			.SELF(gen[7221]),
			.cell_state(gen[7221])
		); 

/******************* CELL 7222 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7222 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7126]),
			.N(gen[7127]),
			.NE(gen[7128]),

			.O(gen[7221]),
			.E(gen[7223]),

			.SO(gen[7316]),
			.S(gen[7317]),
			.SE(gen[7318]),

			.SELF(gen[7222]),
			.cell_state(gen[7222])
		); 

/******************* CELL 7223 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7223 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7127]),
			.N(gen[7128]),
			.NE(gen[7129]),

			.O(gen[7222]),
			.E(gen[7224]),

			.SO(gen[7317]),
			.S(gen[7318]),
			.SE(gen[7319]),

			.SELF(gen[7223]),
			.cell_state(gen[7223])
		); 

/******************* CELL 7224 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7224 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7128]),
			.N(gen[7129]),
			.NE(gen[7130]),

			.O(gen[7223]),
			.E(gen[7225]),

			.SO(gen[7318]),
			.S(gen[7319]),
			.SE(gen[7320]),

			.SELF(gen[7224]),
			.cell_state(gen[7224])
		); 

/******************* CELL 7225 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7225 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7129]),
			.N(gen[7130]),
			.NE(gen[7131]),

			.O(gen[7224]),
			.E(gen[7226]),

			.SO(gen[7319]),
			.S(gen[7320]),
			.SE(gen[7321]),

			.SELF(gen[7225]),
			.cell_state(gen[7225])
		); 

/******************* CELL 7226 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7226 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7130]),
			.N(gen[7131]),
			.NE(gen[7132]),

			.O(gen[7225]),
			.E(gen[7227]),

			.SO(gen[7320]),
			.S(gen[7321]),
			.SE(gen[7322]),

			.SELF(gen[7226]),
			.cell_state(gen[7226])
		); 

/******************* CELL 7227 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7227 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7131]),
			.N(gen[7132]),
			.NE(gen[7133]),

			.O(gen[7226]),
			.E(gen[7228]),

			.SO(gen[7321]),
			.S(gen[7322]),
			.SE(gen[7323]),

			.SELF(gen[7227]),
			.cell_state(gen[7227])
		); 

/******************* CELL 7228 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7228 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7132]),
			.N(gen[7133]),
			.NE(gen[7134]),

			.O(gen[7227]),
			.E(gen[7229]),

			.SO(gen[7322]),
			.S(gen[7323]),
			.SE(gen[7324]),

			.SELF(gen[7228]),
			.cell_state(gen[7228])
		); 

/******************* CELL 7229 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7229 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7133]),
			.N(gen[7134]),
			.NE(gen[7135]),

			.O(gen[7228]),
			.E(gen[7230]),

			.SO(gen[7323]),
			.S(gen[7324]),
			.SE(gen[7325]),

			.SELF(gen[7229]),
			.cell_state(gen[7229])
		); 

/******************* CELL 7230 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7230 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7134]),
			.N(gen[7135]),
			.NE(gen[7136]),

			.O(gen[7229]),
			.E(gen[7231]),

			.SO(gen[7324]),
			.S(gen[7325]),
			.SE(gen[7326]),

			.SELF(gen[7230]),
			.cell_state(gen[7230])
		); 

/******************* CELL 7231 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7231 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7135]),
			.N(gen[7136]),
			.NE(gen[7137]),

			.O(gen[7230]),
			.E(gen[7232]),

			.SO(gen[7325]),
			.S(gen[7326]),
			.SE(gen[7327]),

			.SELF(gen[7231]),
			.cell_state(gen[7231])
		); 

/******************* CELL 7232 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7232 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7136]),
			.N(gen[7137]),
			.NE(gen[7138]),

			.O(gen[7231]),
			.E(gen[7233]),

			.SO(gen[7326]),
			.S(gen[7327]),
			.SE(gen[7328]),

			.SELF(gen[7232]),
			.cell_state(gen[7232])
		); 

/******************* CELL 7233 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7233 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7137]),
			.N(gen[7138]),
			.NE(gen[7139]),

			.O(gen[7232]),
			.E(gen[7234]),

			.SO(gen[7327]),
			.S(gen[7328]),
			.SE(gen[7329]),

			.SELF(gen[7233]),
			.cell_state(gen[7233])
		); 

/******************* CELL 7234 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7234 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7138]),
			.N(gen[7139]),
			.NE(gen[7140]),

			.O(gen[7233]),
			.E(gen[7235]),

			.SO(gen[7328]),
			.S(gen[7329]),
			.SE(gen[7330]),

			.SELF(gen[7234]),
			.cell_state(gen[7234])
		); 

/******************* CELL 7235 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7235 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7139]),
			.N(gen[7140]),
			.NE(gen[7141]),

			.O(gen[7234]),
			.E(gen[7236]),

			.SO(gen[7329]),
			.S(gen[7330]),
			.SE(gen[7331]),

			.SELF(gen[7235]),
			.cell_state(gen[7235])
		); 

/******************* CELL 7236 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7236 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7140]),
			.N(gen[7141]),
			.NE(gen[7142]),

			.O(gen[7235]),
			.E(gen[7237]),

			.SO(gen[7330]),
			.S(gen[7331]),
			.SE(gen[7332]),

			.SELF(gen[7236]),
			.cell_state(gen[7236])
		); 

/******************* CELL 7237 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7237 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7141]),
			.N(gen[7142]),
			.NE(gen[7143]),

			.O(gen[7236]),
			.E(gen[7238]),

			.SO(gen[7331]),
			.S(gen[7332]),
			.SE(gen[7333]),

			.SELF(gen[7237]),
			.cell_state(gen[7237])
		); 

/******************* CELL 7238 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7238 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7142]),
			.N(gen[7143]),
			.NE(gen[7144]),

			.O(gen[7237]),
			.E(gen[7239]),

			.SO(gen[7332]),
			.S(gen[7333]),
			.SE(gen[7334]),

			.SELF(gen[7238]),
			.cell_state(gen[7238])
		); 

/******************* CELL 7239 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7239 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7143]),
			.N(gen[7144]),
			.NE(gen[7145]),

			.O(gen[7238]),
			.E(gen[7240]),

			.SO(gen[7333]),
			.S(gen[7334]),
			.SE(gen[7335]),

			.SELF(gen[7239]),
			.cell_state(gen[7239])
		); 

/******************* CELL 7240 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7240 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7144]),
			.N(gen[7145]),
			.NE(gen[7146]),

			.O(gen[7239]),
			.E(gen[7241]),

			.SO(gen[7334]),
			.S(gen[7335]),
			.SE(gen[7336]),

			.SELF(gen[7240]),
			.cell_state(gen[7240])
		); 

/******************* CELL 7241 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7241 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7145]),
			.N(gen[7146]),
			.NE(gen[7147]),

			.O(gen[7240]),
			.E(gen[7242]),

			.SO(gen[7335]),
			.S(gen[7336]),
			.SE(gen[7337]),

			.SELF(gen[7241]),
			.cell_state(gen[7241])
		); 

/******************* CELL 7242 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7242 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7146]),
			.N(gen[7147]),
			.NE(gen[7148]),

			.O(gen[7241]),
			.E(gen[7243]),

			.SO(gen[7336]),
			.S(gen[7337]),
			.SE(gen[7338]),

			.SELF(gen[7242]),
			.cell_state(gen[7242])
		); 

/******************* CELL 7243 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7243 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7147]),
			.N(gen[7148]),
			.NE(gen[7149]),

			.O(gen[7242]),
			.E(gen[7244]),

			.SO(gen[7337]),
			.S(gen[7338]),
			.SE(gen[7339]),

			.SELF(gen[7243]),
			.cell_state(gen[7243])
		); 

/******************* CELL 7244 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7244 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7148]),
			.N(gen[7149]),
			.NE(gen[7150]),

			.O(gen[7243]),
			.E(gen[7245]),

			.SO(gen[7338]),
			.S(gen[7339]),
			.SE(gen[7340]),

			.SELF(gen[7244]),
			.cell_state(gen[7244])
		); 

/******************* CELL 7245 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7245 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7149]),
			.N(gen[7150]),
			.NE(gen[7151]),

			.O(gen[7244]),
			.E(gen[7246]),

			.SO(gen[7339]),
			.S(gen[7340]),
			.SE(gen[7341]),

			.SELF(gen[7245]),
			.cell_state(gen[7245])
		); 

/******************* CELL 7246 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7246 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7150]),
			.N(gen[7151]),
			.NE(gen[7152]),

			.O(gen[7245]),
			.E(gen[7247]),

			.SO(gen[7340]),
			.S(gen[7341]),
			.SE(gen[7342]),

			.SELF(gen[7246]),
			.cell_state(gen[7246])
		); 

/******************* CELL 7247 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7247 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7151]),
			.N(gen[7152]),
			.NE(gen[7153]),

			.O(gen[7246]),
			.E(gen[7248]),

			.SO(gen[7341]),
			.S(gen[7342]),
			.SE(gen[7343]),

			.SELF(gen[7247]),
			.cell_state(gen[7247])
		); 

/******************* CELL 7248 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7248 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7152]),
			.N(gen[7153]),
			.NE(gen[7154]),

			.O(gen[7247]),
			.E(gen[7249]),

			.SO(gen[7342]),
			.S(gen[7343]),
			.SE(gen[7344]),

			.SELF(gen[7248]),
			.cell_state(gen[7248])
		); 

/******************* CELL 7249 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7249 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7153]),
			.N(gen[7154]),
			.NE(gen[7155]),

			.O(gen[7248]),
			.E(gen[7250]),

			.SO(gen[7343]),
			.S(gen[7344]),
			.SE(gen[7345]),

			.SELF(gen[7249]),
			.cell_state(gen[7249])
		); 

/******************* CELL 7250 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7250 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7154]),
			.N(gen[7155]),
			.NE(gen[7156]),

			.O(gen[7249]),
			.E(gen[7251]),

			.SO(gen[7344]),
			.S(gen[7345]),
			.SE(gen[7346]),

			.SELF(gen[7250]),
			.cell_state(gen[7250])
		); 

/******************* CELL 7251 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7251 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7155]),
			.N(gen[7156]),
			.NE(gen[7157]),

			.O(gen[7250]),
			.E(gen[7252]),

			.SO(gen[7345]),
			.S(gen[7346]),
			.SE(gen[7347]),

			.SELF(gen[7251]),
			.cell_state(gen[7251])
		); 

/******************* CELL 7252 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7252 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7156]),
			.N(gen[7157]),
			.NE(gen[7158]),

			.O(gen[7251]),
			.E(gen[7253]),

			.SO(gen[7346]),
			.S(gen[7347]),
			.SE(gen[7348]),

			.SELF(gen[7252]),
			.cell_state(gen[7252])
		); 

/******************* CELL 7253 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7253 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7157]),
			.N(gen[7158]),
			.NE(gen[7159]),

			.O(gen[7252]),
			.E(gen[7254]),

			.SO(gen[7347]),
			.S(gen[7348]),
			.SE(gen[7349]),

			.SELF(gen[7253]),
			.cell_state(gen[7253])
		); 

/******************* CELL 7254 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7254 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7158]),
			.N(gen[7159]),
			.NE(gen[7160]),

			.O(gen[7253]),
			.E(gen[7255]),

			.SO(gen[7348]),
			.S(gen[7349]),
			.SE(gen[7350]),

			.SELF(gen[7254]),
			.cell_state(gen[7254])
		); 

/******************* CELL 7255 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7255 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7159]),
			.N(gen[7160]),
			.NE(gen[7161]),

			.O(gen[7254]),
			.E(gen[7256]),

			.SO(gen[7349]),
			.S(gen[7350]),
			.SE(gen[7351]),

			.SELF(gen[7255]),
			.cell_state(gen[7255])
		); 

/******************* CELL 7256 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7256 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7160]),
			.N(gen[7161]),
			.NE(gen[7162]),

			.O(gen[7255]),
			.E(gen[7257]),

			.SO(gen[7350]),
			.S(gen[7351]),
			.SE(gen[7352]),

			.SELF(gen[7256]),
			.cell_state(gen[7256])
		); 

/******************* CELL 7257 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7257 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7161]),
			.N(gen[7162]),
			.NE(gen[7163]),

			.O(gen[7256]),
			.E(gen[7258]),

			.SO(gen[7351]),
			.S(gen[7352]),
			.SE(gen[7353]),

			.SELF(gen[7257]),
			.cell_state(gen[7257])
		); 

/******************* CELL 7258 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7258 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7162]),
			.N(gen[7163]),
			.NE(gen[7164]),

			.O(gen[7257]),
			.E(gen[7259]),

			.SO(gen[7352]),
			.S(gen[7353]),
			.SE(gen[7354]),

			.SELF(gen[7258]),
			.cell_state(gen[7258])
		); 

/******************* CELL 7259 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7259 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7163]),
			.N(gen[7164]),
			.NE(gen[7165]),

			.O(gen[7258]),
			.E(gen[7260]),

			.SO(gen[7353]),
			.S(gen[7354]),
			.SE(gen[7355]),

			.SELF(gen[7259]),
			.cell_state(gen[7259])
		); 

/******************* CELL 7260 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7260 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7164]),
			.N(gen[7165]),
			.NE(gen[7166]),

			.O(gen[7259]),
			.E(gen[7261]),

			.SO(gen[7354]),
			.S(gen[7355]),
			.SE(gen[7356]),

			.SELF(gen[7260]),
			.cell_state(gen[7260])
		); 

/******************* CELL 7261 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7261 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7165]),
			.N(gen[7166]),
			.NE(gen[7167]),

			.O(gen[7260]),
			.E(gen[7262]),

			.SO(gen[7355]),
			.S(gen[7356]),
			.SE(gen[7357]),

			.SELF(gen[7261]),
			.cell_state(gen[7261])
		); 

/******************* CELL 7262 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7262 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7166]),
			.N(gen[7167]),
			.NE(gen[7168]),

			.O(gen[7261]),
			.E(gen[7263]),

			.SO(gen[7356]),
			.S(gen[7357]),
			.SE(gen[7358]),

			.SELF(gen[7262]),
			.cell_state(gen[7262])
		); 

/******************* CELL 7263 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7263 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7167]),
			.N(gen[7168]),
			.NE(gen[7169]),

			.O(gen[7262]),
			.E(gen[7264]),

			.SO(gen[7357]),
			.S(gen[7358]),
			.SE(gen[7359]),

			.SELF(gen[7263]),
			.cell_state(gen[7263])
		); 

/******************* CELL 7264 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7264 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7168]),
			.N(gen[7169]),
			.NE(gen[7170]),

			.O(gen[7263]),
			.E(gen[7265]),

			.SO(gen[7358]),
			.S(gen[7359]),
			.SE(gen[7360]),

			.SELF(gen[7264]),
			.cell_state(gen[7264])
		); 

/******************* CELL 7265 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7265 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7169]),
			.N(gen[7170]),
			.NE(gen[7171]),

			.O(gen[7264]),
			.E(gen[7266]),

			.SO(gen[7359]),
			.S(gen[7360]),
			.SE(gen[7361]),

			.SELF(gen[7265]),
			.cell_state(gen[7265])
		); 

/******************* CELL 7266 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7266 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7170]),
			.N(gen[7171]),
			.NE(gen[7172]),

			.O(gen[7265]),
			.E(gen[7267]),

			.SO(gen[7360]),
			.S(gen[7361]),
			.SE(gen[7362]),

			.SELF(gen[7266]),
			.cell_state(gen[7266])
		); 

/******************* CELL 7267 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7267 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7171]),
			.N(gen[7172]),
			.NE(gen[7173]),

			.O(gen[7266]),
			.E(gen[7268]),

			.SO(gen[7361]),
			.S(gen[7362]),
			.SE(gen[7363]),

			.SELF(gen[7267]),
			.cell_state(gen[7267])
		); 

/******************* CELL 7268 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7268 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7172]),
			.N(gen[7173]),
			.NE(gen[7174]),

			.O(gen[7267]),
			.E(gen[7269]),

			.SO(gen[7362]),
			.S(gen[7363]),
			.SE(gen[7364]),

			.SELF(gen[7268]),
			.cell_state(gen[7268])
		); 

/******************* CELL 7269 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7269 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7173]),
			.N(gen[7174]),
			.NE(gen[7175]),

			.O(gen[7268]),
			.E(gen[7270]),

			.SO(gen[7363]),
			.S(gen[7364]),
			.SE(gen[7365]),

			.SELF(gen[7269]),
			.cell_state(gen[7269])
		); 

/******************* CELL 7270 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7270 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7174]),
			.N(gen[7175]),
			.NE(gen[7176]),

			.O(gen[7269]),
			.E(gen[7271]),

			.SO(gen[7364]),
			.S(gen[7365]),
			.SE(gen[7366]),

			.SELF(gen[7270]),
			.cell_state(gen[7270])
		); 

/******************* CELL 7271 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7271 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7175]),
			.N(gen[7176]),
			.NE(gen[7177]),

			.O(gen[7270]),
			.E(gen[7272]),

			.SO(gen[7365]),
			.S(gen[7366]),
			.SE(gen[7367]),

			.SELF(gen[7271]),
			.cell_state(gen[7271])
		); 

/******************* CELL 7272 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7272 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7176]),
			.N(gen[7177]),
			.NE(gen[7178]),

			.O(gen[7271]),
			.E(gen[7273]),

			.SO(gen[7366]),
			.S(gen[7367]),
			.SE(gen[7368]),

			.SELF(gen[7272]),
			.cell_state(gen[7272])
		); 

/******************* CELL 7273 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7273 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7177]),
			.N(gen[7178]),
			.NE(gen[7179]),

			.O(gen[7272]),
			.E(gen[7274]),

			.SO(gen[7367]),
			.S(gen[7368]),
			.SE(gen[7369]),

			.SELF(gen[7273]),
			.cell_state(gen[7273])
		); 

/******************* CELL 7274 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7274 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7178]),
			.N(gen[7179]),
			.NE(gen[7180]),

			.O(gen[7273]),
			.E(gen[7275]),

			.SO(gen[7368]),
			.S(gen[7369]),
			.SE(gen[7370]),

			.SELF(gen[7274]),
			.cell_state(gen[7274])
		); 

/******************* CELL 7275 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7275 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7179]),
			.N(gen[7180]),
			.NE(gen[7181]),

			.O(gen[7274]),
			.E(gen[7276]),

			.SO(gen[7369]),
			.S(gen[7370]),
			.SE(gen[7371]),

			.SELF(gen[7275]),
			.cell_state(gen[7275])
		); 

/******************* CELL 7276 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7276 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7180]),
			.N(gen[7181]),
			.NE(gen[7182]),

			.O(gen[7275]),
			.E(gen[7277]),

			.SO(gen[7370]),
			.S(gen[7371]),
			.SE(gen[7372]),

			.SELF(gen[7276]),
			.cell_state(gen[7276])
		); 

/******************* CELL 7277 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7277 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7181]),
			.N(gen[7182]),
			.NE(gen[7183]),

			.O(gen[7276]),
			.E(gen[7278]),

			.SO(gen[7371]),
			.S(gen[7372]),
			.SE(gen[7373]),

			.SELF(gen[7277]),
			.cell_state(gen[7277])
		); 

/******************* CELL 7278 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7278 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7182]),
			.N(gen[7183]),
			.NE(gen[7184]),

			.O(gen[7277]),
			.E(gen[7279]),

			.SO(gen[7372]),
			.S(gen[7373]),
			.SE(gen[7374]),

			.SELF(gen[7278]),
			.cell_state(gen[7278])
		); 

/******************* CELL 7279 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7279 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7183]),
			.N(gen[7184]),
			.NE(gen[7185]),

			.O(gen[7278]),
			.E(gen[7280]),

			.SO(gen[7373]),
			.S(gen[7374]),
			.SE(gen[7375]),

			.SELF(gen[7279]),
			.cell_state(gen[7279])
		); 

/******************* CELL 7280 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7280 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7184]),
			.N(gen[7185]),
			.NE(gen[7186]),

			.O(gen[7279]),
			.E(gen[7281]),

			.SO(gen[7374]),
			.S(gen[7375]),
			.SE(gen[7376]),

			.SELF(gen[7280]),
			.cell_state(gen[7280])
		); 

/******************* CELL 7281 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7281 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7185]),
			.N(gen[7186]),
			.NE(gen[7187]),

			.O(gen[7280]),
			.E(gen[7282]),

			.SO(gen[7375]),
			.S(gen[7376]),
			.SE(gen[7377]),

			.SELF(gen[7281]),
			.cell_state(gen[7281])
		); 

/******************* CELL 7282 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7282 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7186]),
			.N(gen[7187]),
			.NE(gen[7188]),

			.O(gen[7281]),
			.E(gen[7283]),

			.SO(gen[7376]),
			.S(gen[7377]),
			.SE(gen[7378]),

			.SELF(gen[7282]),
			.cell_state(gen[7282])
		); 

/******************* CELL 7283 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7283 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7187]),
			.N(gen[7188]),
			.NE(gen[7189]),

			.O(gen[7282]),
			.E(gen[7284]),

			.SO(gen[7377]),
			.S(gen[7378]),
			.SE(gen[7379]),

			.SELF(gen[7283]),
			.cell_state(gen[7283])
		); 

/******************* CELL 7284 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7284 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7188]),
			.N(gen[7189]),
			.NE(gen[7190]),

			.O(gen[7283]),
			.E(gen[7285]),

			.SO(gen[7378]),
			.S(gen[7379]),
			.SE(gen[7380]),

			.SELF(gen[7284]),
			.cell_state(gen[7284])
		); 

/******************* CELL 7285 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7285 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7189]),
			.N(gen[7190]),
			.NE(gen[7191]),

			.O(gen[7284]),
			.E(gen[7286]),

			.SO(gen[7379]),
			.S(gen[7380]),
			.SE(gen[7381]),

			.SELF(gen[7285]),
			.cell_state(gen[7285])
		); 

/******************* CELL 7286 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7286 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7190]),
			.N(gen[7191]),
			.NE(gen[7192]),

			.O(gen[7285]),
			.E(gen[7287]),

			.SO(gen[7380]),
			.S(gen[7381]),
			.SE(gen[7382]),

			.SELF(gen[7286]),
			.cell_state(gen[7286])
		); 

/******************* CELL 7287 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7287 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7191]),
			.N(gen[7192]),
			.NE(gen[7193]),

			.O(gen[7286]),
			.E(gen[7288]),

			.SO(gen[7381]),
			.S(gen[7382]),
			.SE(gen[7383]),

			.SELF(gen[7287]),
			.cell_state(gen[7287])
		); 

/******************* CELL 7288 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7288 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7192]),
			.N(gen[7193]),
			.NE(gen[7194]),

			.O(gen[7287]),
			.E(gen[7289]),

			.SO(gen[7382]),
			.S(gen[7383]),
			.SE(gen[7384]),

			.SELF(gen[7288]),
			.cell_state(gen[7288])
		); 

/******************* CELL 7289 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7289 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7193]),
			.N(gen[7194]),
			.NE(gen[7195]),

			.O(gen[7288]),
			.E(gen[7290]),

			.SO(gen[7383]),
			.S(gen[7384]),
			.SE(gen[7385]),

			.SELF(gen[7289]),
			.cell_state(gen[7289])
		); 

/******************* CELL 7290 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7290 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7194]),
			.N(gen[7195]),
			.NE(gen[7196]),

			.O(gen[7289]),
			.E(gen[7291]),

			.SO(gen[7384]),
			.S(gen[7385]),
			.SE(gen[7386]),

			.SELF(gen[7290]),
			.cell_state(gen[7290])
		); 

/******************* CELL 7291 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7291 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7195]),
			.N(gen[7196]),
			.NE(gen[7197]),

			.O(gen[7290]),
			.E(gen[7292]),

			.SO(gen[7385]),
			.S(gen[7386]),
			.SE(gen[7387]),

			.SELF(gen[7291]),
			.cell_state(gen[7291])
		); 

/******************* CELL 7292 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7292 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7196]),
			.N(gen[7197]),
			.NE(gen[7198]),

			.O(gen[7291]),
			.E(gen[7293]),

			.SO(gen[7386]),
			.S(gen[7387]),
			.SE(gen[7388]),

			.SELF(gen[7292]),
			.cell_state(gen[7292])
		); 

/******************* CELL 7293 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7293 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7197]),
			.N(gen[7198]),
			.NE(gen[7199]),

			.O(gen[7292]),
			.E(gen[7294]),

			.SO(gen[7387]),
			.S(gen[7388]),
			.SE(gen[7389]),

			.SELF(gen[7293]),
			.cell_state(gen[7293])
		); 

/******************* CELL 7294 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7294 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7198]),
			.N(gen[7199]),
			.NE(gen[7200]),

			.O(gen[7293]),
			.E(gen[7295]),

			.SO(gen[7388]),
			.S(gen[7389]),
			.SE(gen[7390]),

			.SELF(gen[7294]),
			.cell_state(gen[7294])
		); 

/******************* CELL 7295 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7295 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7199]),
			.N(gen[7200]),
			.NE(gen[7201]),

			.O(gen[7294]),
			.E(gen[7296]),

			.SO(gen[7389]),
			.S(gen[7390]),
			.SE(gen[7391]),

			.SELF(gen[7295]),
			.cell_state(gen[7295])
		); 

/******************* CELL 7296 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7296 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7200]),
			.N(gen[7201]),
			.NE(gen[7202]),

			.O(gen[7295]),
			.E(gen[7297]),

			.SO(gen[7390]),
			.S(gen[7391]),
			.SE(gen[7392]),

			.SELF(gen[7296]),
			.cell_state(gen[7296])
		); 

/******************* CELL 7297 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7297 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7201]),
			.N(gen[7202]),
			.NE(gen[7203]),

			.O(gen[7296]),
			.E(gen[7298]),

			.SO(gen[7391]),
			.S(gen[7392]),
			.SE(gen[7393]),

			.SELF(gen[7297]),
			.cell_state(gen[7297])
		); 

/******************* CELL 7298 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7298 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7202]),
			.N(gen[7203]),
			.NE(gen[7204]),

			.O(gen[7297]),
			.E(gen[7299]),

			.SO(gen[7392]),
			.S(gen[7393]),
			.SE(gen[7394]),

			.SELF(gen[7298]),
			.cell_state(gen[7298])
		); 

/******************* CELL 7299 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7299 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7203]),
			.N(gen[7204]),
			.NE(gen[7205]),

			.O(gen[7298]),
			.E(gen[7300]),

			.SO(gen[7393]),
			.S(gen[7394]),
			.SE(gen[7395]),

			.SELF(gen[7299]),
			.cell_state(gen[7299])
		); 

/******************* CELL 7300 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7300 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7204]),
			.N(gen[7205]),
			.NE(gen[7206]),

			.O(gen[7299]),
			.E(gen[7301]),

			.SO(gen[7394]),
			.S(gen[7395]),
			.SE(gen[7396]),

			.SELF(gen[7300]),
			.cell_state(gen[7300])
		); 

/******************* CELL 7301 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7301 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7205]),
			.N(gen[7206]),
			.NE(gen[7207]),

			.O(gen[7300]),
			.E(gen[7302]),

			.SO(gen[7395]),
			.S(gen[7396]),
			.SE(gen[7397]),

			.SELF(gen[7301]),
			.cell_state(gen[7301])
		); 

/******************* CELL 7302 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7302 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7206]),
			.N(gen[7207]),
			.NE(gen[7208]),

			.O(gen[7301]),
			.E(gen[7303]),

			.SO(gen[7396]),
			.S(gen[7397]),
			.SE(gen[7398]),

			.SELF(gen[7302]),
			.cell_state(gen[7302])
		); 

/******************* CELL 7303 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7303 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7207]),
			.N(gen[7208]),
			.NE(gen[7209]),

			.O(gen[7302]),
			.E(gen[7304]),

			.SO(gen[7397]),
			.S(gen[7398]),
			.SE(gen[7399]),

			.SELF(gen[7303]),
			.cell_state(gen[7303])
		); 

/******************* CELL 7304 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7304 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7208]),
			.N(gen[7209]),
			.NE(gen[7210]),

			.O(gen[7303]),
			.E(gen[7305]),

			.SO(gen[7398]),
			.S(gen[7399]),
			.SE(gen[7400]),

			.SELF(gen[7304]),
			.cell_state(gen[7304])
		); 

/******************* CELL 7305 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7305 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7209]),
			.N(gen[7210]),
			.NE(gen[7211]),

			.O(gen[7304]),
			.E(gen[7306]),

			.SO(gen[7399]),
			.S(gen[7400]),
			.SE(gen[7401]),

			.SELF(gen[7305]),
			.cell_state(gen[7305])
		); 

/******************* CELL 7306 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7306 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7210]),
			.N(gen[7211]),
			.NE(gen[7212]),

			.O(gen[7305]),
			.E(gen[7307]),

			.SO(gen[7400]),
			.S(gen[7401]),
			.SE(gen[7402]),

			.SELF(gen[7306]),
			.cell_state(gen[7306])
		); 

/******************* CELL 7307 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7307 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7211]),
			.N(gen[7212]),
			.NE(gen[7213]),

			.O(gen[7306]),
			.E(gen[7308]),

			.SO(gen[7401]),
			.S(gen[7402]),
			.SE(gen[7403]),

			.SELF(gen[7307]),
			.cell_state(gen[7307])
		); 

/******************* CELL 7308 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7308 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7212]),
			.N(gen[7213]),
			.NE(gen[7214]),

			.O(gen[7307]),
			.E(gen[7309]),

			.SO(gen[7402]),
			.S(gen[7403]),
			.SE(gen[7404]),

			.SELF(gen[7308]),
			.cell_state(gen[7308])
		); 

/******************* CELL 7309 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7309 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7213]),
			.N(gen[7214]),
			.NE(gen[7215]),

			.O(gen[7308]),
			.E(gen[7310]),

			.SO(gen[7403]),
			.S(gen[7404]),
			.SE(gen[7405]),

			.SELF(gen[7309]),
			.cell_state(gen[7309])
		); 

/******************* CELL 7310 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7310 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7214]),
			.N(gen[7215]),
			.NE(gen[7216]),

			.O(gen[7309]),
			.E(gen[7311]),

			.SO(gen[7404]),
			.S(gen[7405]),
			.SE(gen[7406]),

			.SELF(gen[7310]),
			.cell_state(gen[7310])
		); 

/******************* CELL 7311 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7311 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7215]),
			.N(gen[7216]),
			.NE(gen[7217]),

			.O(gen[7310]),
			.E(gen[7312]),

			.SO(gen[7405]),
			.S(gen[7406]),
			.SE(gen[7407]),

			.SELF(gen[7311]),
			.cell_state(gen[7311])
		); 

/******************* CELL 7312 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7312 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7216]),
			.N(gen[7217]),
			.NE(gen[7218]),

			.O(gen[7311]),
			.E(gen[7313]),

			.SO(gen[7406]),
			.S(gen[7407]),
			.SE(gen[7408]),

			.SELF(gen[7312]),
			.cell_state(gen[7312])
		); 

/******************* CELL 7313 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7313 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7217]),
			.N(gen[7218]),
			.NE(gen[7219]),

			.O(gen[7312]),
			.E(gen[7314]),

			.SO(gen[7407]),
			.S(gen[7408]),
			.SE(gen[7409]),

			.SELF(gen[7313]),
			.cell_state(gen[7313])
		); 

/******************* CELL 7314 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7314 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7218]),
			.N(gen[7219]),
			.NE(gen[7218]),

			.O(gen[7313]),
			.E(gen[7313]),

			.SO(gen[7408]),
			.S(gen[7409]),
			.SE(gen[7408]),

			.SELF(gen[7314]),
			.cell_state(gen[7314])
		); 

/******************* CELL 7315 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7315 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7221]),
			.N(gen[7220]),
			.NE(gen[7221]),

			.O(gen[7316]),
			.E(gen[7316]),

			.SO(gen[7411]),
			.S(gen[7410]),
			.SE(gen[7411]),

			.SELF(gen[7315]),
			.cell_state(gen[7315])
		); 

/******************* CELL 7316 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7316 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7220]),
			.N(gen[7221]),
			.NE(gen[7222]),

			.O(gen[7315]),
			.E(gen[7317]),

			.SO(gen[7410]),
			.S(gen[7411]),
			.SE(gen[7412]),

			.SELF(gen[7316]),
			.cell_state(gen[7316])
		); 

/******************* CELL 7317 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7317 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7221]),
			.N(gen[7222]),
			.NE(gen[7223]),

			.O(gen[7316]),
			.E(gen[7318]),

			.SO(gen[7411]),
			.S(gen[7412]),
			.SE(gen[7413]),

			.SELF(gen[7317]),
			.cell_state(gen[7317])
		); 

/******************* CELL 7318 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7318 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7222]),
			.N(gen[7223]),
			.NE(gen[7224]),

			.O(gen[7317]),
			.E(gen[7319]),

			.SO(gen[7412]),
			.S(gen[7413]),
			.SE(gen[7414]),

			.SELF(gen[7318]),
			.cell_state(gen[7318])
		); 

/******************* CELL 7319 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7319 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7223]),
			.N(gen[7224]),
			.NE(gen[7225]),

			.O(gen[7318]),
			.E(gen[7320]),

			.SO(gen[7413]),
			.S(gen[7414]),
			.SE(gen[7415]),

			.SELF(gen[7319]),
			.cell_state(gen[7319])
		); 

/******************* CELL 7320 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7320 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7224]),
			.N(gen[7225]),
			.NE(gen[7226]),

			.O(gen[7319]),
			.E(gen[7321]),

			.SO(gen[7414]),
			.S(gen[7415]),
			.SE(gen[7416]),

			.SELF(gen[7320]),
			.cell_state(gen[7320])
		); 

/******************* CELL 7321 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7321 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7225]),
			.N(gen[7226]),
			.NE(gen[7227]),

			.O(gen[7320]),
			.E(gen[7322]),

			.SO(gen[7415]),
			.S(gen[7416]),
			.SE(gen[7417]),

			.SELF(gen[7321]),
			.cell_state(gen[7321])
		); 

/******************* CELL 7322 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7322 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7226]),
			.N(gen[7227]),
			.NE(gen[7228]),

			.O(gen[7321]),
			.E(gen[7323]),

			.SO(gen[7416]),
			.S(gen[7417]),
			.SE(gen[7418]),

			.SELF(gen[7322]),
			.cell_state(gen[7322])
		); 

/******************* CELL 7323 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7323 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7227]),
			.N(gen[7228]),
			.NE(gen[7229]),

			.O(gen[7322]),
			.E(gen[7324]),

			.SO(gen[7417]),
			.S(gen[7418]),
			.SE(gen[7419]),

			.SELF(gen[7323]),
			.cell_state(gen[7323])
		); 

/******************* CELL 7324 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7324 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7228]),
			.N(gen[7229]),
			.NE(gen[7230]),

			.O(gen[7323]),
			.E(gen[7325]),

			.SO(gen[7418]),
			.S(gen[7419]),
			.SE(gen[7420]),

			.SELF(gen[7324]),
			.cell_state(gen[7324])
		); 

/******************* CELL 7325 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7325 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7229]),
			.N(gen[7230]),
			.NE(gen[7231]),

			.O(gen[7324]),
			.E(gen[7326]),

			.SO(gen[7419]),
			.S(gen[7420]),
			.SE(gen[7421]),

			.SELF(gen[7325]),
			.cell_state(gen[7325])
		); 

/******************* CELL 7326 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7326 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7230]),
			.N(gen[7231]),
			.NE(gen[7232]),

			.O(gen[7325]),
			.E(gen[7327]),

			.SO(gen[7420]),
			.S(gen[7421]),
			.SE(gen[7422]),

			.SELF(gen[7326]),
			.cell_state(gen[7326])
		); 

/******************* CELL 7327 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7327 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7231]),
			.N(gen[7232]),
			.NE(gen[7233]),

			.O(gen[7326]),
			.E(gen[7328]),

			.SO(gen[7421]),
			.S(gen[7422]),
			.SE(gen[7423]),

			.SELF(gen[7327]),
			.cell_state(gen[7327])
		); 

/******************* CELL 7328 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7328 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7232]),
			.N(gen[7233]),
			.NE(gen[7234]),

			.O(gen[7327]),
			.E(gen[7329]),

			.SO(gen[7422]),
			.S(gen[7423]),
			.SE(gen[7424]),

			.SELF(gen[7328]),
			.cell_state(gen[7328])
		); 

/******************* CELL 7329 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7329 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7233]),
			.N(gen[7234]),
			.NE(gen[7235]),

			.O(gen[7328]),
			.E(gen[7330]),

			.SO(gen[7423]),
			.S(gen[7424]),
			.SE(gen[7425]),

			.SELF(gen[7329]),
			.cell_state(gen[7329])
		); 

/******************* CELL 7330 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7330 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7234]),
			.N(gen[7235]),
			.NE(gen[7236]),

			.O(gen[7329]),
			.E(gen[7331]),

			.SO(gen[7424]),
			.S(gen[7425]),
			.SE(gen[7426]),

			.SELF(gen[7330]),
			.cell_state(gen[7330])
		); 

/******************* CELL 7331 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7331 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7235]),
			.N(gen[7236]),
			.NE(gen[7237]),

			.O(gen[7330]),
			.E(gen[7332]),

			.SO(gen[7425]),
			.S(gen[7426]),
			.SE(gen[7427]),

			.SELF(gen[7331]),
			.cell_state(gen[7331])
		); 

/******************* CELL 7332 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7332 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7236]),
			.N(gen[7237]),
			.NE(gen[7238]),

			.O(gen[7331]),
			.E(gen[7333]),

			.SO(gen[7426]),
			.S(gen[7427]),
			.SE(gen[7428]),

			.SELF(gen[7332]),
			.cell_state(gen[7332])
		); 

/******************* CELL 7333 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7333 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7237]),
			.N(gen[7238]),
			.NE(gen[7239]),

			.O(gen[7332]),
			.E(gen[7334]),

			.SO(gen[7427]),
			.S(gen[7428]),
			.SE(gen[7429]),

			.SELF(gen[7333]),
			.cell_state(gen[7333])
		); 

/******************* CELL 7334 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7334 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7238]),
			.N(gen[7239]),
			.NE(gen[7240]),

			.O(gen[7333]),
			.E(gen[7335]),

			.SO(gen[7428]),
			.S(gen[7429]),
			.SE(gen[7430]),

			.SELF(gen[7334]),
			.cell_state(gen[7334])
		); 

/******************* CELL 7335 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7335 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7239]),
			.N(gen[7240]),
			.NE(gen[7241]),

			.O(gen[7334]),
			.E(gen[7336]),

			.SO(gen[7429]),
			.S(gen[7430]),
			.SE(gen[7431]),

			.SELF(gen[7335]),
			.cell_state(gen[7335])
		); 

/******************* CELL 7336 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7336 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7240]),
			.N(gen[7241]),
			.NE(gen[7242]),

			.O(gen[7335]),
			.E(gen[7337]),

			.SO(gen[7430]),
			.S(gen[7431]),
			.SE(gen[7432]),

			.SELF(gen[7336]),
			.cell_state(gen[7336])
		); 

/******************* CELL 7337 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7337 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7241]),
			.N(gen[7242]),
			.NE(gen[7243]),

			.O(gen[7336]),
			.E(gen[7338]),

			.SO(gen[7431]),
			.S(gen[7432]),
			.SE(gen[7433]),

			.SELF(gen[7337]),
			.cell_state(gen[7337])
		); 

/******************* CELL 7338 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7338 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7242]),
			.N(gen[7243]),
			.NE(gen[7244]),

			.O(gen[7337]),
			.E(gen[7339]),

			.SO(gen[7432]),
			.S(gen[7433]),
			.SE(gen[7434]),

			.SELF(gen[7338]),
			.cell_state(gen[7338])
		); 

/******************* CELL 7339 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7339 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7243]),
			.N(gen[7244]),
			.NE(gen[7245]),

			.O(gen[7338]),
			.E(gen[7340]),

			.SO(gen[7433]),
			.S(gen[7434]),
			.SE(gen[7435]),

			.SELF(gen[7339]),
			.cell_state(gen[7339])
		); 

/******************* CELL 7340 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7340 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7244]),
			.N(gen[7245]),
			.NE(gen[7246]),

			.O(gen[7339]),
			.E(gen[7341]),

			.SO(gen[7434]),
			.S(gen[7435]),
			.SE(gen[7436]),

			.SELF(gen[7340]),
			.cell_state(gen[7340])
		); 

/******************* CELL 7341 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7341 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7245]),
			.N(gen[7246]),
			.NE(gen[7247]),

			.O(gen[7340]),
			.E(gen[7342]),

			.SO(gen[7435]),
			.S(gen[7436]),
			.SE(gen[7437]),

			.SELF(gen[7341]),
			.cell_state(gen[7341])
		); 

/******************* CELL 7342 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7342 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7246]),
			.N(gen[7247]),
			.NE(gen[7248]),

			.O(gen[7341]),
			.E(gen[7343]),

			.SO(gen[7436]),
			.S(gen[7437]),
			.SE(gen[7438]),

			.SELF(gen[7342]),
			.cell_state(gen[7342])
		); 

/******************* CELL 7343 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7343 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7247]),
			.N(gen[7248]),
			.NE(gen[7249]),

			.O(gen[7342]),
			.E(gen[7344]),

			.SO(gen[7437]),
			.S(gen[7438]),
			.SE(gen[7439]),

			.SELF(gen[7343]),
			.cell_state(gen[7343])
		); 

/******************* CELL 7344 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7344 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7248]),
			.N(gen[7249]),
			.NE(gen[7250]),

			.O(gen[7343]),
			.E(gen[7345]),

			.SO(gen[7438]),
			.S(gen[7439]),
			.SE(gen[7440]),

			.SELF(gen[7344]),
			.cell_state(gen[7344])
		); 

/******************* CELL 7345 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7345 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7249]),
			.N(gen[7250]),
			.NE(gen[7251]),

			.O(gen[7344]),
			.E(gen[7346]),

			.SO(gen[7439]),
			.S(gen[7440]),
			.SE(gen[7441]),

			.SELF(gen[7345]),
			.cell_state(gen[7345])
		); 

/******************* CELL 7346 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7346 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7250]),
			.N(gen[7251]),
			.NE(gen[7252]),

			.O(gen[7345]),
			.E(gen[7347]),

			.SO(gen[7440]),
			.S(gen[7441]),
			.SE(gen[7442]),

			.SELF(gen[7346]),
			.cell_state(gen[7346])
		); 

/******************* CELL 7347 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7347 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7251]),
			.N(gen[7252]),
			.NE(gen[7253]),

			.O(gen[7346]),
			.E(gen[7348]),

			.SO(gen[7441]),
			.S(gen[7442]),
			.SE(gen[7443]),

			.SELF(gen[7347]),
			.cell_state(gen[7347])
		); 

/******************* CELL 7348 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7348 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7252]),
			.N(gen[7253]),
			.NE(gen[7254]),

			.O(gen[7347]),
			.E(gen[7349]),

			.SO(gen[7442]),
			.S(gen[7443]),
			.SE(gen[7444]),

			.SELF(gen[7348]),
			.cell_state(gen[7348])
		); 

/******************* CELL 7349 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7349 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7253]),
			.N(gen[7254]),
			.NE(gen[7255]),

			.O(gen[7348]),
			.E(gen[7350]),

			.SO(gen[7443]),
			.S(gen[7444]),
			.SE(gen[7445]),

			.SELF(gen[7349]),
			.cell_state(gen[7349])
		); 

/******************* CELL 7350 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7350 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7254]),
			.N(gen[7255]),
			.NE(gen[7256]),

			.O(gen[7349]),
			.E(gen[7351]),

			.SO(gen[7444]),
			.S(gen[7445]),
			.SE(gen[7446]),

			.SELF(gen[7350]),
			.cell_state(gen[7350])
		); 

/******************* CELL 7351 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7351 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7255]),
			.N(gen[7256]),
			.NE(gen[7257]),

			.O(gen[7350]),
			.E(gen[7352]),

			.SO(gen[7445]),
			.S(gen[7446]),
			.SE(gen[7447]),

			.SELF(gen[7351]),
			.cell_state(gen[7351])
		); 

/******************* CELL 7352 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7352 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7256]),
			.N(gen[7257]),
			.NE(gen[7258]),

			.O(gen[7351]),
			.E(gen[7353]),

			.SO(gen[7446]),
			.S(gen[7447]),
			.SE(gen[7448]),

			.SELF(gen[7352]),
			.cell_state(gen[7352])
		); 

/******************* CELL 7353 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7353 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7257]),
			.N(gen[7258]),
			.NE(gen[7259]),

			.O(gen[7352]),
			.E(gen[7354]),

			.SO(gen[7447]),
			.S(gen[7448]),
			.SE(gen[7449]),

			.SELF(gen[7353]),
			.cell_state(gen[7353])
		); 

/******************* CELL 7354 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7354 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7258]),
			.N(gen[7259]),
			.NE(gen[7260]),

			.O(gen[7353]),
			.E(gen[7355]),

			.SO(gen[7448]),
			.S(gen[7449]),
			.SE(gen[7450]),

			.SELF(gen[7354]),
			.cell_state(gen[7354])
		); 

/******************* CELL 7355 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7355 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7259]),
			.N(gen[7260]),
			.NE(gen[7261]),

			.O(gen[7354]),
			.E(gen[7356]),

			.SO(gen[7449]),
			.S(gen[7450]),
			.SE(gen[7451]),

			.SELF(gen[7355]),
			.cell_state(gen[7355])
		); 

/******************* CELL 7356 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7356 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7260]),
			.N(gen[7261]),
			.NE(gen[7262]),

			.O(gen[7355]),
			.E(gen[7357]),

			.SO(gen[7450]),
			.S(gen[7451]),
			.SE(gen[7452]),

			.SELF(gen[7356]),
			.cell_state(gen[7356])
		); 

/******************* CELL 7357 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7357 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7261]),
			.N(gen[7262]),
			.NE(gen[7263]),

			.O(gen[7356]),
			.E(gen[7358]),

			.SO(gen[7451]),
			.S(gen[7452]),
			.SE(gen[7453]),

			.SELF(gen[7357]),
			.cell_state(gen[7357])
		); 

/******************* CELL 7358 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7358 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7262]),
			.N(gen[7263]),
			.NE(gen[7264]),

			.O(gen[7357]),
			.E(gen[7359]),

			.SO(gen[7452]),
			.S(gen[7453]),
			.SE(gen[7454]),

			.SELF(gen[7358]),
			.cell_state(gen[7358])
		); 

/******************* CELL 7359 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7359 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7263]),
			.N(gen[7264]),
			.NE(gen[7265]),

			.O(gen[7358]),
			.E(gen[7360]),

			.SO(gen[7453]),
			.S(gen[7454]),
			.SE(gen[7455]),

			.SELF(gen[7359]),
			.cell_state(gen[7359])
		); 

/******************* CELL 7360 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7360 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7264]),
			.N(gen[7265]),
			.NE(gen[7266]),

			.O(gen[7359]),
			.E(gen[7361]),

			.SO(gen[7454]),
			.S(gen[7455]),
			.SE(gen[7456]),

			.SELF(gen[7360]),
			.cell_state(gen[7360])
		); 

/******************* CELL 7361 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7361 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7265]),
			.N(gen[7266]),
			.NE(gen[7267]),

			.O(gen[7360]),
			.E(gen[7362]),

			.SO(gen[7455]),
			.S(gen[7456]),
			.SE(gen[7457]),

			.SELF(gen[7361]),
			.cell_state(gen[7361])
		); 

/******************* CELL 7362 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7362 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7266]),
			.N(gen[7267]),
			.NE(gen[7268]),

			.O(gen[7361]),
			.E(gen[7363]),

			.SO(gen[7456]),
			.S(gen[7457]),
			.SE(gen[7458]),

			.SELF(gen[7362]),
			.cell_state(gen[7362])
		); 

/******************* CELL 7363 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7363 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7267]),
			.N(gen[7268]),
			.NE(gen[7269]),

			.O(gen[7362]),
			.E(gen[7364]),

			.SO(gen[7457]),
			.S(gen[7458]),
			.SE(gen[7459]),

			.SELF(gen[7363]),
			.cell_state(gen[7363])
		); 

/******************* CELL 7364 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7364 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7268]),
			.N(gen[7269]),
			.NE(gen[7270]),

			.O(gen[7363]),
			.E(gen[7365]),

			.SO(gen[7458]),
			.S(gen[7459]),
			.SE(gen[7460]),

			.SELF(gen[7364]),
			.cell_state(gen[7364])
		); 

/******************* CELL 7365 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7365 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7269]),
			.N(gen[7270]),
			.NE(gen[7271]),

			.O(gen[7364]),
			.E(gen[7366]),

			.SO(gen[7459]),
			.S(gen[7460]),
			.SE(gen[7461]),

			.SELF(gen[7365]),
			.cell_state(gen[7365])
		); 

/******************* CELL 7366 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7366 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7270]),
			.N(gen[7271]),
			.NE(gen[7272]),

			.O(gen[7365]),
			.E(gen[7367]),

			.SO(gen[7460]),
			.S(gen[7461]),
			.SE(gen[7462]),

			.SELF(gen[7366]),
			.cell_state(gen[7366])
		); 

/******************* CELL 7367 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7367 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7271]),
			.N(gen[7272]),
			.NE(gen[7273]),

			.O(gen[7366]),
			.E(gen[7368]),

			.SO(gen[7461]),
			.S(gen[7462]),
			.SE(gen[7463]),

			.SELF(gen[7367]),
			.cell_state(gen[7367])
		); 

/******************* CELL 7368 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7368 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7272]),
			.N(gen[7273]),
			.NE(gen[7274]),

			.O(gen[7367]),
			.E(gen[7369]),

			.SO(gen[7462]),
			.S(gen[7463]),
			.SE(gen[7464]),

			.SELF(gen[7368]),
			.cell_state(gen[7368])
		); 

/******************* CELL 7369 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7369 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7273]),
			.N(gen[7274]),
			.NE(gen[7275]),

			.O(gen[7368]),
			.E(gen[7370]),

			.SO(gen[7463]),
			.S(gen[7464]),
			.SE(gen[7465]),

			.SELF(gen[7369]),
			.cell_state(gen[7369])
		); 

/******************* CELL 7370 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7370 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7274]),
			.N(gen[7275]),
			.NE(gen[7276]),

			.O(gen[7369]),
			.E(gen[7371]),

			.SO(gen[7464]),
			.S(gen[7465]),
			.SE(gen[7466]),

			.SELF(gen[7370]),
			.cell_state(gen[7370])
		); 

/******************* CELL 7371 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7371 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7275]),
			.N(gen[7276]),
			.NE(gen[7277]),

			.O(gen[7370]),
			.E(gen[7372]),

			.SO(gen[7465]),
			.S(gen[7466]),
			.SE(gen[7467]),

			.SELF(gen[7371]),
			.cell_state(gen[7371])
		); 

/******************* CELL 7372 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7372 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7276]),
			.N(gen[7277]),
			.NE(gen[7278]),

			.O(gen[7371]),
			.E(gen[7373]),

			.SO(gen[7466]),
			.S(gen[7467]),
			.SE(gen[7468]),

			.SELF(gen[7372]),
			.cell_state(gen[7372])
		); 

/******************* CELL 7373 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7373 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7277]),
			.N(gen[7278]),
			.NE(gen[7279]),

			.O(gen[7372]),
			.E(gen[7374]),

			.SO(gen[7467]),
			.S(gen[7468]),
			.SE(gen[7469]),

			.SELF(gen[7373]),
			.cell_state(gen[7373])
		); 

/******************* CELL 7374 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7374 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7278]),
			.N(gen[7279]),
			.NE(gen[7280]),

			.O(gen[7373]),
			.E(gen[7375]),

			.SO(gen[7468]),
			.S(gen[7469]),
			.SE(gen[7470]),

			.SELF(gen[7374]),
			.cell_state(gen[7374])
		); 

/******************* CELL 7375 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7375 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7279]),
			.N(gen[7280]),
			.NE(gen[7281]),

			.O(gen[7374]),
			.E(gen[7376]),

			.SO(gen[7469]),
			.S(gen[7470]),
			.SE(gen[7471]),

			.SELF(gen[7375]),
			.cell_state(gen[7375])
		); 

/******************* CELL 7376 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7376 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7280]),
			.N(gen[7281]),
			.NE(gen[7282]),

			.O(gen[7375]),
			.E(gen[7377]),

			.SO(gen[7470]),
			.S(gen[7471]),
			.SE(gen[7472]),

			.SELF(gen[7376]),
			.cell_state(gen[7376])
		); 

/******************* CELL 7377 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7377 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7281]),
			.N(gen[7282]),
			.NE(gen[7283]),

			.O(gen[7376]),
			.E(gen[7378]),

			.SO(gen[7471]),
			.S(gen[7472]),
			.SE(gen[7473]),

			.SELF(gen[7377]),
			.cell_state(gen[7377])
		); 

/******************* CELL 7378 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7378 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7282]),
			.N(gen[7283]),
			.NE(gen[7284]),

			.O(gen[7377]),
			.E(gen[7379]),

			.SO(gen[7472]),
			.S(gen[7473]),
			.SE(gen[7474]),

			.SELF(gen[7378]),
			.cell_state(gen[7378])
		); 

/******************* CELL 7379 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7379 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7283]),
			.N(gen[7284]),
			.NE(gen[7285]),

			.O(gen[7378]),
			.E(gen[7380]),

			.SO(gen[7473]),
			.S(gen[7474]),
			.SE(gen[7475]),

			.SELF(gen[7379]),
			.cell_state(gen[7379])
		); 

/******************* CELL 7380 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7380 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7284]),
			.N(gen[7285]),
			.NE(gen[7286]),

			.O(gen[7379]),
			.E(gen[7381]),

			.SO(gen[7474]),
			.S(gen[7475]),
			.SE(gen[7476]),

			.SELF(gen[7380]),
			.cell_state(gen[7380])
		); 

/******************* CELL 7381 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7381 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7285]),
			.N(gen[7286]),
			.NE(gen[7287]),

			.O(gen[7380]),
			.E(gen[7382]),

			.SO(gen[7475]),
			.S(gen[7476]),
			.SE(gen[7477]),

			.SELF(gen[7381]),
			.cell_state(gen[7381])
		); 

/******************* CELL 7382 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7382 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7286]),
			.N(gen[7287]),
			.NE(gen[7288]),

			.O(gen[7381]),
			.E(gen[7383]),

			.SO(gen[7476]),
			.S(gen[7477]),
			.SE(gen[7478]),

			.SELF(gen[7382]),
			.cell_state(gen[7382])
		); 

/******************* CELL 7383 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7383 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7287]),
			.N(gen[7288]),
			.NE(gen[7289]),

			.O(gen[7382]),
			.E(gen[7384]),

			.SO(gen[7477]),
			.S(gen[7478]),
			.SE(gen[7479]),

			.SELF(gen[7383]),
			.cell_state(gen[7383])
		); 

/******************* CELL 7384 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7384 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7288]),
			.N(gen[7289]),
			.NE(gen[7290]),

			.O(gen[7383]),
			.E(gen[7385]),

			.SO(gen[7478]),
			.S(gen[7479]),
			.SE(gen[7480]),

			.SELF(gen[7384]),
			.cell_state(gen[7384])
		); 

/******************* CELL 7385 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7385 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7289]),
			.N(gen[7290]),
			.NE(gen[7291]),

			.O(gen[7384]),
			.E(gen[7386]),

			.SO(gen[7479]),
			.S(gen[7480]),
			.SE(gen[7481]),

			.SELF(gen[7385]),
			.cell_state(gen[7385])
		); 

/******************* CELL 7386 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7386 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7290]),
			.N(gen[7291]),
			.NE(gen[7292]),

			.O(gen[7385]),
			.E(gen[7387]),

			.SO(gen[7480]),
			.S(gen[7481]),
			.SE(gen[7482]),

			.SELF(gen[7386]),
			.cell_state(gen[7386])
		); 

/******************* CELL 7387 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7387 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7291]),
			.N(gen[7292]),
			.NE(gen[7293]),

			.O(gen[7386]),
			.E(gen[7388]),

			.SO(gen[7481]),
			.S(gen[7482]),
			.SE(gen[7483]),

			.SELF(gen[7387]),
			.cell_state(gen[7387])
		); 

/******************* CELL 7388 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7388 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7292]),
			.N(gen[7293]),
			.NE(gen[7294]),

			.O(gen[7387]),
			.E(gen[7389]),

			.SO(gen[7482]),
			.S(gen[7483]),
			.SE(gen[7484]),

			.SELF(gen[7388]),
			.cell_state(gen[7388])
		); 

/******************* CELL 7389 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7389 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7293]),
			.N(gen[7294]),
			.NE(gen[7295]),

			.O(gen[7388]),
			.E(gen[7390]),

			.SO(gen[7483]),
			.S(gen[7484]),
			.SE(gen[7485]),

			.SELF(gen[7389]),
			.cell_state(gen[7389])
		); 

/******************* CELL 7390 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7390 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7294]),
			.N(gen[7295]),
			.NE(gen[7296]),

			.O(gen[7389]),
			.E(gen[7391]),

			.SO(gen[7484]),
			.S(gen[7485]),
			.SE(gen[7486]),

			.SELF(gen[7390]),
			.cell_state(gen[7390])
		); 

/******************* CELL 7391 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7391 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7295]),
			.N(gen[7296]),
			.NE(gen[7297]),

			.O(gen[7390]),
			.E(gen[7392]),

			.SO(gen[7485]),
			.S(gen[7486]),
			.SE(gen[7487]),

			.SELF(gen[7391]),
			.cell_state(gen[7391])
		); 

/******************* CELL 7392 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7392 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7296]),
			.N(gen[7297]),
			.NE(gen[7298]),

			.O(gen[7391]),
			.E(gen[7393]),

			.SO(gen[7486]),
			.S(gen[7487]),
			.SE(gen[7488]),

			.SELF(gen[7392]),
			.cell_state(gen[7392])
		); 

/******************* CELL 7393 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7393 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7297]),
			.N(gen[7298]),
			.NE(gen[7299]),

			.O(gen[7392]),
			.E(gen[7394]),

			.SO(gen[7487]),
			.S(gen[7488]),
			.SE(gen[7489]),

			.SELF(gen[7393]),
			.cell_state(gen[7393])
		); 

/******************* CELL 7394 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7394 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7298]),
			.N(gen[7299]),
			.NE(gen[7300]),

			.O(gen[7393]),
			.E(gen[7395]),

			.SO(gen[7488]),
			.S(gen[7489]),
			.SE(gen[7490]),

			.SELF(gen[7394]),
			.cell_state(gen[7394])
		); 

/******************* CELL 7395 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7395 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7299]),
			.N(gen[7300]),
			.NE(gen[7301]),

			.O(gen[7394]),
			.E(gen[7396]),

			.SO(gen[7489]),
			.S(gen[7490]),
			.SE(gen[7491]),

			.SELF(gen[7395]),
			.cell_state(gen[7395])
		); 

/******************* CELL 7396 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7396 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7300]),
			.N(gen[7301]),
			.NE(gen[7302]),

			.O(gen[7395]),
			.E(gen[7397]),

			.SO(gen[7490]),
			.S(gen[7491]),
			.SE(gen[7492]),

			.SELF(gen[7396]),
			.cell_state(gen[7396])
		); 

/******************* CELL 7397 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7397 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7301]),
			.N(gen[7302]),
			.NE(gen[7303]),

			.O(gen[7396]),
			.E(gen[7398]),

			.SO(gen[7491]),
			.S(gen[7492]),
			.SE(gen[7493]),

			.SELF(gen[7397]),
			.cell_state(gen[7397])
		); 

/******************* CELL 7398 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7398 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7302]),
			.N(gen[7303]),
			.NE(gen[7304]),

			.O(gen[7397]),
			.E(gen[7399]),

			.SO(gen[7492]),
			.S(gen[7493]),
			.SE(gen[7494]),

			.SELF(gen[7398]),
			.cell_state(gen[7398])
		); 

/******************* CELL 7399 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7399 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7303]),
			.N(gen[7304]),
			.NE(gen[7305]),

			.O(gen[7398]),
			.E(gen[7400]),

			.SO(gen[7493]),
			.S(gen[7494]),
			.SE(gen[7495]),

			.SELF(gen[7399]),
			.cell_state(gen[7399])
		); 

/******************* CELL 7400 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7400 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7304]),
			.N(gen[7305]),
			.NE(gen[7306]),

			.O(gen[7399]),
			.E(gen[7401]),

			.SO(gen[7494]),
			.S(gen[7495]),
			.SE(gen[7496]),

			.SELF(gen[7400]),
			.cell_state(gen[7400])
		); 

/******************* CELL 7401 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7401 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7305]),
			.N(gen[7306]),
			.NE(gen[7307]),

			.O(gen[7400]),
			.E(gen[7402]),

			.SO(gen[7495]),
			.S(gen[7496]),
			.SE(gen[7497]),

			.SELF(gen[7401]),
			.cell_state(gen[7401])
		); 

/******************* CELL 7402 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7402 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7306]),
			.N(gen[7307]),
			.NE(gen[7308]),

			.O(gen[7401]),
			.E(gen[7403]),

			.SO(gen[7496]),
			.S(gen[7497]),
			.SE(gen[7498]),

			.SELF(gen[7402]),
			.cell_state(gen[7402])
		); 

/******************* CELL 7403 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7403 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7307]),
			.N(gen[7308]),
			.NE(gen[7309]),

			.O(gen[7402]),
			.E(gen[7404]),

			.SO(gen[7497]),
			.S(gen[7498]),
			.SE(gen[7499]),

			.SELF(gen[7403]),
			.cell_state(gen[7403])
		); 

/******************* CELL 7404 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7404 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7308]),
			.N(gen[7309]),
			.NE(gen[7310]),

			.O(gen[7403]),
			.E(gen[7405]),

			.SO(gen[7498]),
			.S(gen[7499]),
			.SE(gen[7500]),

			.SELF(gen[7404]),
			.cell_state(gen[7404])
		); 

/******************* CELL 7405 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7405 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7309]),
			.N(gen[7310]),
			.NE(gen[7311]),

			.O(gen[7404]),
			.E(gen[7406]),

			.SO(gen[7499]),
			.S(gen[7500]),
			.SE(gen[7501]),

			.SELF(gen[7405]),
			.cell_state(gen[7405])
		); 

/******************* CELL 7406 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7406 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7310]),
			.N(gen[7311]),
			.NE(gen[7312]),

			.O(gen[7405]),
			.E(gen[7407]),

			.SO(gen[7500]),
			.S(gen[7501]),
			.SE(gen[7502]),

			.SELF(gen[7406]),
			.cell_state(gen[7406])
		); 

/******************* CELL 7407 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7407 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7311]),
			.N(gen[7312]),
			.NE(gen[7313]),

			.O(gen[7406]),
			.E(gen[7408]),

			.SO(gen[7501]),
			.S(gen[7502]),
			.SE(gen[7503]),

			.SELF(gen[7407]),
			.cell_state(gen[7407])
		); 

/******************* CELL 7408 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7408 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7312]),
			.N(gen[7313]),
			.NE(gen[7314]),

			.O(gen[7407]),
			.E(gen[7409]),

			.SO(gen[7502]),
			.S(gen[7503]),
			.SE(gen[7504]),

			.SELF(gen[7408]),
			.cell_state(gen[7408])
		); 

/******************* CELL 7409 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7409 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7313]),
			.N(gen[7314]),
			.NE(gen[7313]),

			.O(gen[7408]),
			.E(gen[7408]),

			.SO(gen[7503]),
			.S(gen[7504]),
			.SE(gen[7503]),

			.SELF(gen[7409]),
			.cell_state(gen[7409])
		); 

/******************* CELL 7410 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7410 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7316]),
			.N(gen[7315]),
			.NE(gen[7316]),

			.O(gen[7411]),
			.E(gen[7411]),

			.SO(gen[7506]),
			.S(gen[7505]),
			.SE(gen[7506]),

			.SELF(gen[7410]),
			.cell_state(gen[7410])
		); 

/******************* CELL 7411 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7411 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7315]),
			.N(gen[7316]),
			.NE(gen[7317]),

			.O(gen[7410]),
			.E(gen[7412]),

			.SO(gen[7505]),
			.S(gen[7506]),
			.SE(gen[7507]),

			.SELF(gen[7411]),
			.cell_state(gen[7411])
		); 

/******************* CELL 7412 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7412 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7316]),
			.N(gen[7317]),
			.NE(gen[7318]),

			.O(gen[7411]),
			.E(gen[7413]),

			.SO(gen[7506]),
			.S(gen[7507]),
			.SE(gen[7508]),

			.SELF(gen[7412]),
			.cell_state(gen[7412])
		); 

/******************* CELL 7413 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7413 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7317]),
			.N(gen[7318]),
			.NE(gen[7319]),

			.O(gen[7412]),
			.E(gen[7414]),

			.SO(gen[7507]),
			.S(gen[7508]),
			.SE(gen[7509]),

			.SELF(gen[7413]),
			.cell_state(gen[7413])
		); 

/******************* CELL 7414 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7414 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7318]),
			.N(gen[7319]),
			.NE(gen[7320]),

			.O(gen[7413]),
			.E(gen[7415]),

			.SO(gen[7508]),
			.S(gen[7509]),
			.SE(gen[7510]),

			.SELF(gen[7414]),
			.cell_state(gen[7414])
		); 

/******************* CELL 7415 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7415 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7319]),
			.N(gen[7320]),
			.NE(gen[7321]),

			.O(gen[7414]),
			.E(gen[7416]),

			.SO(gen[7509]),
			.S(gen[7510]),
			.SE(gen[7511]),

			.SELF(gen[7415]),
			.cell_state(gen[7415])
		); 

/******************* CELL 7416 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7416 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7320]),
			.N(gen[7321]),
			.NE(gen[7322]),

			.O(gen[7415]),
			.E(gen[7417]),

			.SO(gen[7510]),
			.S(gen[7511]),
			.SE(gen[7512]),

			.SELF(gen[7416]),
			.cell_state(gen[7416])
		); 

/******************* CELL 7417 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7417 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7321]),
			.N(gen[7322]),
			.NE(gen[7323]),

			.O(gen[7416]),
			.E(gen[7418]),

			.SO(gen[7511]),
			.S(gen[7512]),
			.SE(gen[7513]),

			.SELF(gen[7417]),
			.cell_state(gen[7417])
		); 

/******************* CELL 7418 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7418 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7322]),
			.N(gen[7323]),
			.NE(gen[7324]),

			.O(gen[7417]),
			.E(gen[7419]),

			.SO(gen[7512]),
			.S(gen[7513]),
			.SE(gen[7514]),

			.SELF(gen[7418]),
			.cell_state(gen[7418])
		); 

/******************* CELL 7419 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7419 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7323]),
			.N(gen[7324]),
			.NE(gen[7325]),

			.O(gen[7418]),
			.E(gen[7420]),

			.SO(gen[7513]),
			.S(gen[7514]),
			.SE(gen[7515]),

			.SELF(gen[7419]),
			.cell_state(gen[7419])
		); 

/******************* CELL 7420 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7420 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7324]),
			.N(gen[7325]),
			.NE(gen[7326]),

			.O(gen[7419]),
			.E(gen[7421]),

			.SO(gen[7514]),
			.S(gen[7515]),
			.SE(gen[7516]),

			.SELF(gen[7420]),
			.cell_state(gen[7420])
		); 

/******************* CELL 7421 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7421 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7325]),
			.N(gen[7326]),
			.NE(gen[7327]),

			.O(gen[7420]),
			.E(gen[7422]),

			.SO(gen[7515]),
			.S(gen[7516]),
			.SE(gen[7517]),

			.SELF(gen[7421]),
			.cell_state(gen[7421])
		); 

/******************* CELL 7422 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7422 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7326]),
			.N(gen[7327]),
			.NE(gen[7328]),

			.O(gen[7421]),
			.E(gen[7423]),

			.SO(gen[7516]),
			.S(gen[7517]),
			.SE(gen[7518]),

			.SELF(gen[7422]),
			.cell_state(gen[7422])
		); 

/******************* CELL 7423 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7423 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7327]),
			.N(gen[7328]),
			.NE(gen[7329]),

			.O(gen[7422]),
			.E(gen[7424]),

			.SO(gen[7517]),
			.S(gen[7518]),
			.SE(gen[7519]),

			.SELF(gen[7423]),
			.cell_state(gen[7423])
		); 

/******************* CELL 7424 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7424 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7328]),
			.N(gen[7329]),
			.NE(gen[7330]),

			.O(gen[7423]),
			.E(gen[7425]),

			.SO(gen[7518]),
			.S(gen[7519]),
			.SE(gen[7520]),

			.SELF(gen[7424]),
			.cell_state(gen[7424])
		); 

/******************* CELL 7425 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7425 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7329]),
			.N(gen[7330]),
			.NE(gen[7331]),

			.O(gen[7424]),
			.E(gen[7426]),

			.SO(gen[7519]),
			.S(gen[7520]),
			.SE(gen[7521]),

			.SELF(gen[7425]),
			.cell_state(gen[7425])
		); 

/******************* CELL 7426 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7426 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7330]),
			.N(gen[7331]),
			.NE(gen[7332]),

			.O(gen[7425]),
			.E(gen[7427]),

			.SO(gen[7520]),
			.S(gen[7521]),
			.SE(gen[7522]),

			.SELF(gen[7426]),
			.cell_state(gen[7426])
		); 

/******************* CELL 7427 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7427 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7331]),
			.N(gen[7332]),
			.NE(gen[7333]),

			.O(gen[7426]),
			.E(gen[7428]),

			.SO(gen[7521]),
			.S(gen[7522]),
			.SE(gen[7523]),

			.SELF(gen[7427]),
			.cell_state(gen[7427])
		); 

/******************* CELL 7428 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7428 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7332]),
			.N(gen[7333]),
			.NE(gen[7334]),

			.O(gen[7427]),
			.E(gen[7429]),

			.SO(gen[7522]),
			.S(gen[7523]),
			.SE(gen[7524]),

			.SELF(gen[7428]),
			.cell_state(gen[7428])
		); 

/******************* CELL 7429 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7429 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7333]),
			.N(gen[7334]),
			.NE(gen[7335]),

			.O(gen[7428]),
			.E(gen[7430]),

			.SO(gen[7523]),
			.S(gen[7524]),
			.SE(gen[7525]),

			.SELF(gen[7429]),
			.cell_state(gen[7429])
		); 

/******************* CELL 7430 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7430 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7334]),
			.N(gen[7335]),
			.NE(gen[7336]),

			.O(gen[7429]),
			.E(gen[7431]),

			.SO(gen[7524]),
			.S(gen[7525]),
			.SE(gen[7526]),

			.SELF(gen[7430]),
			.cell_state(gen[7430])
		); 

/******************* CELL 7431 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7431 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7335]),
			.N(gen[7336]),
			.NE(gen[7337]),

			.O(gen[7430]),
			.E(gen[7432]),

			.SO(gen[7525]),
			.S(gen[7526]),
			.SE(gen[7527]),

			.SELF(gen[7431]),
			.cell_state(gen[7431])
		); 

/******************* CELL 7432 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7432 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7336]),
			.N(gen[7337]),
			.NE(gen[7338]),

			.O(gen[7431]),
			.E(gen[7433]),

			.SO(gen[7526]),
			.S(gen[7527]),
			.SE(gen[7528]),

			.SELF(gen[7432]),
			.cell_state(gen[7432])
		); 

/******************* CELL 7433 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7433 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7337]),
			.N(gen[7338]),
			.NE(gen[7339]),

			.O(gen[7432]),
			.E(gen[7434]),

			.SO(gen[7527]),
			.S(gen[7528]),
			.SE(gen[7529]),

			.SELF(gen[7433]),
			.cell_state(gen[7433])
		); 

/******************* CELL 7434 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7434 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7338]),
			.N(gen[7339]),
			.NE(gen[7340]),

			.O(gen[7433]),
			.E(gen[7435]),

			.SO(gen[7528]),
			.S(gen[7529]),
			.SE(gen[7530]),

			.SELF(gen[7434]),
			.cell_state(gen[7434])
		); 

/******************* CELL 7435 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7435 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7339]),
			.N(gen[7340]),
			.NE(gen[7341]),

			.O(gen[7434]),
			.E(gen[7436]),

			.SO(gen[7529]),
			.S(gen[7530]),
			.SE(gen[7531]),

			.SELF(gen[7435]),
			.cell_state(gen[7435])
		); 

/******************* CELL 7436 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7436 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7340]),
			.N(gen[7341]),
			.NE(gen[7342]),

			.O(gen[7435]),
			.E(gen[7437]),

			.SO(gen[7530]),
			.S(gen[7531]),
			.SE(gen[7532]),

			.SELF(gen[7436]),
			.cell_state(gen[7436])
		); 

/******************* CELL 7437 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7437 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7341]),
			.N(gen[7342]),
			.NE(gen[7343]),

			.O(gen[7436]),
			.E(gen[7438]),

			.SO(gen[7531]),
			.S(gen[7532]),
			.SE(gen[7533]),

			.SELF(gen[7437]),
			.cell_state(gen[7437])
		); 

/******************* CELL 7438 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7438 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7342]),
			.N(gen[7343]),
			.NE(gen[7344]),

			.O(gen[7437]),
			.E(gen[7439]),

			.SO(gen[7532]),
			.S(gen[7533]),
			.SE(gen[7534]),

			.SELF(gen[7438]),
			.cell_state(gen[7438])
		); 

/******************* CELL 7439 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7439 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7343]),
			.N(gen[7344]),
			.NE(gen[7345]),

			.O(gen[7438]),
			.E(gen[7440]),

			.SO(gen[7533]),
			.S(gen[7534]),
			.SE(gen[7535]),

			.SELF(gen[7439]),
			.cell_state(gen[7439])
		); 

/******************* CELL 7440 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7440 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7344]),
			.N(gen[7345]),
			.NE(gen[7346]),

			.O(gen[7439]),
			.E(gen[7441]),

			.SO(gen[7534]),
			.S(gen[7535]),
			.SE(gen[7536]),

			.SELF(gen[7440]),
			.cell_state(gen[7440])
		); 

/******************* CELL 7441 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7441 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7345]),
			.N(gen[7346]),
			.NE(gen[7347]),

			.O(gen[7440]),
			.E(gen[7442]),

			.SO(gen[7535]),
			.S(gen[7536]),
			.SE(gen[7537]),

			.SELF(gen[7441]),
			.cell_state(gen[7441])
		); 

/******************* CELL 7442 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7442 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7346]),
			.N(gen[7347]),
			.NE(gen[7348]),

			.O(gen[7441]),
			.E(gen[7443]),

			.SO(gen[7536]),
			.S(gen[7537]),
			.SE(gen[7538]),

			.SELF(gen[7442]),
			.cell_state(gen[7442])
		); 

/******************* CELL 7443 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7443 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7347]),
			.N(gen[7348]),
			.NE(gen[7349]),

			.O(gen[7442]),
			.E(gen[7444]),

			.SO(gen[7537]),
			.S(gen[7538]),
			.SE(gen[7539]),

			.SELF(gen[7443]),
			.cell_state(gen[7443])
		); 

/******************* CELL 7444 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7444 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7348]),
			.N(gen[7349]),
			.NE(gen[7350]),

			.O(gen[7443]),
			.E(gen[7445]),

			.SO(gen[7538]),
			.S(gen[7539]),
			.SE(gen[7540]),

			.SELF(gen[7444]),
			.cell_state(gen[7444])
		); 

/******************* CELL 7445 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7445 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7349]),
			.N(gen[7350]),
			.NE(gen[7351]),

			.O(gen[7444]),
			.E(gen[7446]),

			.SO(gen[7539]),
			.S(gen[7540]),
			.SE(gen[7541]),

			.SELF(gen[7445]),
			.cell_state(gen[7445])
		); 

/******************* CELL 7446 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7446 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7350]),
			.N(gen[7351]),
			.NE(gen[7352]),

			.O(gen[7445]),
			.E(gen[7447]),

			.SO(gen[7540]),
			.S(gen[7541]),
			.SE(gen[7542]),

			.SELF(gen[7446]),
			.cell_state(gen[7446])
		); 

/******************* CELL 7447 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7447 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7351]),
			.N(gen[7352]),
			.NE(gen[7353]),

			.O(gen[7446]),
			.E(gen[7448]),

			.SO(gen[7541]),
			.S(gen[7542]),
			.SE(gen[7543]),

			.SELF(gen[7447]),
			.cell_state(gen[7447])
		); 

/******************* CELL 7448 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7448 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7352]),
			.N(gen[7353]),
			.NE(gen[7354]),

			.O(gen[7447]),
			.E(gen[7449]),

			.SO(gen[7542]),
			.S(gen[7543]),
			.SE(gen[7544]),

			.SELF(gen[7448]),
			.cell_state(gen[7448])
		); 

/******************* CELL 7449 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7449 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7353]),
			.N(gen[7354]),
			.NE(gen[7355]),

			.O(gen[7448]),
			.E(gen[7450]),

			.SO(gen[7543]),
			.S(gen[7544]),
			.SE(gen[7545]),

			.SELF(gen[7449]),
			.cell_state(gen[7449])
		); 

/******************* CELL 7450 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7450 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7354]),
			.N(gen[7355]),
			.NE(gen[7356]),

			.O(gen[7449]),
			.E(gen[7451]),

			.SO(gen[7544]),
			.S(gen[7545]),
			.SE(gen[7546]),

			.SELF(gen[7450]),
			.cell_state(gen[7450])
		); 

/******************* CELL 7451 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7451 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7355]),
			.N(gen[7356]),
			.NE(gen[7357]),

			.O(gen[7450]),
			.E(gen[7452]),

			.SO(gen[7545]),
			.S(gen[7546]),
			.SE(gen[7547]),

			.SELF(gen[7451]),
			.cell_state(gen[7451])
		); 

/******************* CELL 7452 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7452 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7356]),
			.N(gen[7357]),
			.NE(gen[7358]),

			.O(gen[7451]),
			.E(gen[7453]),

			.SO(gen[7546]),
			.S(gen[7547]),
			.SE(gen[7548]),

			.SELF(gen[7452]),
			.cell_state(gen[7452])
		); 

/******************* CELL 7453 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7453 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7357]),
			.N(gen[7358]),
			.NE(gen[7359]),

			.O(gen[7452]),
			.E(gen[7454]),

			.SO(gen[7547]),
			.S(gen[7548]),
			.SE(gen[7549]),

			.SELF(gen[7453]),
			.cell_state(gen[7453])
		); 

/******************* CELL 7454 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7454 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7358]),
			.N(gen[7359]),
			.NE(gen[7360]),

			.O(gen[7453]),
			.E(gen[7455]),

			.SO(gen[7548]),
			.S(gen[7549]),
			.SE(gen[7550]),

			.SELF(gen[7454]),
			.cell_state(gen[7454])
		); 

/******************* CELL 7455 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7455 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7359]),
			.N(gen[7360]),
			.NE(gen[7361]),

			.O(gen[7454]),
			.E(gen[7456]),

			.SO(gen[7549]),
			.S(gen[7550]),
			.SE(gen[7551]),

			.SELF(gen[7455]),
			.cell_state(gen[7455])
		); 

/******************* CELL 7456 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7456 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7360]),
			.N(gen[7361]),
			.NE(gen[7362]),

			.O(gen[7455]),
			.E(gen[7457]),

			.SO(gen[7550]),
			.S(gen[7551]),
			.SE(gen[7552]),

			.SELF(gen[7456]),
			.cell_state(gen[7456])
		); 

/******************* CELL 7457 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7457 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7361]),
			.N(gen[7362]),
			.NE(gen[7363]),

			.O(gen[7456]),
			.E(gen[7458]),

			.SO(gen[7551]),
			.S(gen[7552]),
			.SE(gen[7553]),

			.SELF(gen[7457]),
			.cell_state(gen[7457])
		); 

/******************* CELL 7458 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7458 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7362]),
			.N(gen[7363]),
			.NE(gen[7364]),

			.O(gen[7457]),
			.E(gen[7459]),

			.SO(gen[7552]),
			.S(gen[7553]),
			.SE(gen[7554]),

			.SELF(gen[7458]),
			.cell_state(gen[7458])
		); 

/******************* CELL 7459 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7459 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7363]),
			.N(gen[7364]),
			.NE(gen[7365]),

			.O(gen[7458]),
			.E(gen[7460]),

			.SO(gen[7553]),
			.S(gen[7554]),
			.SE(gen[7555]),

			.SELF(gen[7459]),
			.cell_state(gen[7459])
		); 

/******************* CELL 7460 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7460 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7364]),
			.N(gen[7365]),
			.NE(gen[7366]),

			.O(gen[7459]),
			.E(gen[7461]),

			.SO(gen[7554]),
			.S(gen[7555]),
			.SE(gen[7556]),

			.SELF(gen[7460]),
			.cell_state(gen[7460])
		); 

/******************* CELL 7461 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7461 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7365]),
			.N(gen[7366]),
			.NE(gen[7367]),

			.O(gen[7460]),
			.E(gen[7462]),

			.SO(gen[7555]),
			.S(gen[7556]),
			.SE(gen[7557]),

			.SELF(gen[7461]),
			.cell_state(gen[7461])
		); 

/******************* CELL 7462 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7462 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7366]),
			.N(gen[7367]),
			.NE(gen[7368]),

			.O(gen[7461]),
			.E(gen[7463]),

			.SO(gen[7556]),
			.S(gen[7557]),
			.SE(gen[7558]),

			.SELF(gen[7462]),
			.cell_state(gen[7462])
		); 

/******************* CELL 7463 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7463 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7367]),
			.N(gen[7368]),
			.NE(gen[7369]),

			.O(gen[7462]),
			.E(gen[7464]),

			.SO(gen[7557]),
			.S(gen[7558]),
			.SE(gen[7559]),

			.SELF(gen[7463]),
			.cell_state(gen[7463])
		); 

/******************* CELL 7464 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7464 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7368]),
			.N(gen[7369]),
			.NE(gen[7370]),

			.O(gen[7463]),
			.E(gen[7465]),

			.SO(gen[7558]),
			.S(gen[7559]),
			.SE(gen[7560]),

			.SELF(gen[7464]),
			.cell_state(gen[7464])
		); 

/******************* CELL 7465 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7465 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7369]),
			.N(gen[7370]),
			.NE(gen[7371]),

			.O(gen[7464]),
			.E(gen[7466]),

			.SO(gen[7559]),
			.S(gen[7560]),
			.SE(gen[7561]),

			.SELF(gen[7465]),
			.cell_state(gen[7465])
		); 

/******************* CELL 7466 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7466 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7370]),
			.N(gen[7371]),
			.NE(gen[7372]),

			.O(gen[7465]),
			.E(gen[7467]),

			.SO(gen[7560]),
			.S(gen[7561]),
			.SE(gen[7562]),

			.SELF(gen[7466]),
			.cell_state(gen[7466])
		); 

/******************* CELL 7467 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7467 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7371]),
			.N(gen[7372]),
			.NE(gen[7373]),

			.O(gen[7466]),
			.E(gen[7468]),

			.SO(gen[7561]),
			.S(gen[7562]),
			.SE(gen[7563]),

			.SELF(gen[7467]),
			.cell_state(gen[7467])
		); 

/******************* CELL 7468 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7468 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7372]),
			.N(gen[7373]),
			.NE(gen[7374]),

			.O(gen[7467]),
			.E(gen[7469]),

			.SO(gen[7562]),
			.S(gen[7563]),
			.SE(gen[7564]),

			.SELF(gen[7468]),
			.cell_state(gen[7468])
		); 

/******************* CELL 7469 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7469 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7373]),
			.N(gen[7374]),
			.NE(gen[7375]),

			.O(gen[7468]),
			.E(gen[7470]),

			.SO(gen[7563]),
			.S(gen[7564]),
			.SE(gen[7565]),

			.SELF(gen[7469]),
			.cell_state(gen[7469])
		); 

/******************* CELL 7470 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7470 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7374]),
			.N(gen[7375]),
			.NE(gen[7376]),

			.O(gen[7469]),
			.E(gen[7471]),

			.SO(gen[7564]),
			.S(gen[7565]),
			.SE(gen[7566]),

			.SELF(gen[7470]),
			.cell_state(gen[7470])
		); 

/******************* CELL 7471 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7471 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7375]),
			.N(gen[7376]),
			.NE(gen[7377]),

			.O(gen[7470]),
			.E(gen[7472]),

			.SO(gen[7565]),
			.S(gen[7566]),
			.SE(gen[7567]),

			.SELF(gen[7471]),
			.cell_state(gen[7471])
		); 

/******************* CELL 7472 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7472 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7376]),
			.N(gen[7377]),
			.NE(gen[7378]),

			.O(gen[7471]),
			.E(gen[7473]),

			.SO(gen[7566]),
			.S(gen[7567]),
			.SE(gen[7568]),

			.SELF(gen[7472]),
			.cell_state(gen[7472])
		); 

/******************* CELL 7473 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7473 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7377]),
			.N(gen[7378]),
			.NE(gen[7379]),

			.O(gen[7472]),
			.E(gen[7474]),

			.SO(gen[7567]),
			.S(gen[7568]),
			.SE(gen[7569]),

			.SELF(gen[7473]),
			.cell_state(gen[7473])
		); 

/******************* CELL 7474 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7474 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7378]),
			.N(gen[7379]),
			.NE(gen[7380]),

			.O(gen[7473]),
			.E(gen[7475]),

			.SO(gen[7568]),
			.S(gen[7569]),
			.SE(gen[7570]),

			.SELF(gen[7474]),
			.cell_state(gen[7474])
		); 

/******************* CELL 7475 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7475 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7379]),
			.N(gen[7380]),
			.NE(gen[7381]),

			.O(gen[7474]),
			.E(gen[7476]),

			.SO(gen[7569]),
			.S(gen[7570]),
			.SE(gen[7571]),

			.SELF(gen[7475]),
			.cell_state(gen[7475])
		); 

/******************* CELL 7476 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7476 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7380]),
			.N(gen[7381]),
			.NE(gen[7382]),

			.O(gen[7475]),
			.E(gen[7477]),

			.SO(gen[7570]),
			.S(gen[7571]),
			.SE(gen[7572]),

			.SELF(gen[7476]),
			.cell_state(gen[7476])
		); 

/******************* CELL 7477 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7477 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7381]),
			.N(gen[7382]),
			.NE(gen[7383]),

			.O(gen[7476]),
			.E(gen[7478]),

			.SO(gen[7571]),
			.S(gen[7572]),
			.SE(gen[7573]),

			.SELF(gen[7477]),
			.cell_state(gen[7477])
		); 

/******************* CELL 7478 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7478 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7382]),
			.N(gen[7383]),
			.NE(gen[7384]),

			.O(gen[7477]),
			.E(gen[7479]),

			.SO(gen[7572]),
			.S(gen[7573]),
			.SE(gen[7574]),

			.SELF(gen[7478]),
			.cell_state(gen[7478])
		); 

/******************* CELL 7479 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7479 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7383]),
			.N(gen[7384]),
			.NE(gen[7385]),

			.O(gen[7478]),
			.E(gen[7480]),

			.SO(gen[7573]),
			.S(gen[7574]),
			.SE(gen[7575]),

			.SELF(gen[7479]),
			.cell_state(gen[7479])
		); 

/******************* CELL 7480 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7480 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7384]),
			.N(gen[7385]),
			.NE(gen[7386]),

			.O(gen[7479]),
			.E(gen[7481]),

			.SO(gen[7574]),
			.S(gen[7575]),
			.SE(gen[7576]),

			.SELF(gen[7480]),
			.cell_state(gen[7480])
		); 

/******************* CELL 7481 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7481 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7385]),
			.N(gen[7386]),
			.NE(gen[7387]),

			.O(gen[7480]),
			.E(gen[7482]),

			.SO(gen[7575]),
			.S(gen[7576]),
			.SE(gen[7577]),

			.SELF(gen[7481]),
			.cell_state(gen[7481])
		); 

/******************* CELL 7482 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7482 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7386]),
			.N(gen[7387]),
			.NE(gen[7388]),

			.O(gen[7481]),
			.E(gen[7483]),

			.SO(gen[7576]),
			.S(gen[7577]),
			.SE(gen[7578]),

			.SELF(gen[7482]),
			.cell_state(gen[7482])
		); 

/******************* CELL 7483 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7483 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7387]),
			.N(gen[7388]),
			.NE(gen[7389]),

			.O(gen[7482]),
			.E(gen[7484]),

			.SO(gen[7577]),
			.S(gen[7578]),
			.SE(gen[7579]),

			.SELF(gen[7483]),
			.cell_state(gen[7483])
		); 

/******************* CELL 7484 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7484 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7388]),
			.N(gen[7389]),
			.NE(gen[7390]),

			.O(gen[7483]),
			.E(gen[7485]),

			.SO(gen[7578]),
			.S(gen[7579]),
			.SE(gen[7580]),

			.SELF(gen[7484]),
			.cell_state(gen[7484])
		); 

/******************* CELL 7485 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7485 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7389]),
			.N(gen[7390]),
			.NE(gen[7391]),

			.O(gen[7484]),
			.E(gen[7486]),

			.SO(gen[7579]),
			.S(gen[7580]),
			.SE(gen[7581]),

			.SELF(gen[7485]),
			.cell_state(gen[7485])
		); 

/******************* CELL 7486 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7486 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7390]),
			.N(gen[7391]),
			.NE(gen[7392]),

			.O(gen[7485]),
			.E(gen[7487]),

			.SO(gen[7580]),
			.S(gen[7581]),
			.SE(gen[7582]),

			.SELF(gen[7486]),
			.cell_state(gen[7486])
		); 

/******************* CELL 7487 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7487 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7391]),
			.N(gen[7392]),
			.NE(gen[7393]),

			.O(gen[7486]),
			.E(gen[7488]),

			.SO(gen[7581]),
			.S(gen[7582]),
			.SE(gen[7583]),

			.SELF(gen[7487]),
			.cell_state(gen[7487])
		); 

/******************* CELL 7488 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7488 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7392]),
			.N(gen[7393]),
			.NE(gen[7394]),

			.O(gen[7487]),
			.E(gen[7489]),

			.SO(gen[7582]),
			.S(gen[7583]),
			.SE(gen[7584]),

			.SELF(gen[7488]),
			.cell_state(gen[7488])
		); 

/******************* CELL 7489 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7489 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7393]),
			.N(gen[7394]),
			.NE(gen[7395]),

			.O(gen[7488]),
			.E(gen[7490]),

			.SO(gen[7583]),
			.S(gen[7584]),
			.SE(gen[7585]),

			.SELF(gen[7489]),
			.cell_state(gen[7489])
		); 

/******************* CELL 7490 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7490 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7394]),
			.N(gen[7395]),
			.NE(gen[7396]),

			.O(gen[7489]),
			.E(gen[7491]),

			.SO(gen[7584]),
			.S(gen[7585]),
			.SE(gen[7586]),

			.SELF(gen[7490]),
			.cell_state(gen[7490])
		); 

/******************* CELL 7491 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7491 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7395]),
			.N(gen[7396]),
			.NE(gen[7397]),

			.O(gen[7490]),
			.E(gen[7492]),

			.SO(gen[7585]),
			.S(gen[7586]),
			.SE(gen[7587]),

			.SELF(gen[7491]),
			.cell_state(gen[7491])
		); 

/******************* CELL 7492 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7492 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7396]),
			.N(gen[7397]),
			.NE(gen[7398]),

			.O(gen[7491]),
			.E(gen[7493]),

			.SO(gen[7586]),
			.S(gen[7587]),
			.SE(gen[7588]),

			.SELF(gen[7492]),
			.cell_state(gen[7492])
		); 

/******************* CELL 7493 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7493 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7397]),
			.N(gen[7398]),
			.NE(gen[7399]),

			.O(gen[7492]),
			.E(gen[7494]),

			.SO(gen[7587]),
			.S(gen[7588]),
			.SE(gen[7589]),

			.SELF(gen[7493]),
			.cell_state(gen[7493])
		); 

/******************* CELL 7494 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7494 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7398]),
			.N(gen[7399]),
			.NE(gen[7400]),

			.O(gen[7493]),
			.E(gen[7495]),

			.SO(gen[7588]),
			.S(gen[7589]),
			.SE(gen[7590]),

			.SELF(gen[7494]),
			.cell_state(gen[7494])
		); 

/******************* CELL 7495 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7495 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7399]),
			.N(gen[7400]),
			.NE(gen[7401]),

			.O(gen[7494]),
			.E(gen[7496]),

			.SO(gen[7589]),
			.S(gen[7590]),
			.SE(gen[7591]),

			.SELF(gen[7495]),
			.cell_state(gen[7495])
		); 

/******************* CELL 7496 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7496 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7400]),
			.N(gen[7401]),
			.NE(gen[7402]),

			.O(gen[7495]),
			.E(gen[7497]),

			.SO(gen[7590]),
			.S(gen[7591]),
			.SE(gen[7592]),

			.SELF(gen[7496]),
			.cell_state(gen[7496])
		); 

/******************* CELL 7497 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7497 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7401]),
			.N(gen[7402]),
			.NE(gen[7403]),

			.O(gen[7496]),
			.E(gen[7498]),

			.SO(gen[7591]),
			.S(gen[7592]),
			.SE(gen[7593]),

			.SELF(gen[7497]),
			.cell_state(gen[7497])
		); 

/******************* CELL 7498 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7498 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7402]),
			.N(gen[7403]),
			.NE(gen[7404]),

			.O(gen[7497]),
			.E(gen[7499]),

			.SO(gen[7592]),
			.S(gen[7593]),
			.SE(gen[7594]),

			.SELF(gen[7498]),
			.cell_state(gen[7498])
		); 

/******************* CELL 7499 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7499 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7403]),
			.N(gen[7404]),
			.NE(gen[7405]),

			.O(gen[7498]),
			.E(gen[7500]),

			.SO(gen[7593]),
			.S(gen[7594]),
			.SE(gen[7595]),

			.SELF(gen[7499]),
			.cell_state(gen[7499])
		); 

/******************* CELL 7500 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7500 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7404]),
			.N(gen[7405]),
			.NE(gen[7406]),

			.O(gen[7499]),
			.E(gen[7501]),

			.SO(gen[7594]),
			.S(gen[7595]),
			.SE(gen[7596]),

			.SELF(gen[7500]),
			.cell_state(gen[7500])
		); 

/******************* CELL 7501 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7501 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7405]),
			.N(gen[7406]),
			.NE(gen[7407]),

			.O(gen[7500]),
			.E(gen[7502]),

			.SO(gen[7595]),
			.S(gen[7596]),
			.SE(gen[7597]),

			.SELF(gen[7501]),
			.cell_state(gen[7501])
		); 

/******************* CELL 7502 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7502 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7406]),
			.N(gen[7407]),
			.NE(gen[7408]),

			.O(gen[7501]),
			.E(gen[7503]),

			.SO(gen[7596]),
			.S(gen[7597]),
			.SE(gen[7598]),

			.SELF(gen[7502]),
			.cell_state(gen[7502])
		); 

/******************* CELL 7503 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7503 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7407]),
			.N(gen[7408]),
			.NE(gen[7409]),

			.O(gen[7502]),
			.E(gen[7504]),

			.SO(gen[7597]),
			.S(gen[7598]),
			.SE(gen[7599]),

			.SELF(gen[7503]),
			.cell_state(gen[7503])
		); 

/******************* CELL 7504 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7504 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7408]),
			.N(gen[7409]),
			.NE(gen[7408]),

			.O(gen[7503]),
			.E(gen[7503]),

			.SO(gen[7598]),
			.S(gen[7599]),
			.SE(gen[7598]),

			.SELF(gen[7504]),
			.cell_state(gen[7504])
		); 

/******************* CELL 7505 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7505 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7411]),
			.N(gen[7410]),
			.NE(gen[7411]),

			.O(gen[7506]),
			.E(gen[7506]),

			.SO(gen[7601]),
			.S(gen[7600]),
			.SE(gen[7601]),

			.SELF(gen[7505]),
			.cell_state(gen[7505])
		); 

/******************* CELL 7506 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7506 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7410]),
			.N(gen[7411]),
			.NE(gen[7412]),

			.O(gen[7505]),
			.E(gen[7507]),

			.SO(gen[7600]),
			.S(gen[7601]),
			.SE(gen[7602]),

			.SELF(gen[7506]),
			.cell_state(gen[7506])
		); 

/******************* CELL 7507 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7507 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7411]),
			.N(gen[7412]),
			.NE(gen[7413]),

			.O(gen[7506]),
			.E(gen[7508]),

			.SO(gen[7601]),
			.S(gen[7602]),
			.SE(gen[7603]),

			.SELF(gen[7507]),
			.cell_state(gen[7507])
		); 

/******************* CELL 7508 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7508 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7412]),
			.N(gen[7413]),
			.NE(gen[7414]),

			.O(gen[7507]),
			.E(gen[7509]),

			.SO(gen[7602]),
			.S(gen[7603]),
			.SE(gen[7604]),

			.SELF(gen[7508]),
			.cell_state(gen[7508])
		); 

/******************* CELL 7509 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7509 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7413]),
			.N(gen[7414]),
			.NE(gen[7415]),

			.O(gen[7508]),
			.E(gen[7510]),

			.SO(gen[7603]),
			.S(gen[7604]),
			.SE(gen[7605]),

			.SELF(gen[7509]),
			.cell_state(gen[7509])
		); 

/******************* CELL 7510 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7510 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7414]),
			.N(gen[7415]),
			.NE(gen[7416]),

			.O(gen[7509]),
			.E(gen[7511]),

			.SO(gen[7604]),
			.S(gen[7605]),
			.SE(gen[7606]),

			.SELF(gen[7510]),
			.cell_state(gen[7510])
		); 

/******************* CELL 7511 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7511 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7415]),
			.N(gen[7416]),
			.NE(gen[7417]),

			.O(gen[7510]),
			.E(gen[7512]),

			.SO(gen[7605]),
			.S(gen[7606]),
			.SE(gen[7607]),

			.SELF(gen[7511]),
			.cell_state(gen[7511])
		); 

/******************* CELL 7512 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7512 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7416]),
			.N(gen[7417]),
			.NE(gen[7418]),

			.O(gen[7511]),
			.E(gen[7513]),

			.SO(gen[7606]),
			.S(gen[7607]),
			.SE(gen[7608]),

			.SELF(gen[7512]),
			.cell_state(gen[7512])
		); 

/******************* CELL 7513 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7513 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7417]),
			.N(gen[7418]),
			.NE(gen[7419]),

			.O(gen[7512]),
			.E(gen[7514]),

			.SO(gen[7607]),
			.S(gen[7608]),
			.SE(gen[7609]),

			.SELF(gen[7513]),
			.cell_state(gen[7513])
		); 

/******************* CELL 7514 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7514 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7418]),
			.N(gen[7419]),
			.NE(gen[7420]),

			.O(gen[7513]),
			.E(gen[7515]),

			.SO(gen[7608]),
			.S(gen[7609]),
			.SE(gen[7610]),

			.SELF(gen[7514]),
			.cell_state(gen[7514])
		); 

/******************* CELL 7515 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7515 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7419]),
			.N(gen[7420]),
			.NE(gen[7421]),

			.O(gen[7514]),
			.E(gen[7516]),

			.SO(gen[7609]),
			.S(gen[7610]),
			.SE(gen[7611]),

			.SELF(gen[7515]),
			.cell_state(gen[7515])
		); 

/******************* CELL 7516 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7516 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7420]),
			.N(gen[7421]),
			.NE(gen[7422]),

			.O(gen[7515]),
			.E(gen[7517]),

			.SO(gen[7610]),
			.S(gen[7611]),
			.SE(gen[7612]),

			.SELF(gen[7516]),
			.cell_state(gen[7516])
		); 

/******************* CELL 7517 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7517 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7421]),
			.N(gen[7422]),
			.NE(gen[7423]),

			.O(gen[7516]),
			.E(gen[7518]),

			.SO(gen[7611]),
			.S(gen[7612]),
			.SE(gen[7613]),

			.SELF(gen[7517]),
			.cell_state(gen[7517])
		); 

/******************* CELL 7518 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7518 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7422]),
			.N(gen[7423]),
			.NE(gen[7424]),

			.O(gen[7517]),
			.E(gen[7519]),

			.SO(gen[7612]),
			.S(gen[7613]),
			.SE(gen[7614]),

			.SELF(gen[7518]),
			.cell_state(gen[7518])
		); 

/******************* CELL 7519 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7519 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7423]),
			.N(gen[7424]),
			.NE(gen[7425]),

			.O(gen[7518]),
			.E(gen[7520]),

			.SO(gen[7613]),
			.S(gen[7614]),
			.SE(gen[7615]),

			.SELF(gen[7519]),
			.cell_state(gen[7519])
		); 

/******************* CELL 7520 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7520 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7424]),
			.N(gen[7425]),
			.NE(gen[7426]),

			.O(gen[7519]),
			.E(gen[7521]),

			.SO(gen[7614]),
			.S(gen[7615]),
			.SE(gen[7616]),

			.SELF(gen[7520]),
			.cell_state(gen[7520])
		); 

/******************* CELL 7521 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7521 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7425]),
			.N(gen[7426]),
			.NE(gen[7427]),

			.O(gen[7520]),
			.E(gen[7522]),

			.SO(gen[7615]),
			.S(gen[7616]),
			.SE(gen[7617]),

			.SELF(gen[7521]),
			.cell_state(gen[7521])
		); 

/******************* CELL 7522 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7522 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7426]),
			.N(gen[7427]),
			.NE(gen[7428]),

			.O(gen[7521]),
			.E(gen[7523]),

			.SO(gen[7616]),
			.S(gen[7617]),
			.SE(gen[7618]),

			.SELF(gen[7522]),
			.cell_state(gen[7522])
		); 

/******************* CELL 7523 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7523 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7427]),
			.N(gen[7428]),
			.NE(gen[7429]),

			.O(gen[7522]),
			.E(gen[7524]),

			.SO(gen[7617]),
			.S(gen[7618]),
			.SE(gen[7619]),

			.SELF(gen[7523]),
			.cell_state(gen[7523])
		); 

/******************* CELL 7524 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7524 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7428]),
			.N(gen[7429]),
			.NE(gen[7430]),

			.O(gen[7523]),
			.E(gen[7525]),

			.SO(gen[7618]),
			.S(gen[7619]),
			.SE(gen[7620]),

			.SELF(gen[7524]),
			.cell_state(gen[7524])
		); 

/******************* CELL 7525 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7525 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7429]),
			.N(gen[7430]),
			.NE(gen[7431]),

			.O(gen[7524]),
			.E(gen[7526]),

			.SO(gen[7619]),
			.S(gen[7620]),
			.SE(gen[7621]),

			.SELF(gen[7525]),
			.cell_state(gen[7525])
		); 

/******************* CELL 7526 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7526 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7430]),
			.N(gen[7431]),
			.NE(gen[7432]),

			.O(gen[7525]),
			.E(gen[7527]),

			.SO(gen[7620]),
			.S(gen[7621]),
			.SE(gen[7622]),

			.SELF(gen[7526]),
			.cell_state(gen[7526])
		); 

/******************* CELL 7527 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7527 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7431]),
			.N(gen[7432]),
			.NE(gen[7433]),

			.O(gen[7526]),
			.E(gen[7528]),

			.SO(gen[7621]),
			.S(gen[7622]),
			.SE(gen[7623]),

			.SELF(gen[7527]),
			.cell_state(gen[7527])
		); 

/******************* CELL 7528 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7528 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7432]),
			.N(gen[7433]),
			.NE(gen[7434]),

			.O(gen[7527]),
			.E(gen[7529]),

			.SO(gen[7622]),
			.S(gen[7623]),
			.SE(gen[7624]),

			.SELF(gen[7528]),
			.cell_state(gen[7528])
		); 

/******************* CELL 7529 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7529 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7433]),
			.N(gen[7434]),
			.NE(gen[7435]),

			.O(gen[7528]),
			.E(gen[7530]),

			.SO(gen[7623]),
			.S(gen[7624]),
			.SE(gen[7625]),

			.SELF(gen[7529]),
			.cell_state(gen[7529])
		); 

/******************* CELL 7530 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7530 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7434]),
			.N(gen[7435]),
			.NE(gen[7436]),

			.O(gen[7529]),
			.E(gen[7531]),

			.SO(gen[7624]),
			.S(gen[7625]),
			.SE(gen[7626]),

			.SELF(gen[7530]),
			.cell_state(gen[7530])
		); 

/******************* CELL 7531 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7531 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7435]),
			.N(gen[7436]),
			.NE(gen[7437]),

			.O(gen[7530]),
			.E(gen[7532]),

			.SO(gen[7625]),
			.S(gen[7626]),
			.SE(gen[7627]),

			.SELF(gen[7531]),
			.cell_state(gen[7531])
		); 

/******************* CELL 7532 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7532 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7436]),
			.N(gen[7437]),
			.NE(gen[7438]),

			.O(gen[7531]),
			.E(gen[7533]),

			.SO(gen[7626]),
			.S(gen[7627]),
			.SE(gen[7628]),

			.SELF(gen[7532]),
			.cell_state(gen[7532])
		); 

/******************* CELL 7533 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7533 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7437]),
			.N(gen[7438]),
			.NE(gen[7439]),

			.O(gen[7532]),
			.E(gen[7534]),

			.SO(gen[7627]),
			.S(gen[7628]),
			.SE(gen[7629]),

			.SELF(gen[7533]),
			.cell_state(gen[7533])
		); 

/******************* CELL 7534 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7534 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7438]),
			.N(gen[7439]),
			.NE(gen[7440]),

			.O(gen[7533]),
			.E(gen[7535]),

			.SO(gen[7628]),
			.S(gen[7629]),
			.SE(gen[7630]),

			.SELF(gen[7534]),
			.cell_state(gen[7534])
		); 

/******************* CELL 7535 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7535 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7439]),
			.N(gen[7440]),
			.NE(gen[7441]),

			.O(gen[7534]),
			.E(gen[7536]),

			.SO(gen[7629]),
			.S(gen[7630]),
			.SE(gen[7631]),

			.SELF(gen[7535]),
			.cell_state(gen[7535])
		); 

/******************* CELL 7536 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7536 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7440]),
			.N(gen[7441]),
			.NE(gen[7442]),

			.O(gen[7535]),
			.E(gen[7537]),

			.SO(gen[7630]),
			.S(gen[7631]),
			.SE(gen[7632]),

			.SELF(gen[7536]),
			.cell_state(gen[7536])
		); 

/******************* CELL 7537 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7537 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7441]),
			.N(gen[7442]),
			.NE(gen[7443]),

			.O(gen[7536]),
			.E(gen[7538]),

			.SO(gen[7631]),
			.S(gen[7632]),
			.SE(gen[7633]),

			.SELF(gen[7537]),
			.cell_state(gen[7537])
		); 

/******************* CELL 7538 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7538 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7442]),
			.N(gen[7443]),
			.NE(gen[7444]),

			.O(gen[7537]),
			.E(gen[7539]),

			.SO(gen[7632]),
			.S(gen[7633]),
			.SE(gen[7634]),

			.SELF(gen[7538]),
			.cell_state(gen[7538])
		); 

/******************* CELL 7539 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7539 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7443]),
			.N(gen[7444]),
			.NE(gen[7445]),

			.O(gen[7538]),
			.E(gen[7540]),

			.SO(gen[7633]),
			.S(gen[7634]),
			.SE(gen[7635]),

			.SELF(gen[7539]),
			.cell_state(gen[7539])
		); 

/******************* CELL 7540 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7540 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7444]),
			.N(gen[7445]),
			.NE(gen[7446]),

			.O(gen[7539]),
			.E(gen[7541]),

			.SO(gen[7634]),
			.S(gen[7635]),
			.SE(gen[7636]),

			.SELF(gen[7540]),
			.cell_state(gen[7540])
		); 

/******************* CELL 7541 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7541 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7445]),
			.N(gen[7446]),
			.NE(gen[7447]),

			.O(gen[7540]),
			.E(gen[7542]),

			.SO(gen[7635]),
			.S(gen[7636]),
			.SE(gen[7637]),

			.SELF(gen[7541]),
			.cell_state(gen[7541])
		); 

/******************* CELL 7542 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7542 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7446]),
			.N(gen[7447]),
			.NE(gen[7448]),

			.O(gen[7541]),
			.E(gen[7543]),

			.SO(gen[7636]),
			.S(gen[7637]),
			.SE(gen[7638]),

			.SELF(gen[7542]),
			.cell_state(gen[7542])
		); 

/******************* CELL 7543 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7543 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7447]),
			.N(gen[7448]),
			.NE(gen[7449]),

			.O(gen[7542]),
			.E(gen[7544]),

			.SO(gen[7637]),
			.S(gen[7638]),
			.SE(gen[7639]),

			.SELF(gen[7543]),
			.cell_state(gen[7543])
		); 

/******************* CELL 7544 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7544 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7448]),
			.N(gen[7449]),
			.NE(gen[7450]),

			.O(gen[7543]),
			.E(gen[7545]),

			.SO(gen[7638]),
			.S(gen[7639]),
			.SE(gen[7640]),

			.SELF(gen[7544]),
			.cell_state(gen[7544])
		); 

/******************* CELL 7545 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7545 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7449]),
			.N(gen[7450]),
			.NE(gen[7451]),

			.O(gen[7544]),
			.E(gen[7546]),

			.SO(gen[7639]),
			.S(gen[7640]),
			.SE(gen[7641]),

			.SELF(gen[7545]),
			.cell_state(gen[7545])
		); 

/******************* CELL 7546 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7546 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7450]),
			.N(gen[7451]),
			.NE(gen[7452]),

			.O(gen[7545]),
			.E(gen[7547]),

			.SO(gen[7640]),
			.S(gen[7641]),
			.SE(gen[7642]),

			.SELF(gen[7546]),
			.cell_state(gen[7546])
		); 

/******************* CELL 7547 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7547 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7451]),
			.N(gen[7452]),
			.NE(gen[7453]),

			.O(gen[7546]),
			.E(gen[7548]),

			.SO(gen[7641]),
			.S(gen[7642]),
			.SE(gen[7643]),

			.SELF(gen[7547]),
			.cell_state(gen[7547])
		); 

/******************* CELL 7548 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7548 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7452]),
			.N(gen[7453]),
			.NE(gen[7454]),

			.O(gen[7547]),
			.E(gen[7549]),

			.SO(gen[7642]),
			.S(gen[7643]),
			.SE(gen[7644]),

			.SELF(gen[7548]),
			.cell_state(gen[7548])
		); 

/******************* CELL 7549 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7549 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7453]),
			.N(gen[7454]),
			.NE(gen[7455]),

			.O(gen[7548]),
			.E(gen[7550]),

			.SO(gen[7643]),
			.S(gen[7644]),
			.SE(gen[7645]),

			.SELF(gen[7549]),
			.cell_state(gen[7549])
		); 

/******************* CELL 7550 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7550 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7454]),
			.N(gen[7455]),
			.NE(gen[7456]),

			.O(gen[7549]),
			.E(gen[7551]),

			.SO(gen[7644]),
			.S(gen[7645]),
			.SE(gen[7646]),

			.SELF(gen[7550]),
			.cell_state(gen[7550])
		); 

/******************* CELL 7551 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7551 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7455]),
			.N(gen[7456]),
			.NE(gen[7457]),

			.O(gen[7550]),
			.E(gen[7552]),

			.SO(gen[7645]),
			.S(gen[7646]),
			.SE(gen[7647]),

			.SELF(gen[7551]),
			.cell_state(gen[7551])
		); 

/******************* CELL 7552 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7552 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7456]),
			.N(gen[7457]),
			.NE(gen[7458]),

			.O(gen[7551]),
			.E(gen[7553]),

			.SO(gen[7646]),
			.S(gen[7647]),
			.SE(gen[7648]),

			.SELF(gen[7552]),
			.cell_state(gen[7552])
		); 

/******************* CELL 7553 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7553 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7457]),
			.N(gen[7458]),
			.NE(gen[7459]),

			.O(gen[7552]),
			.E(gen[7554]),

			.SO(gen[7647]),
			.S(gen[7648]),
			.SE(gen[7649]),

			.SELF(gen[7553]),
			.cell_state(gen[7553])
		); 

/******************* CELL 7554 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7554 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7458]),
			.N(gen[7459]),
			.NE(gen[7460]),

			.O(gen[7553]),
			.E(gen[7555]),

			.SO(gen[7648]),
			.S(gen[7649]),
			.SE(gen[7650]),

			.SELF(gen[7554]),
			.cell_state(gen[7554])
		); 

/******************* CELL 7555 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7555 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7459]),
			.N(gen[7460]),
			.NE(gen[7461]),

			.O(gen[7554]),
			.E(gen[7556]),

			.SO(gen[7649]),
			.S(gen[7650]),
			.SE(gen[7651]),

			.SELF(gen[7555]),
			.cell_state(gen[7555])
		); 

/******************* CELL 7556 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7556 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7460]),
			.N(gen[7461]),
			.NE(gen[7462]),

			.O(gen[7555]),
			.E(gen[7557]),

			.SO(gen[7650]),
			.S(gen[7651]),
			.SE(gen[7652]),

			.SELF(gen[7556]),
			.cell_state(gen[7556])
		); 

/******************* CELL 7557 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7557 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7461]),
			.N(gen[7462]),
			.NE(gen[7463]),

			.O(gen[7556]),
			.E(gen[7558]),

			.SO(gen[7651]),
			.S(gen[7652]),
			.SE(gen[7653]),

			.SELF(gen[7557]),
			.cell_state(gen[7557])
		); 

/******************* CELL 7558 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7558 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7462]),
			.N(gen[7463]),
			.NE(gen[7464]),

			.O(gen[7557]),
			.E(gen[7559]),

			.SO(gen[7652]),
			.S(gen[7653]),
			.SE(gen[7654]),

			.SELF(gen[7558]),
			.cell_state(gen[7558])
		); 

/******************* CELL 7559 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7559 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7463]),
			.N(gen[7464]),
			.NE(gen[7465]),

			.O(gen[7558]),
			.E(gen[7560]),

			.SO(gen[7653]),
			.S(gen[7654]),
			.SE(gen[7655]),

			.SELF(gen[7559]),
			.cell_state(gen[7559])
		); 

/******************* CELL 7560 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7560 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7464]),
			.N(gen[7465]),
			.NE(gen[7466]),

			.O(gen[7559]),
			.E(gen[7561]),

			.SO(gen[7654]),
			.S(gen[7655]),
			.SE(gen[7656]),

			.SELF(gen[7560]),
			.cell_state(gen[7560])
		); 

/******************* CELL 7561 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7561 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7465]),
			.N(gen[7466]),
			.NE(gen[7467]),

			.O(gen[7560]),
			.E(gen[7562]),

			.SO(gen[7655]),
			.S(gen[7656]),
			.SE(gen[7657]),

			.SELF(gen[7561]),
			.cell_state(gen[7561])
		); 

/******************* CELL 7562 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7562 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7466]),
			.N(gen[7467]),
			.NE(gen[7468]),

			.O(gen[7561]),
			.E(gen[7563]),

			.SO(gen[7656]),
			.S(gen[7657]),
			.SE(gen[7658]),

			.SELF(gen[7562]),
			.cell_state(gen[7562])
		); 

/******************* CELL 7563 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7563 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7467]),
			.N(gen[7468]),
			.NE(gen[7469]),

			.O(gen[7562]),
			.E(gen[7564]),

			.SO(gen[7657]),
			.S(gen[7658]),
			.SE(gen[7659]),

			.SELF(gen[7563]),
			.cell_state(gen[7563])
		); 

/******************* CELL 7564 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7564 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7468]),
			.N(gen[7469]),
			.NE(gen[7470]),

			.O(gen[7563]),
			.E(gen[7565]),

			.SO(gen[7658]),
			.S(gen[7659]),
			.SE(gen[7660]),

			.SELF(gen[7564]),
			.cell_state(gen[7564])
		); 

/******************* CELL 7565 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7565 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7469]),
			.N(gen[7470]),
			.NE(gen[7471]),

			.O(gen[7564]),
			.E(gen[7566]),

			.SO(gen[7659]),
			.S(gen[7660]),
			.SE(gen[7661]),

			.SELF(gen[7565]),
			.cell_state(gen[7565])
		); 

/******************* CELL 7566 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7566 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7470]),
			.N(gen[7471]),
			.NE(gen[7472]),

			.O(gen[7565]),
			.E(gen[7567]),

			.SO(gen[7660]),
			.S(gen[7661]),
			.SE(gen[7662]),

			.SELF(gen[7566]),
			.cell_state(gen[7566])
		); 

/******************* CELL 7567 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7567 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7471]),
			.N(gen[7472]),
			.NE(gen[7473]),

			.O(gen[7566]),
			.E(gen[7568]),

			.SO(gen[7661]),
			.S(gen[7662]),
			.SE(gen[7663]),

			.SELF(gen[7567]),
			.cell_state(gen[7567])
		); 

/******************* CELL 7568 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7568 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7472]),
			.N(gen[7473]),
			.NE(gen[7474]),

			.O(gen[7567]),
			.E(gen[7569]),

			.SO(gen[7662]),
			.S(gen[7663]),
			.SE(gen[7664]),

			.SELF(gen[7568]),
			.cell_state(gen[7568])
		); 

/******************* CELL 7569 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7569 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7473]),
			.N(gen[7474]),
			.NE(gen[7475]),

			.O(gen[7568]),
			.E(gen[7570]),

			.SO(gen[7663]),
			.S(gen[7664]),
			.SE(gen[7665]),

			.SELF(gen[7569]),
			.cell_state(gen[7569])
		); 

/******************* CELL 7570 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7570 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7474]),
			.N(gen[7475]),
			.NE(gen[7476]),

			.O(gen[7569]),
			.E(gen[7571]),

			.SO(gen[7664]),
			.S(gen[7665]),
			.SE(gen[7666]),

			.SELF(gen[7570]),
			.cell_state(gen[7570])
		); 

/******************* CELL 7571 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7571 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7475]),
			.N(gen[7476]),
			.NE(gen[7477]),

			.O(gen[7570]),
			.E(gen[7572]),

			.SO(gen[7665]),
			.S(gen[7666]),
			.SE(gen[7667]),

			.SELF(gen[7571]),
			.cell_state(gen[7571])
		); 

/******************* CELL 7572 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7572 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7476]),
			.N(gen[7477]),
			.NE(gen[7478]),

			.O(gen[7571]),
			.E(gen[7573]),

			.SO(gen[7666]),
			.S(gen[7667]),
			.SE(gen[7668]),

			.SELF(gen[7572]),
			.cell_state(gen[7572])
		); 

/******************* CELL 7573 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7573 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7477]),
			.N(gen[7478]),
			.NE(gen[7479]),

			.O(gen[7572]),
			.E(gen[7574]),

			.SO(gen[7667]),
			.S(gen[7668]),
			.SE(gen[7669]),

			.SELF(gen[7573]),
			.cell_state(gen[7573])
		); 

/******************* CELL 7574 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7574 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7478]),
			.N(gen[7479]),
			.NE(gen[7480]),

			.O(gen[7573]),
			.E(gen[7575]),

			.SO(gen[7668]),
			.S(gen[7669]),
			.SE(gen[7670]),

			.SELF(gen[7574]),
			.cell_state(gen[7574])
		); 

/******************* CELL 7575 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7575 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7479]),
			.N(gen[7480]),
			.NE(gen[7481]),

			.O(gen[7574]),
			.E(gen[7576]),

			.SO(gen[7669]),
			.S(gen[7670]),
			.SE(gen[7671]),

			.SELF(gen[7575]),
			.cell_state(gen[7575])
		); 

/******************* CELL 7576 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7576 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7480]),
			.N(gen[7481]),
			.NE(gen[7482]),

			.O(gen[7575]),
			.E(gen[7577]),

			.SO(gen[7670]),
			.S(gen[7671]),
			.SE(gen[7672]),

			.SELF(gen[7576]),
			.cell_state(gen[7576])
		); 

/******************* CELL 7577 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7577 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7481]),
			.N(gen[7482]),
			.NE(gen[7483]),

			.O(gen[7576]),
			.E(gen[7578]),

			.SO(gen[7671]),
			.S(gen[7672]),
			.SE(gen[7673]),

			.SELF(gen[7577]),
			.cell_state(gen[7577])
		); 

/******************* CELL 7578 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7578 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7482]),
			.N(gen[7483]),
			.NE(gen[7484]),

			.O(gen[7577]),
			.E(gen[7579]),

			.SO(gen[7672]),
			.S(gen[7673]),
			.SE(gen[7674]),

			.SELF(gen[7578]),
			.cell_state(gen[7578])
		); 

/******************* CELL 7579 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7579 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7483]),
			.N(gen[7484]),
			.NE(gen[7485]),

			.O(gen[7578]),
			.E(gen[7580]),

			.SO(gen[7673]),
			.S(gen[7674]),
			.SE(gen[7675]),

			.SELF(gen[7579]),
			.cell_state(gen[7579])
		); 

/******************* CELL 7580 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7580 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7484]),
			.N(gen[7485]),
			.NE(gen[7486]),

			.O(gen[7579]),
			.E(gen[7581]),

			.SO(gen[7674]),
			.S(gen[7675]),
			.SE(gen[7676]),

			.SELF(gen[7580]),
			.cell_state(gen[7580])
		); 

/******************* CELL 7581 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7581 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7485]),
			.N(gen[7486]),
			.NE(gen[7487]),

			.O(gen[7580]),
			.E(gen[7582]),

			.SO(gen[7675]),
			.S(gen[7676]),
			.SE(gen[7677]),

			.SELF(gen[7581]),
			.cell_state(gen[7581])
		); 

/******************* CELL 7582 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7582 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7486]),
			.N(gen[7487]),
			.NE(gen[7488]),

			.O(gen[7581]),
			.E(gen[7583]),

			.SO(gen[7676]),
			.S(gen[7677]),
			.SE(gen[7678]),

			.SELF(gen[7582]),
			.cell_state(gen[7582])
		); 

/******************* CELL 7583 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7583 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7487]),
			.N(gen[7488]),
			.NE(gen[7489]),

			.O(gen[7582]),
			.E(gen[7584]),

			.SO(gen[7677]),
			.S(gen[7678]),
			.SE(gen[7679]),

			.SELF(gen[7583]),
			.cell_state(gen[7583])
		); 

/******************* CELL 7584 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7584 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7488]),
			.N(gen[7489]),
			.NE(gen[7490]),

			.O(gen[7583]),
			.E(gen[7585]),

			.SO(gen[7678]),
			.S(gen[7679]),
			.SE(gen[7680]),

			.SELF(gen[7584]),
			.cell_state(gen[7584])
		); 

/******************* CELL 7585 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7585 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7489]),
			.N(gen[7490]),
			.NE(gen[7491]),

			.O(gen[7584]),
			.E(gen[7586]),

			.SO(gen[7679]),
			.S(gen[7680]),
			.SE(gen[7681]),

			.SELF(gen[7585]),
			.cell_state(gen[7585])
		); 

/******************* CELL 7586 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7586 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7490]),
			.N(gen[7491]),
			.NE(gen[7492]),

			.O(gen[7585]),
			.E(gen[7587]),

			.SO(gen[7680]),
			.S(gen[7681]),
			.SE(gen[7682]),

			.SELF(gen[7586]),
			.cell_state(gen[7586])
		); 

/******************* CELL 7587 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7587 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7491]),
			.N(gen[7492]),
			.NE(gen[7493]),

			.O(gen[7586]),
			.E(gen[7588]),

			.SO(gen[7681]),
			.S(gen[7682]),
			.SE(gen[7683]),

			.SELF(gen[7587]),
			.cell_state(gen[7587])
		); 

/******************* CELL 7588 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7588 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7492]),
			.N(gen[7493]),
			.NE(gen[7494]),

			.O(gen[7587]),
			.E(gen[7589]),

			.SO(gen[7682]),
			.S(gen[7683]),
			.SE(gen[7684]),

			.SELF(gen[7588]),
			.cell_state(gen[7588])
		); 

/******************* CELL 7589 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7589 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7493]),
			.N(gen[7494]),
			.NE(gen[7495]),

			.O(gen[7588]),
			.E(gen[7590]),

			.SO(gen[7683]),
			.S(gen[7684]),
			.SE(gen[7685]),

			.SELF(gen[7589]),
			.cell_state(gen[7589])
		); 

/******************* CELL 7590 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7590 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7494]),
			.N(gen[7495]),
			.NE(gen[7496]),

			.O(gen[7589]),
			.E(gen[7591]),

			.SO(gen[7684]),
			.S(gen[7685]),
			.SE(gen[7686]),

			.SELF(gen[7590]),
			.cell_state(gen[7590])
		); 

/******************* CELL 7591 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7591 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7495]),
			.N(gen[7496]),
			.NE(gen[7497]),

			.O(gen[7590]),
			.E(gen[7592]),

			.SO(gen[7685]),
			.S(gen[7686]),
			.SE(gen[7687]),

			.SELF(gen[7591]),
			.cell_state(gen[7591])
		); 

/******************* CELL 7592 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7592 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7496]),
			.N(gen[7497]),
			.NE(gen[7498]),

			.O(gen[7591]),
			.E(gen[7593]),

			.SO(gen[7686]),
			.S(gen[7687]),
			.SE(gen[7688]),

			.SELF(gen[7592]),
			.cell_state(gen[7592])
		); 

/******************* CELL 7593 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7593 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7497]),
			.N(gen[7498]),
			.NE(gen[7499]),

			.O(gen[7592]),
			.E(gen[7594]),

			.SO(gen[7687]),
			.S(gen[7688]),
			.SE(gen[7689]),

			.SELF(gen[7593]),
			.cell_state(gen[7593])
		); 

/******************* CELL 7594 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7594 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7498]),
			.N(gen[7499]),
			.NE(gen[7500]),

			.O(gen[7593]),
			.E(gen[7595]),

			.SO(gen[7688]),
			.S(gen[7689]),
			.SE(gen[7690]),

			.SELF(gen[7594]),
			.cell_state(gen[7594])
		); 

/******************* CELL 7595 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7595 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7499]),
			.N(gen[7500]),
			.NE(gen[7501]),

			.O(gen[7594]),
			.E(gen[7596]),

			.SO(gen[7689]),
			.S(gen[7690]),
			.SE(gen[7691]),

			.SELF(gen[7595]),
			.cell_state(gen[7595])
		); 

/******************* CELL 7596 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7596 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7500]),
			.N(gen[7501]),
			.NE(gen[7502]),

			.O(gen[7595]),
			.E(gen[7597]),

			.SO(gen[7690]),
			.S(gen[7691]),
			.SE(gen[7692]),

			.SELF(gen[7596]),
			.cell_state(gen[7596])
		); 

/******************* CELL 7597 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7597 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7501]),
			.N(gen[7502]),
			.NE(gen[7503]),

			.O(gen[7596]),
			.E(gen[7598]),

			.SO(gen[7691]),
			.S(gen[7692]),
			.SE(gen[7693]),

			.SELF(gen[7597]),
			.cell_state(gen[7597])
		); 

/******************* CELL 7598 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7598 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7502]),
			.N(gen[7503]),
			.NE(gen[7504]),

			.O(gen[7597]),
			.E(gen[7599]),

			.SO(gen[7692]),
			.S(gen[7693]),
			.SE(gen[7694]),

			.SELF(gen[7598]),
			.cell_state(gen[7598])
		); 

/******************* CELL 7599 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7599 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7503]),
			.N(gen[7504]),
			.NE(gen[7503]),

			.O(gen[7598]),
			.E(gen[7598]),

			.SO(gen[7693]),
			.S(gen[7694]),
			.SE(gen[7693]),

			.SELF(gen[7599]),
			.cell_state(gen[7599])
		); 

/******************* CELL 7600 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7600 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7506]),
			.N(gen[7505]),
			.NE(gen[7506]),

			.O(gen[7601]),
			.E(gen[7601]),

			.SO(gen[7696]),
			.S(gen[7695]),
			.SE(gen[7696]),

			.SELF(gen[7600]),
			.cell_state(gen[7600])
		); 

/******************* CELL 7601 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7601 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7505]),
			.N(gen[7506]),
			.NE(gen[7507]),

			.O(gen[7600]),
			.E(gen[7602]),

			.SO(gen[7695]),
			.S(gen[7696]),
			.SE(gen[7697]),

			.SELF(gen[7601]),
			.cell_state(gen[7601])
		); 

/******************* CELL 7602 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7602 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7506]),
			.N(gen[7507]),
			.NE(gen[7508]),

			.O(gen[7601]),
			.E(gen[7603]),

			.SO(gen[7696]),
			.S(gen[7697]),
			.SE(gen[7698]),

			.SELF(gen[7602]),
			.cell_state(gen[7602])
		); 

/******************* CELL 7603 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7603 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7507]),
			.N(gen[7508]),
			.NE(gen[7509]),

			.O(gen[7602]),
			.E(gen[7604]),

			.SO(gen[7697]),
			.S(gen[7698]),
			.SE(gen[7699]),

			.SELF(gen[7603]),
			.cell_state(gen[7603])
		); 

/******************* CELL 7604 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7604 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7508]),
			.N(gen[7509]),
			.NE(gen[7510]),

			.O(gen[7603]),
			.E(gen[7605]),

			.SO(gen[7698]),
			.S(gen[7699]),
			.SE(gen[7700]),

			.SELF(gen[7604]),
			.cell_state(gen[7604])
		); 

/******************* CELL 7605 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7605 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7509]),
			.N(gen[7510]),
			.NE(gen[7511]),

			.O(gen[7604]),
			.E(gen[7606]),

			.SO(gen[7699]),
			.S(gen[7700]),
			.SE(gen[7701]),

			.SELF(gen[7605]),
			.cell_state(gen[7605])
		); 

/******************* CELL 7606 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7606 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7510]),
			.N(gen[7511]),
			.NE(gen[7512]),

			.O(gen[7605]),
			.E(gen[7607]),

			.SO(gen[7700]),
			.S(gen[7701]),
			.SE(gen[7702]),

			.SELF(gen[7606]),
			.cell_state(gen[7606])
		); 

/******************* CELL 7607 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7607 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7511]),
			.N(gen[7512]),
			.NE(gen[7513]),

			.O(gen[7606]),
			.E(gen[7608]),

			.SO(gen[7701]),
			.S(gen[7702]),
			.SE(gen[7703]),

			.SELF(gen[7607]),
			.cell_state(gen[7607])
		); 

/******************* CELL 7608 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7608 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7512]),
			.N(gen[7513]),
			.NE(gen[7514]),

			.O(gen[7607]),
			.E(gen[7609]),

			.SO(gen[7702]),
			.S(gen[7703]),
			.SE(gen[7704]),

			.SELF(gen[7608]),
			.cell_state(gen[7608])
		); 

/******************* CELL 7609 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7609 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7513]),
			.N(gen[7514]),
			.NE(gen[7515]),

			.O(gen[7608]),
			.E(gen[7610]),

			.SO(gen[7703]),
			.S(gen[7704]),
			.SE(gen[7705]),

			.SELF(gen[7609]),
			.cell_state(gen[7609])
		); 

/******************* CELL 7610 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7610 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7514]),
			.N(gen[7515]),
			.NE(gen[7516]),

			.O(gen[7609]),
			.E(gen[7611]),

			.SO(gen[7704]),
			.S(gen[7705]),
			.SE(gen[7706]),

			.SELF(gen[7610]),
			.cell_state(gen[7610])
		); 

/******************* CELL 7611 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7611 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7515]),
			.N(gen[7516]),
			.NE(gen[7517]),

			.O(gen[7610]),
			.E(gen[7612]),

			.SO(gen[7705]),
			.S(gen[7706]),
			.SE(gen[7707]),

			.SELF(gen[7611]),
			.cell_state(gen[7611])
		); 

/******************* CELL 7612 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7612 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7516]),
			.N(gen[7517]),
			.NE(gen[7518]),

			.O(gen[7611]),
			.E(gen[7613]),

			.SO(gen[7706]),
			.S(gen[7707]),
			.SE(gen[7708]),

			.SELF(gen[7612]),
			.cell_state(gen[7612])
		); 

/******************* CELL 7613 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7613 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7517]),
			.N(gen[7518]),
			.NE(gen[7519]),

			.O(gen[7612]),
			.E(gen[7614]),

			.SO(gen[7707]),
			.S(gen[7708]),
			.SE(gen[7709]),

			.SELF(gen[7613]),
			.cell_state(gen[7613])
		); 

/******************* CELL 7614 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7614 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7518]),
			.N(gen[7519]),
			.NE(gen[7520]),

			.O(gen[7613]),
			.E(gen[7615]),

			.SO(gen[7708]),
			.S(gen[7709]),
			.SE(gen[7710]),

			.SELF(gen[7614]),
			.cell_state(gen[7614])
		); 

/******************* CELL 7615 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7615 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7519]),
			.N(gen[7520]),
			.NE(gen[7521]),

			.O(gen[7614]),
			.E(gen[7616]),

			.SO(gen[7709]),
			.S(gen[7710]),
			.SE(gen[7711]),

			.SELF(gen[7615]),
			.cell_state(gen[7615])
		); 

/******************* CELL 7616 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7616 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7520]),
			.N(gen[7521]),
			.NE(gen[7522]),

			.O(gen[7615]),
			.E(gen[7617]),

			.SO(gen[7710]),
			.S(gen[7711]),
			.SE(gen[7712]),

			.SELF(gen[7616]),
			.cell_state(gen[7616])
		); 

/******************* CELL 7617 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7617 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7521]),
			.N(gen[7522]),
			.NE(gen[7523]),

			.O(gen[7616]),
			.E(gen[7618]),

			.SO(gen[7711]),
			.S(gen[7712]),
			.SE(gen[7713]),

			.SELF(gen[7617]),
			.cell_state(gen[7617])
		); 

/******************* CELL 7618 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7618 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7522]),
			.N(gen[7523]),
			.NE(gen[7524]),

			.O(gen[7617]),
			.E(gen[7619]),

			.SO(gen[7712]),
			.S(gen[7713]),
			.SE(gen[7714]),

			.SELF(gen[7618]),
			.cell_state(gen[7618])
		); 

/******************* CELL 7619 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7619 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7523]),
			.N(gen[7524]),
			.NE(gen[7525]),

			.O(gen[7618]),
			.E(gen[7620]),

			.SO(gen[7713]),
			.S(gen[7714]),
			.SE(gen[7715]),

			.SELF(gen[7619]),
			.cell_state(gen[7619])
		); 

/******************* CELL 7620 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7620 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7524]),
			.N(gen[7525]),
			.NE(gen[7526]),

			.O(gen[7619]),
			.E(gen[7621]),

			.SO(gen[7714]),
			.S(gen[7715]),
			.SE(gen[7716]),

			.SELF(gen[7620]),
			.cell_state(gen[7620])
		); 

/******************* CELL 7621 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7621 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7525]),
			.N(gen[7526]),
			.NE(gen[7527]),

			.O(gen[7620]),
			.E(gen[7622]),

			.SO(gen[7715]),
			.S(gen[7716]),
			.SE(gen[7717]),

			.SELF(gen[7621]),
			.cell_state(gen[7621])
		); 

/******************* CELL 7622 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7622 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7526]),
			.N(gen[7527]),
			.NE(gen[7528]),

			.O(gen[7621]),
			.E(gen[7623]),

			.SO(gen[7716]),
			.S(gen[7717]),
			.SE(gen[7718]),

			.SELF(gen[7622]),
			.cell_state(gen[7622])
		); 

/******************* CELL 7623 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7623 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7527]),
			.N(gen[7528]),
			.NE(gen[7529]),

			.O(gen[7622]),
			.E(gen[7624]),

			.SO(gen[7717]),
			.S(gen[7718]),
			.SE(gen[7719]),

			.SELF(gen[7623]),
			.cell_state(gen[7623])
		); 

/******************* CELL 7624 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7624 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7528]),
			.N(gen[7529]),
			.NE(gen[7530]),

			.O(gen[7623]),
			.E(gen[7625]),

			.SO(gen[7718]),
			.S(gen[7719]),
			.SE(gen[7720]),

			.SELF(gen[7624]),
			.cell_state(gen[7624])
		); 

/******************* CELL 7625 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7625 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7529]),
			.N(gen[7530]),
			.NE(gen[7531]),

			.O(gen[7624]),
			.E(gen[7626]),

			.SO(gen[7719]),
			.S(gen[7720]),
			.SE(gen[7721]),

			.SELF(gen[7625]),
			.cell_state(gen[7625])
		); 

/******************* CELL 7626 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7626 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7530]),
			.N(gen[7531]),
			.NE(gen[7532]),

			.O(gen[7625]),
			.E(gen[7627]),

			.SO(gen[7720]),
			.S(gen[7721]),
			.SE(gen[7722]),

			.SELF(gen[7626]),
			.cell_state(gen[7626])
		); 

/******************* CELL 7627 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7627 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7531]),
			.N(gen[7532]),
			.NE(gen[7533]),

			.O(gen[7626]),
			.E(gen[7628]),

			.SO(gen[7721]),
			.S(gen[7722]),
			.SE(gen[7723]),

			.SELF(gen[7627]),
			.cell_state(gen[7627])
		); 

/******************* CELL 7628 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7628 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7532]),
			.N(gen[7533]),
			.NE(gen[7534]),

			.O(gen[7627]),
			.E(gen[7629]),

			.SO(gen[7722]),
			.S(gen[7723]),
			.SE(gen[7724]),

			.SELF(gen[7628]),
			.cell_state(gen[7628])
		); 

/******************* CELL 7629 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7629 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7533]),
			.N(gen[7534]),
			.NE(gen[7535]),

			.O(gen[7628]),
			.E(gen[7630]),

			.SO(gen[7723]),
			.S(gen[7724]),
			.SE(gen[7725]),

			.SELF(gen[7629]),
			.cell_state(gen[7629])
		); 

/******************* CELL 7630 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7630 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7534]),
			.N(gen[7535]),
			.NE(gen[7536]),

			.O(gen[7629]),
			.E(gen[7631]),

			.SO(gen[7724]),
			.S(gen[7725]),
			.SE(gen[7726]),

			.SELF(gen[7630]),
			.cell_state(gen[7630])
		); 

/******************* CELL 7631 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7631 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7535]),
			.N(gen[7536]),
			.NE(gen[7537]),

			.O(gen[7630]),
			.E(gen[7632]),

			.SO(gen[7725]),
			.S(gen[7726]),
			.SE(gen[7727]),

			.SELF(gen[7631]),
			.cell_state(gen[7631])
		); 

/******************* CELL 7632 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7632 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7536]),
			.N(gen[7537]),
			.NE(gen[7538]),

			.O(gen[7631]),
			.E(gen[7633]),

			.SO(gen[7726]),
			.S(gen[7727]),
			.SE(gen[7728]),

			.SELF(gen[7632]),
			.cell_state(gen[7632])
		); 

/******************* CELL 7633 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7633 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7537]),
			.N(gen[7538]),
			.NE(gen[7539]),

			.O(gen[7632]),
			.E(gen[7634]),

			.SO(gen[7727]),
			.S(gen[7728]),
			.SE(gen[7729]),

			.SELF(gen[7633]),
			.cell_state(gen[7633])
		); 

/******************* CELL 7634 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7634 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7538]),
			.N(gen[7539]),
			.NE(gen[7540]),

			.O(gen[7633]),
			.E(gen[7635]),

			.SO(gen[7728]),
			.S(gen[7729]),
			.SE(gen[7730]),

			.SELF(gen[7634]),
			.cell_state(gen[7634])
		); 

/******************* CELL 7635 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7635 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7539]),
			.N(gen[7540]),
			.NE(gen[7541]),

			.O(gen[7634]),
			.E(gen[7636]),

			.SO(gen[7729]),
			.S(gen[7730]),
			.SE(gen[7731]),

			.SELF(gen[7635]),
			.cell_state(gen[7635])
		); 

/******************* CELL 7636 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7636 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7540]),
			.N(gen[7541]),
			.NE(gen[7542]),

			.O(gen[7635]),
			.E(gen[7637]),

			.SO(gen[7730]),
			.S(gen[7731]),
			.SE(gen[7732]),

			.SELF(gen[7636]),
			.cell_state(gen[7636])
		); 

/******************* CELL 7637 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7637 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7541]),
			.N(gen[7542]),
			.NE(gen[7543]),

			.O(gen[7636]),
			.E(gen[7638]),

			.SO(gen[7731]),
			.S(gen[7732]),
			.SE(gen[7733]),

			.SELF(gen[7637]),
			.cell_state(gen[7637])
		); 

/******************* CELL 7638 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7638 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7542]),
			.N(gen[7543]),
			.NE(gen[7544]),

			.O(gen[7637]),
			.E(gen[7639]),

			.SO(gen[7732]),
			.S(gen[7733]),
			.SE(gen[7734]),

			.SELF(gen[7638]),
			.cell_state(gen[7638])
		); 

/******************* CELL 7639 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7639 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7543]),
			.N(gen[7544]),
			.NE(gen[7545]),

			.O(gen[7638]),
			.E(gen[7640]),

			.SO(gen[7733]),
			.S(gen[7734]),
			.SE(gen[7735]),

			.SELF(gen[7639]),
			.cell_state(gen[7639])
		); 

/******************* CELL 7640 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7640 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7544]),
			.N(gen[7545]),
			.NE(gen[7546]),

			.O(gen[7639]),
			.E(gen[7641]),

			.SO(gen[7734]),
			.S(gen[7735]),
			.SE(gen[7736]),

			.SELF(gen[7640]),
			.cell_state(gen[7640])
		); 

/******************* CELL 7641 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7641 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7545]),
			.N(gen[7546]),
			.NE(gen[7547]),

			.O(gen[7640]),
			.E(gen[7642]),

			.SO(gen[7735]),
			.S(gen[7736]),
			.SE(gen[7737]),

			.SELF(gen[7641]),
			.cell_state(gen[7641])
		); 

/******************* CELL 7642 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7642 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7546]),
			.N(gen[7547]),
			.NE(gen[7548]),

			.O(gen[7641]),
			.E(gen[7643]),

			.SO(gen[7736]),
			.S(gen[7737]),
			.SE(gen[7738]),

			.SELF(gen[7642]),
			.cell_state(gen[7642])
		); 

/******************* CELL 7643 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7643 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7547]),
			.N(gen[7548]),
			.NE(gen[7549]),

			.O(gen[7642]),
			.E(gen[7644]),

			.SO(gen[7737]),
			.S(gen[7738]),
			.SE(gen[7739]),

			.SELF(gen[7643]),
			.cell_state(gen[7643])
		); 

/******************* CELL 7644 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7644 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7548]),
			.N(gen[7549]),
			.NE(gen[7550]),

			.O(gen[7643]),
			.E(gen[7645]),

			.SO(gen[7738]),
			.S(gen[7739]),
			.SE(gen[7740]),

			.SELF(gen[7644]),
			.cell_state(gen[7644])
		); 

/******************* CELL 7645 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7645 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7549]),
			.N(gen[7550]),
			.NE(gen[7551]),

			.O(gen[7644]),
			.E(gen[7646]),

			.SO(gen[7739]),
			.S(gen[7740]),
			.SE(gen[7741]),

			.SELF(gen[7645]),
			.cell_state(gen[7645])
		); 

/******************* CELL 7646 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7646 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7550]),
			.N(gen[7551]),
			.NE(gen[7552]),

			.O(gen[7645]),
			.E(gen[7647]),

			.SO(gen[7740]),
			.S(gen[7741]),
			.SE(gen[7742]),

			.SELF(gen[7646]),
			.cell_state(gen[7646])
		); 

/******************* CELL 7647 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7647 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7551]),
			.N(gen[7552]),
			.NE(gen[7553]),

			.O(gen[7646]),
			.E(gen[7648]),

			.SO(gen[7741]),
			.S(gen[7742]),
			.SE(gen[7743]),

			.SELF(gen[7647]),
			.cell_state(gen[7647])
		); 

/******************* CELL 7648 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7648 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7552]),
			.N(gen[7553]),
			.NE(gen[7554]),

			.O(gen[7647]),
			.E(gen[7649]),

			.SO(gen[7742]),
			.S(gen[7743]),
			.SE(gen[7744]),

			.SELF(gen[7648]),
			.cell_state(gen[7648])
		); 

/******************* CELL 7649 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7649 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7553]),
			.N(gen[7554]),
			.NE(gen[7555]),

			.O(gen[7648]),
			.E(gen[7650]),

			.SO(gen[7743]),
			.S(gen[7744]),
			.SE(gen[7745]),

			.SELF(gen[7649]),
			.cell_state(gen[7649])
		); 

/******************* CELL 7650 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7650 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7554]),
			.N(gen[7555]),
			.NE(gen[7556]),

			.O(gen[7649]),
			.E(gen[7651]),

			.SO(gen[7744]),
			.S(gen[7745]),
			.SE(gen[7746]),

			.SELF(gen[7650]),
			.cell_state(gen[7650])
		); 

/******************* CELL 7651 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7651 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7555]),
			.N(gen[7556]),
			.NE(gen[7557]),

			.O(gen[7650]),
			.E(gen[7652]),

			.SO(gen[7745]),
			.S(gen[7746]),
			.SE(gen[7747]),

			.SELF(gen[7651]),
			.cell_state(gen[7651])
		); 

/******************* CELL 7652 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7652 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7556]),
			.N(gen[7557]),
			.NE(gen[7558]),

			.O(gen[7651]),
			.E(gen[7653]),

			.SO(gen[7746]),
			.S(gen[7747]),
			.SE(gen[7748]),

			.SELF(gen[7652]),
			.cell_state(gen[7652])
		); 

/******************* CELL 7653 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7653 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7557]),
			.N(gen[7558]),
			.NE(gen[7559]),

			.O(gen[7652]),
			.E(gen[7654]),

			.SO(gen[7747]),
			.S(gen[7748]),
			.SE(gen[7749]),

			.SELF(gen[7653]),
			.cell_state(gen[7653])
		); 

/******************* CELL 7654 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7654 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7558]),
			.N(gen[7559]),
			.NE(gen[7560]),

			.O(gen[7653]),
			.E(gen[7655]),

			.SO(gen[7748]),
			.S(gen[7749]),
			.SE(gen[7750]),

			.SELF(gen[7654]),
			.cell_state(gen[7654])
		); 

/******************* CELL 7655 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7655 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7559]),
			.N(gen[7560]),
			.NE(gen[7561]),

			.O(gen[7654]),
			.E(gen[7656]),

			.SO(gen[7749]),
			.S(gen[7750]),
			.SE(gen[7751]),

			.SELF(gen[7655]),
			.cell_state(gen[7655])
		); 

/******************* CELL 7656 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7656 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7560]),
			.N(gen[7561]),
			.NE(gen[7562]),

			.O(gen[7655]),
			.E(gen[7657]),

			.SO(gen[7750]),
			.S(gen[7751]),
			.SE(gen[7752]),

			.SELF(gen[7656]),
			.cell_state(gen[7656])
		); 

/******************* CELL 7657 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7657 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7561]),
			.N(gen[7562]),
			.NE(gen[7563]),

			.O(gen[7656]),
			.E(gen[7658]),

			.SO(gen[7751]),
			.S(gen[7752]),
			.SE(gen[7753]),

			.SELF(gen[7657]),
			.cell_state(gen[7657])
		); 

/******************* CELL 7658 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7658 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7562]),
			.N(gen[7563]),
			.NE(gen[7564]),

			.O(gen[7657]),
			.E(gen[7659]),

			.SO(gen[7752]),
			.S(gen[7753]),
			.SE(gen[7754]),

			.SELF(gen[7658]),
			.cell_state(gen[7658])
		); 

/******************* CELL 7659 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7659 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7563]),
			.N(gen[7564]),
			.NE(gen[7565]),

			.O(gen[7658]),
			.E(gen[7660]),

			.SO(gen[7753]),
			.S(gen[7754]),
			.SE(gen[7755]),

			.SELF(gen[7659]),
			.cell_state(gen[7659])
		); 

/******************* CELL 7660 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7660 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7564]),
			.N(gen[7565]),
			.NE(gen[7566]),

			.O(gen[7659]),
			.E(gen[7661]),

			.SO(gen[7754]),
			.S(gen[7755]),
			.SE(gen[7756]),

			.SELF(gen[7660]),
			.cell_state(gen[7660])
		); 

/******************* CELL 7661 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7661 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7565]),
			.N(gen[7566]),
			.NE(gen[7567]),

			.O(gen[7660]),
			.E(gen[7662]),

			.SO(gen[7755]),
			.S(gen[7756]),
			.SE(gen[7757]),

			.SELF(gen[7661]),
			.cell_state(gen[7661])
		); 

/******************* CELL 7662 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7662 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7566]),
			.N(gen[7567]),
			.NE(gen[7568]),

			.O(gen[7661]),
			.E(gen[7663]),

			.SO(gen[7756]),
			.S(gen[7757]),
			.SE(gen[7758]),

			.SELF(gen[7662]),
			.cell_state(gen[7662])
		); 

/******************* CELL 7663 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7663 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7567]),
			.N(gen[7568]),
			.NE(gen[7569]),

			.O(gen[7662]),
			.E(gen[7664]),

			.SO(gen[7757]),
			.S(gen[7758]),
			.SE(gen[7759]),

			.SELF(gen[7663]),
			.cell_state(gen[7663])
		); 

/******************* CELL 7664 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7664 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7568]),
			.N(gen[7569]),
			.NE(gen[7570]),

			.O(gen[7663]),
			.E(gen[7665]),

			.SO(gen[7758]),
			.S(gen[7759]),
			.SE(gen[7760]),

			.SELF(gen[7664]),
			.cell_state(gen[7664])
		); 

/******************* CELL 7665 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7665 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7569]),
			.N(gen[7570]),
			.NE(gen[7571]),

			.O(gen[7664]),
			.E(gen[7666]),

			.SO(gen[7759]),
			.S(gen[7760]),
			.SE(gen[7761]),

			.SELF(gen[7665]),
			.cell_state(gen[7665])
		); 

/******************* CELL 7666 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7666 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7570]),
			.N(gen[7571]),
			.NE(gen[7572]),

			.O(gen[7665]),
			.E(gen[7667]),

			.SO(gen[7760]),
			.S(gen[7761]),
			.SE(gen[7762]),

			.SELF(gen[7666]),
			.cell_state(gen[7666])
		); 

/******************* CELL 7667 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7667 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7571]),
			.N(gen[7572]),
			.NE(gen[7573]),

			.O(gen[7666]),
			.E(gen[7668]),

			.SO(gen[7761]),
			.S(gen[7762]),
			.SE(gen[7763]),

			.SELF(gen[7667]),
			.cell_state(gen[7667])
		); 

/******************* CELL 7668 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7668 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7572]),
			.N(gen[7573]),
			.NE(gen[7574]),

			.O(gen[7667]),
			.E(gen[7669]),

			.SO(gen[7762]),
			.S(gen[7763]),
			.SE(gen[7764]),

			.SELF(gen[7668]),
			.cell_state(gen[7668])
		); 

/******************* CELL 7669 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7669 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7573]),
			.N(gen[7574]),
			.NE(gen[7575]),

			.O(gen[7668]),
			.E(gen[7670]),

			.SO(gen[7763]),
			.S(gen[7764]),
			.SE(gen[7765]),

			.SELF(gen[7669]),
			.cell_state(gen[7669])
		); 

/******************* CELL 7670 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7670 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7574]),
			.N(gen[7575]),
			.NE(gen[7576]),

			.O(gen[7669]),
			.E(gen[7671]),

			.SO(gen[7764]),
			.S(gen[7765]),
			.SE(gen[7766]),

			.SELF(gen[7670]),
			.cell_state(gen[7670])
		); 

/******************* CELL 7671 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7671 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7575]),
			.N(gen[7576]),
			.NE(gen[7577]),

			.O(gen[7670]),
			.E(gen[7672]),

			.SO(gen[7765]),
			.S(gen[7766]),
			.SE(gen[7767]),

			.SELF(gen[7671]),
			.cell_state(gen[7671])
		); 

/******************* CELL 7672 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7672 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7576]),
			.N(gen[7577]),
			.NE(gen[7578]),

			.O(gen[7671]),
			.E(gen[7673]),

			.SO(gen[7766]),
			.S(gen[7767]),
			.SE(gen[7768]),

			.SELF(gen[7672]),
			.cell_state(gen[7672])
		); 

/******************* CELL 7673 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7673 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7577]),
			.N(gen[7578]),
			.NE(gen[7579]),

			.O(gen[7672]),
			.E(gen[7674]),

			.SO(gen[7767]),
			.S(gen[7768]),
			.SE(gen[7769]),

			.SELF(gen[7673]),
			.cell_state(gen[7673])
		); 

/******************* CELL 7674 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7674 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7578]),
			.N(gen[7579]),
			.NE(gen[7580]),

			.O(gen[7673]),
			.E(gen[7675]),

			.SO(gen[7768]),
			.S(gen[7769]),
			.SE(gen[7770]),

			.SELF(gen[7674]),
			.cell_state(gen[7674])
		); 

/******************* CELL 7675 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7675 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7579]),
			.N(gen[7580]),
			.NE(gen[7581]),

			.O(gen[7674]),
			.E(gen[7676]),

			.SO(gen[7769]),
			.S(gen[7770]),
			.SE(gen[7771]),

			.SELF(gen[7675]),
			.cell_state(gen[7675])
		); 

/******************* CELL 7676 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7676 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7580]),
			.N(gen[7581]),
			.NE(gen[7582]),

			.O(gen[7675]),
			.E(gen[7677]),

			.SO(gen[7770]),
			.S(gen[7771]),
			.SE(gen[7772]),

			.SELF(gen[7676]),
			.cell_state(gen[7676])
		); 

/******************* CELL 7677 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7677 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7581]),
			.N(gen[7582]),
			.NE(gen[7583]),

			.O(gen[7676]),
			.E(gen[7678]),

			.SO(gen[7771]),
			.S(gen[7772]),
			.SE(gen[7773]),

			.SELF(gen[7677]),
			.cell_state(gen[7677])
		); 

/******************* CELL 7678 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7678 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7582]),
			.N(gen[7583]),
			.NE(gen[7584]),

			.O(gen[7677]),
			.E(gen[7679]),

			.SO(gen[7772]),
			.S(gen[7773]),
			.SE(gen[7774]),

			.SELF(gen[7678]),
			.cell_state(gen[7678])
		); 

/******************* CELL 7679 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7679 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7583]),
			.N(gen[7584]),
			.NE(gen[7585]),

			.O(gen[7678]),
			.E(gen[7680]),

			.SO(gen[7773]),
			.S(gen[7774]),
			.SE(gen[7775]),

			.SELF(gen[7679]),
			.cell_state(gen[7679])
		); 

/******************* CELL 7680 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7680 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7584]),
			.N(gen[7585]),
			.NE(gen[7586]),

			.O(gen[7679]),
			.E(gen[7681]),

			.SO(gen[7774]),
			.S(gen[7775]),
			.SE(gen[7776]),

			.SELF(gen[7680]),
			.cell_state(gen[7680])
		); 

/******************* CELL 7681 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7681 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7585]),
			.N(gen[7586]),
			.NE(gen[7587]),

			.O(gen[7680]),
			.E(gen[7682]),

			.SO(gen[7775]),
			.S(gen[7776]),
			.SE(gen[7777]),

			.SELF(gen[7681]),
			.cell_state(gen[7681])
		); 

/******************* CELL 7682 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7682 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7586]),
			.N(gen[7587]),
			.NE(gen[7588]),

			.O(gen[7681]),
			.E(gen[7683]),

			.SO(gen[7776]),
			.S(gen[7777]),
			.SE(gen[7778]),

			.SELF(gen[7682]),
			.cell_state(gen[7682])
		); 

/******************* CELL 7683 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7683 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7587]),
			.N(gen[7588]),
			.NE(gen[7589]),

			.O(gen[7682]),
			.E(gen[7684]),

			.SO(gen[7777]),
			.S(gen[7778]),
			.SE(gen[7779]),

			.SELF(gen[7683]),
			.cell_state(gen[7683])
		); 

/******************* CELL 7684 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7684 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7588]),
			.N(gen[7589]),
			.NE(gen[7590]),

			.O(gen[7683]),
			.E(gen[7685]),

			.SO(gen[7778]),
			.S(gen[7779]),
			.SE(gen[7780]),

			.SELF(gen[7684]),
			.cell_state(gen[7684])
		); 

/******************* CELL 7685 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7685 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7589]),
			.N(gen[7590]),
			.NE(gen[7591]),

			.O(gen[7684]),
			.E(gen[7686]),

			.SO(gen[7779]),
			.S(gen[7780]),
			.SE(gen[7781]),

			.SELF(gen[7685]),
			.cell_state(gen[7685])
		); 

/******************* CELL 7686 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7686 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7590]),
			.N(gen[7591]),
			.NE(gen[7592]),

			.O(gen[7685]),
			.E(gen[7687]),

			.SO(gen[7780]),
			.S(gen[7781]),
			.SE(gen[7782]),

			.SELF(gen[7686]),
			.cell_state(gen[7686])
		); 

/******************* CELL 7687 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7687 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7591]),
			.N(gen[7592]),
			.NE(gen[7593]),

			.O(gen[7686]),
			.E(gen[7688]),

			.SO(gen[7781]),
			.S(gen[7782]),
			.SE(gen[7783]),

			.SELF(gen[7687]),
			.cell_state(gen[7687])
		); 

/******************* CELL 7688 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7688 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7592]),
			.N(gen[7593]),
			.NE(gen[7594]),

			.O(gen[7687]),
			.E(gen[7689]),

			.SO(gen[7782]),
			.S(gen[7783]),
			.SE(gen[7784]),

			.SELF(gen[7688]),
			.cell_state(gen[7688])
		); 

/******************* CELL 7689 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7689 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7593]),
			.N(gen[7594]),
			.NE(gen[7595]),

			.O(gen[7688]),
			.E(gen[7690]),

			.SO(gen[7783]),
			.S(gen[7784]),
			.SE(gen[7785]),

			.SELF(gen[7689]),
			.cell_state(gen[7689])
		); 

/******************* CELL 7690 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7690 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7594]),
			.N(gen[7595]),
			.NE(gen[7596]),

			.O(gen[7689]),
			.E(gen[7691]),

			.SO(gen[7784]),
			.S(gen[7785]),
			.SE(gen[7786]),

			.SELF(gen[7690]),
			.cell_state(gen[7690])
		); 

/******************* CELL 7691 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7691 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7595]),
			.N(gen[7596]),
			.NE(gen[7597]),

			.O(gen[7690]),
			.E(gen[7692]),

			.SO(gen[7785]),
			.S(gen[7786]),
			.SE(gen[7787]),

			.SELF(gen[7691]),
			.cell_state(gen[7691])
		); 

/******************* CELL 7692 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7692 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7596]),
			.N(gen[7597]),
			.NE(gen[7598]),

			.O(gen[7691]),
			.E(gen[7693]),

			.SO(gen[7786]),
			.S(gen[7787]),
			.SE(gen[7788]),

			.SELF(gen[7692]),
			.cell_state(gen[7692])
		); 

/******************* CELL 7693 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7693 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7597]),
			.N(gen[7598]),
			.NE(gen[7599]),

			.O(gen[7692]),
			.E(gen[7694]),

			.SO(gen[7787]),
			.S(gen[7788]),
			.SE(gen[7789]),

			.SELF(gen[7693]),
			.cell_state(gen[7693])
		); 

/******************* CELL 7694 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7694 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7598]),
			.N(gen[7599]),
			.NE(gen[7598]),

			.O(gen[7693]),
			.E(gen[7693]),

			.SO(gen[7788]),
			.S(gen[7789]),
			.SE(gen[7788]),

			.SELF(gen[7694]),
			.cell_state(gen[7694])
		); 

/******************* CELL 7695 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7695 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7601]),
			.N(gen[7600]),
			.NE(gen[7601]),

			.O(gen[7696]),
			.E(gen[7696]),

			.SO(gen[7791]),
			.S(gen[7790]),
			.SE(gen[7791]),

			.SELF(gen[7695]),
			.cell_state(gen[7695])
		); 

/******************* CELL 7696 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7696 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7600]),
			.N(gen[7601]),
			.NE(gen[7602]),

			.O(gen[7695]),
			.E(gen[7697]),

			.SO(gen[7790]),
			.S(gen[7791]),
			.SE(gen[7792]),

			.SELF(gen[7696]),
			.cell_state(gen[7696])
		); 

/******************* CELL 7697 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7697 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7601]),
			.N(gen[7602]),
			.NE(gen[7603]),

			.O(gen[7696]),
			.E(gen[7698]),

			.SO(gen[7791]),
			.S(gen[7792]),
			.SE(gen[7793]),

			.SELF(gen[7697]),
			.cell_state(gen[7697])
		); 

/******************* CELL 7698 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7698 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7602]),
			.N(gen[7603]),
			.NE(gen[7604]),

			.O(gen[7697]),
			.E(gen[7699]),

			.SO(gen[7792]),
			.S(gen[7793]),
			.SE(gen[7794]),

			.SELF(gen[7698]),
			.cell_state(gen[7698])
		); 

/******************* CELL 7699 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7699 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7603]),
			.N(gen[7604]),
			.NE(gen[7605]),

			.O(gen[7698]),
			.E(gen[7700]),

			.SO(gen[7793]),
			.S(gen[7794]),
			.SE(gen[7795]),

			.SELF(gen[7699]),
			.cell_state(gen[7699])
		); 

/******************* CELL 7700 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7700 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7604]),
			.N(gen[7605]),
			.NE(gen[7606]),

			.O(gen[7699]),
			.E(gen[7701]),

			.SO(gen[7794]),
			.S(gen[7795]),
			.SE(gen[7796]),

			.SELF(gen[7700]),
			.cell_state(gen[7700])
		); 

/******************* CELL 7701 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7701 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7605]),
			.N(gen[7606]),
			.NE(gen[7607]),

			.O(gen[7700]),
			.E(gen[7702]),

			.SO(gen[7795]),
			.S(gen[7796]),
			.SE(gen[7797]),

			.SELF(gen[7701]),
			.cell_state(gen[7701])
		); 

/******************* CELL 7702 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7702 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7606]),
			.N(gen[7607]),
			.NE(gen[7608]),

			.O(gen[7701]),
			.E(gen[7703]),

			.SO(gen[7796]),
			.S(gen[7797]),
			.SE(gen[7798]),

			.SELF(gen[7702]),
			.cell_state(gen[7702])
		); 

/******************* CELL 7703 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7703 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7607]),
			.N(gen[7608]),
			.NE(gen[7609]),

			.O(gen[7702]),
			.E(gen[7704]),

			.SO(gen[7797]),
			.S(gen[7798]),
			.SE(gen[7799]),

			.SELF(gen[7703]),
			.cell_state(gen[7703])
		); 

/******************* CELL 7704 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7704 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7608]),
			.N(gen[7609]),
			.NE(gen[7610]),

			.O(gen[7703]),
			.E(gen[7705]),

			.SO(gen[7798]),
			.S(gen[7799]),
			.SE(gen[7800]),

			.SELF(gen[7704]),
			.cell_state(gen[7704])
		); 

/******************* CELL 7705 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7705 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7609]),
			.N(gen[7610]),
			.NE(gen[7611]),

			.O(gen[7704]),
			.E(gen[7706]),

			.SO(gen[7799]),
			.S(gen[7800]),
			.SE(gen[7801]),

			.SELF(gen[7705]),
			.cell_state(gen[7705])
		); 

/******************* CELL 7706 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7706 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7610]),
			.N(gen[7611]),
			.NE(gen[7612]),

			.O(gen[7705]),
			.E(gen[7707]),

			.SO(gen[7800]),
			.S(gen[7801]),
			.SE(gen[7802]),

			.SELF(gen[7706]),
			.cell_state(gen[7706])
		); 

/******************* CELL 7707 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7707 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7611]),
			.N(gen[7612]),
			.NE(gen[7613]),

			.O(gen[7706]),
			.E(gen[7708]),

			.SO(gen[7801]),
			.S(gen[7802]),
			.SE(gen[7803]),

			.SELF(gen[7707]),
			.cell_state(gen[7707])
		); 

/******************* CELL 7708 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7708 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7612]),
			.N(gen[7613]),
			.NE(gen[7614]),

			.O(gen[7707]),
			.E(gen[7709]),

			.SO(gen[7802]),
			.S(gen[7803]),
			.SE(gen[7804]),

			.SELF(gen[7708]),
			.cell_state(gen[7708])
		); 

/******************* CELL 7709 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7709 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7613]),
			.N(gen[7614]),
			.NE(gen[7615]),

			.O(gen[7708]),
			.E(gen[7710]),

			.SO(gen[7803]),
			.S(gen[7804]),
			.SE(gen[7805]),

			.SELF(gen[7709]),
			.cell_state(gen[7709])
		); 

/******************* CELL 7710 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7710 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7614]),
			.N(gen[7615]),
			.NE(gen[7616]),

			.O(gen[7709]),
			.E(gen[7711]),

			.SO(gen[7804]),
			.S(gen[7805]),
			.SE(gen[7806]),

			.SELF(gen[7710]),
			.cell_state(gen[7710])
		); 

/******************* CELL 7711 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7711 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7615]),
			.N(gen[7616]),
			.NE(gen[7617]),

			.O(gen[7710]),
			.E(gen[7712]),

			.SO(gen[7805]),
			.S(gen[7806]),
			.SE(gen[7807]),

			.SELF(gen[7711]),
			.cell_state(gen[7711])
		); 

/******************* CELL 7712 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7712 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7616]),
			.N(gen[7617]),
			.NE(gen[7618]),

			.O(gen[7711]),
			.E(gen[7713]),

			.SO(gen[7806]),
			.S(gen[7807]),
			.SE(gen[7808]),

			.SELF(gen[7712]),
			.cell_state(gen[7712])
		); 

/******************* CELL 7713 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7713 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7617]),
			.N(gen[7618]),
			.NE(gen[7619]),

			.O(gen[7712]),
			.E(gen[7714]),

			.SO(gen[7807]),
			.S(gen[7808]),
			.SE(gen[7809]),

			.SELF(gen[7713]),
			.cell_state(gen[7713])
		); 

/******************* CELL 7714 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7714 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7618]),
			.N(gen[7619]),
			.NE(gen[7620]),

			.O(gen[7713]),
			.E(gen[7715]),

			.SO(gen[7808]),
			.S(gen[7809]),
			.SE(gen[7810]),

			.SELF(gen[7714]),
			.cell_state(gen[7714])
		); 

/******************* CELL 7715 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7715 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7619]),
			.N(gen[7620]),
			.NE(gen[7621]),

			.O(gen[7714]),
			.E(gen[7716]),

			.SO(gen[7809]),
			.S(gen[7810]),
			.SE(gen[7811]),

			.SELF(gen[7715]),
			.cell_state(gen[7715])
		); 

/******************* CELL 7716 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7716 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7620]),
			.N(gen[7621]),
			.NE(gen[7622]),

			.O(gen[7715]),
			.E(gen[7717]),

			.SO(gen[7810]),
			.S(gen[7811]),
			.SE(gen[7812]),

			.SELF(gen[7716]),
			.cell_state(gen[7716])
		); 

/******************* CELL 7717 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7717 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7621]),
			.N(gen[7622]),
			.NE(gen[7623]),

			.O(gen[7716]),
			.E(gen[7718]),

			.SO(gen[7811]),
			.S(gen[7812]),
			.SE(gen[7813]),

			.SELF(gen[7717]),
			.cell_state(gen[7717])
		); 

/******************* CELL 7718 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7718 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7622]),
			.N(gen[7623]),
			.NE(gen[7624]),

			.O(gen[7717]),
			.E(gen[7719]),

			.SO(gen[7812]),
			.S(gen[7813]),
			.SE(gen[7814]),

			.SELF(gen[7718]),
			.cell_state(gen[7718])
		); 

/******************* CELL 7719 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7719 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7623]),
			.N(gen[7624]),
			.NE(gen[7625]),

			.O(gen[7718]),
			.E(gen[7720]),

			.SO(gen[7813]),
			.S(gen[7814]),
			.SE(gen[7815]),

			.SELF(gen[7719]),
			.cell_state(gen[7719])
		); 

/******************* CELL 7720 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7720 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7624]),
			.N(gen[7625]),
			.NE(gen[7626]),

			.O(gen[7719]),
			.E(gen[7721]),

			.SO(gen[7814]),
			.S(gen[7815]),
			.SE(gen[7816]),

			.SELF(gen[7720]),
			.cell_state(gen[7720])
		); 

/******************* CELL 7721 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7721 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7625]),
			.N(gen[7626]),
			.NE(gen[7627]),

			.O(gen[7720]),
			.E(gen[7722]),

			.SO(gen[7815]),
			.S(gen[7816]),
			.SE(gen[7817]),

			.SELF(gen[7721]),
			.cell_state(gen[7721])
		); 

/******************* CELL 7722 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7722 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7626]),
			.N(gen[7627]),
			.NE(gen[7628]),

			.O(gen[7721]),
			.E(gen[7723]),

			.SO(gen[7816]),
			.S(gen[7817]),
			.SE(gen[7818]),

			.SELF(gen[7722]),
			.cell_state(gen[7722])
		); 

/******************* CELL 7723 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7723 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7627]),
			.N(gen[7628]),
			.NE(gen[7629]),

			.O(gen[7722]),
			.E(gen[7724]),

			.SO(gen[7817]),
			.S(gen[7818]),
			.SE(gen[7819]),

			.SELF(gen[7723]),
			.cell_state(gen[7723])
		); 

/******************* CELL 7724 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7724 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7628]),
			.N(gen[7629]),
			.NE(gen[7630]),

			.O(gen[7723]),
			.E(gen[7725]),

			.SO(gen[7818]),
			.S(gen[7819]),
			.SE(gen[7820]),

			.SELF(gen[7724]),
			.cell_state(gen[7724])
		); 

/******************* CELL 7725 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7725 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7629]),
			.N(gen[7630]),
			.NE(gen[7631]),

			.O(gen[7724]),
			.E(gen[7726]),

			.SO(gen[7819]),
			.S(gen[7820]),
			.SE(gen[7821]),

			.SELF(gen[7725]),
			.cell_state(gen[7725])
		); 

/******************* CELL 7726 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7726 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7630]),
			.N(gen[7631]),
			.NE(gen[7632]),

			.O(gen[7725]),
			.E(gen[7727]),

			.SO(gen[7820]),
			.S(gen[7821]),
			.SE(gen[7822]),

			.SELF(gen[7726]),
			.cell_state(gen[7726])
		); 

/******************* CELL 7727 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7727 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7631]),
			.N(gen[7632]),
			.NE(gen[7633]),

			.O(gen[7726]),
			.E(gen[7728]),

			.SO(gen[7821]),
			.S(gen[7822]),
			.SE(gen[7823]),

			.SELF(gen[7727]),
			.cell_state(gen[7727])
		); 

/******************* CELL 7728 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7728 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7632]),
			.N(gen[7633]),
			.NE(gen[7634]),

			.O(gen[7727]),
			.E(gen[7729]),

			.SO(gen[7822]),
			.S(gen[7823]),
			.SE(gen[7824]),

			.SELF(gen[7728]),
			.cell_state(gen[7728])
		); 

/******************* CELL 7729 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7729 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7633]),
			.N(gen[7634]),
			.NE(gen[7635]),

			.O(gen[7728]),
			.E(gen[7730]),

			.SO(gen[7823]),
			.S(gen[7824]),
			.SE(gen[7825]),

			.SELF(gen[7729]),
			.cell_state(gen[7729])
		); 

/******************* CELL 7730 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7730 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7634]),
			.N(gen[7635]),
			.NE(gen[7636]),

			.O(gen[7729]),
			.E(gen[7731]),

			.SO(gen[7824]),
			.S(gen[7825]),
			.SE(gen[7826]),

			.SELF(gen[7730]),
			.cell_state(gen[7730])
		); 

/******************* CELL 7731 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7731 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7635]),
			.N(gen[7636]),
			.NE(gen[7637]),

			.O(gen[7730]),
			.E(gen[7732]),

			.SO(gen[7825]),
			.S(gen[7826]),
			.SE(gen[7827]),

			.SELF(gen[7731]),
			.cell_state(gen[7731])
		); 

/******************* CELL 7732 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7732 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7636]),
			.N(gen[7637]),
			.NE(gen[7638]),

			.O(gen[7731]),
			.E(gen[7733]),

			.SO(gen[7826]),
			.S(gen[7827]),
			.SE(gen[7828]),

			.SELF(gen[7732]),
			.cell_state(gen[7732])
		); 

/******************* CELL 7733 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7733 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7637]),
			.N(gen[7638]),
			.NE(gen[7639]),

			.O(gen[7732]),
			.E(gen[7734]),

			.SO(gen[7827]),
			.S(gen[7828]),
			.SE(gen[7829]),

			.SELF(gen[7733]),
			.cell_state(gen[7733])
		); 

/******************* CELL 7734 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7734 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7638]),
			.N(gen[7639]),
			.NE(gen[7640]),

			.O(gen[7733]),
			.E(gen[7735]),

			.SO(gen[7828]),
			.S(gen[7829]),
			.SE(gen[7830]),

			.SELF(gen[7734]),
			.cell_state(gen[7734])
		); 

/******************* CELL 7735 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7735 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7639]),
			.N(gen[7640]),
			.NE(gen[7641]),

			.O(gen[7734]),
			.E(gen[7736]),

			.SO(gen[7829]),
			.S(gen[7830]),
			.SE(gen[7831]),

			.SELF(gen[7735]),
			.cell_state(gen[7735])
		); 

/******************* CELL 7736 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7736 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7640]),
			.N(gen[7641]),
			.NE(gen[7642]),

			.O(gen[7735]),
			.E(gen[7737]),

			.SO(gen[7830]),
			.S(gen[7831]),
			.SE(gen[7832]),

			.SELF(gen[7736]),
			.cell_state(gen[7736])
		); 

/******************* CELL 7737 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7737 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7641]),
			.N(gen[7642]),
			.NE(gen[7643]),

			.O(gen[7736]),
			.E(gen[7738]),

			.SO(gen[7831]),
			.S(gen[7832]),
			.SE(gen[7833]),

			.SELF(gen[7737]),
			.cell_state(gen[7737])
		); 

/******************* CELL 7738 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7738 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7642]),
			.N(gen[7643]),
			.NE(gen[7644]),

			.O(gen[7737]),
			.E(gen[7739]),

			.SO(gen[7832]),
			.S(gen[7833]),
			.SE(gen[7834]),

			.SELF(gen[7738]),
			.cell_state(gen[7738])
		); 

/******************* CELL 7739 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7739 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7643]),
			.N(gen[7644]),
			.NE(gen[7645]),

			.O(gen[7738]),
			.E(gen[7740]),

			.SO(gen[7833]),
			.S(gen[7834]),
			.SE(gen[7835]),

			.SELF(gen[7739]),
			.cell_state(gen[7739])
		); 

/******************* CELL 7740 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7740 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7644]),
			.N(gen[7645]),
			.NE(gen[7646]),

			.O(gen[7739]),
			.E(gen[7741]),

			.SO(gen[7834]),
			.S(gen[7835]),
			.SE(gen[7836]),

			.SELF(gen[7740]),
			.cell_state(gen[7740])
		); 

/******************* CELL 7741 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7741 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7645]),
			.N(gen[7646]),
			.NE(gen[7647]),

			.O(gen[7740]),
			.E(gen[7742]),

			.SO(gen[7835]),
			.S(gen[7836]),
			.SE(gen[7837]),

			.SELF(gen[7741]),
			.cell_state(gen[7741])
		); 

/******************* CELL 7742 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7742 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7646]),
			.N(gen[7647]),
			.NE(gen[7648]),

			.O(gen[7741]),
			.E(gen[7743]),

			.SO(gen[7836]),
			.S(gen[7837]),
			.SE(gen[7838]),

			.SELF(gen[7742]),
			.cell_state(gen[7742])
		); 

/******************* CELL 7743 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7743 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7647]),
			.N(gen[7648]),
			.NE(gen[7649]),

			.O(gen[7742]),
			.E(gen[7744]),

			.SO(gen[7837]),
			.S(gen[7838]),
			.SE(gen[7839]),

			.SELF(gen[7743]),
			.cell_state(gen[7743])
		); 

/******************* CELL 7744 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7744 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7648]),
			.N(gen[7649]),
			.NE(gen[7650]),

			.O(gen[7743]),
			.E(gen[7745]),

			.SO(gen[7838]),
			.S(gen[7839]),
			.SE(gen[7840]),

			.SELF(gen[7744]),
			.cell_state(gen[7744])
		); 

/******************* CELL 7745 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7745 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7649]),
			.N(gen[7650]),
			.NE(gen[7651]),

			.O(gen[7744]),
			.E(gen[7746]),

			.SO(gen[7839]),
			.S(gen[7840]),
			.SE(gen[7841]),

			.SELF(gen[7745]),
			.cell_state(gen[7745])
		); 

/******************* CELL 7746 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7746 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7650]),
			.N(gen[7651]),
			.NE(gen[7652]),

			.O(gen[7745]),
			.E(gen[7747]),

			.SO(gen[7840]),
			.S(gen[7841]),
			.SE(gen[7842]),

			.SELF(gen[7746]),
			.cell_state(gen[7746])
		); 

/******************* CELL 7747 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7747 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7651]),
			.N(gen[7652]),
			.NE(gen[7653]),

			.O(gen[7746]),
			.E(gen[7748]),

			.SO(gen[7841]),
			.S(gen[7842]),
			.SE(gen[7843]),

			.SELF(gen[7747]),
			.cell_state(gen[7747])
		); 

/******************* CELL 7748 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7748 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7652]),
			.N(gen[7653]),
			.NE(gen[7654]),

			.O(gen[7747]),
			.E(gen[7749]),

			.SO(gen[7842]),
			.S(gen[7843]),
			.SE(gen[7844]),

			.SELF(gen[7748]),
			.cell_state(gen[7748])
		); 

/******************* CELL 7749 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7749 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7653]),
			.N(gen[7654]),
			.NE(gen[7655]),

			.O(gen[7748]),
			.E(gen[7750]),

			.SO(gen[7843]),
			.S(gen[7844]),
			.SE(gen[7845]),

			.SELF(gen[7749]),
			.cell_state(gen[7749])
		); 

/******************* CELL 7750 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7750 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7654]),
			.N(gen[7655]),
			.NE(gen[7656]),

			.O(gen[7749]),
			.E(gen[7751]),

			.SO(gen[7844]),
			.S(gen[7845]),
			.SE(gen[7846]),

			.SELF(gen[7750]),
			.cell_state(gen[7750])
		); 

/******************* CELL 7751 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7751 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7655]),
			.N(gen[7656]),
			.NE(gen[7657]),

			.O(gen[7750]),
			.E(gen[7752]),

			.SO(gen[7845]),
			.S(gen[7846]),
			.SE(gen[7847]),

			.SELF(gen[7751]),
			.cell_state(gen[7751])
		); 

/******************* CELL 7752 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7752 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7656]),
			.N(gen[7657]),
			.NE(gen[7658]),

			.O(gen[7751]),
			.E(gen[7753]),

			.SO(gen[7846]),
			.S(gen[7847]),
			.SE(gen[7848]),

			.SELF(gen[7752]),
			.cell_state(gen[7752])
		); 

/******************* CELL 7753 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7753 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7657]),
			.N(gen[7658]),
			.NE(gen[7659]),

			.O(gen[7752]),
			.E(gen[7754]),

			.SO(gen[7847]),
			.S(gen[7848]),
			.SE(gen[7849]),

			.SELF(gen[7753]),
			.cell_state(gen[7753])
		); 

/******************* CELL 7754 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7754 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7658]),
			.N(gen[7659]),
			.NE(gen[7660]),

			.O(gen[7753]),
			.E(gen[7755]),

			.SO(gen[7848]),
			.S(gen[7849]),
			.SE(gen[7850]),

			.SELF(gen[7754]),
			.cell_state(gen[7754])
		); 

/******************* CELL 7755 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7755 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7659]),
			.N(gen[7660]),
			.NE(gen[7661]),

			.O(gen[7754]),
			.E(gen[7756]),

			.SO(gen[7849]),
			.S(gen[7850]),
			.SE(gen[7851]),

			.SELF(gen[7755]),
			.cell_state(gen[7755])
		); 

/******************* CELL 7756 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7756 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7660]),
			.N(gen[7661]),
			.NE(gen[7662]),

			.O(gen[7755]),
			.E(gen[7757]),

			.SO(gen[7850]),
			.S(gen[7851]),
			.SE(gen[7852]),

			.SELF(gen[7756]),
			.cell_state(gen[7756])
		); 

/******************* CELL 7757 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7757 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7661]),
			.N(gen[7662]),
			.NE(gen[7663]),

			.O(gen[7756]),
			.E(gen[7758]),

			.SO(gen[7851]),
			.S(gen[7852]),
			.SE(gen[7853]),

			.SELF(gen[7757]),
			.cell_state(gen[7757])
		); 

/******************* CELL 7758 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7758 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7662]),
			.N(gen[7663]),
			.NE(gen[7664]),

			.O(gen[7757]),
			.E(gen[7759]),

			.SO(gen[7852]),
			.S(gen[7853]),
			.SE(gen[7854]),

			.SELF(gen[7758]),
			.cell_state(gen[7758])
		); 

/******************* CELL 7759 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7759 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7663]),
			.N(gen[7664]),
			.NE(gen[7665]),

			.O(gen[7758]),
			.E(gen[7760]),

			.SO(gen[7853]),
			.S(gen[7854]),
			.SE(gen[7855]),

			.SELF(gen[7759]),
			.cell_state(gen[7759])
		); 

/******************* CELL 7760 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7760 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7664]),
			.N(gen[7665]),
			.NE(gen[7666]),

			.O(gen[7759]),
			.E(gen[7761]),

			.SO(gen[7854]),
			.S(gen[7855]),
			.SE(gen[7856]),

			.SELF(gen[7760]),
			.cell_state(gen[7760])
		); 

/******************* CELL 7761 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7761 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7665]),
			.N(gen[7666]),
			.NE(gen[7667]),

			.O(gen[7760]),
			.E(gen[7762]),

			.SO(gen[7855]),
			.S(gen[7856]),
			.SE(gen[7857]),

			.SELF(gen[7761]),
			.cell_state(gen[7761])
		); 

/******************* CELL 7762 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7762 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7666]),
			.N(gen[7667]),
			.NE(gen[7668]),

			.O(gen[7761]),
			.E(gen[7763]),

			.SO(gen[7856]),
			.S(gen[7857]),
			.SE(gen[7858]),

			.SELF(gen[7762]),
			.cell_state(gen[7762])
		); 

/******************* CELL 7763 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7763 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7667]),
			.N(gen[7668]),
			.NE(gen[7669]),

			.O(gen[7762]),
			.E(gen[7764]),

			.SO(gen[7857]),
			.S(gen[7858]),
			.SE(gen[7859]),

			.SELF(gen[7763]),
			.cell_state(gen[7763])
		); 

/******************* CELL 7764 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7764 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7668]),
			.N(gen[7669]),
			.NE(gen[7670]),

			.O(gen[7763]),
			.E(gen[7765]),

			.SO(gen[7858]),
			.S(gen[7859]),
			.SE(gen[7860]),

			.SELF(gen[7764]),
			.cell_state(gen[7764])
		); 

/******************* CELL 7765 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7765 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7669]),
			.N(gen[7670]),
			.NE(gen[7671]),

			.O(gen[7764]),
			.E(gen[7766]),

			.SO(gen[7859]),
			.S(gen[7860]),
			.SE(gen[7861]),

			.SELF(gen[7765]),
			.cell_state(gen[7765])
		); 

/******************* CELL 7766 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7766 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7670]),
			.N(gen[7671]),
			.NE(gen[7672]),

			.O(gen[7765]),
			.E(gen[7767]),

			.SO(gen[7860]),
			.S(gen[7861]),
			.SE(gen[7862]),

			.SELF(gen[7766]),
			.cell_state(gen[7766])
		); 

/******************* CELL 7767 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7767 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7671]),
			.N(gen[7672]),
			.NE(gen[7673]),

			.O(gen[7766]),
			.E(gen[7768]),

			.SO(gen[7861]),
			.S(gen[7862]),
			.SE(gen[7863]),

			.SELF(gen[7767]),
			.cell_state(gen[7767])
		); 

/******************* CELL 7768 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7768 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7672]),
			.N(gen[7673]),
			.NE(gen[7674]),

			.O(gen[7767]),
			.E(gen[7769]),

			.SO(gen[7862]),
			.S(gen[7863]),
			.SE(gen[7864]),

			.SELF(gen[7768]),
			.cell_state(gen[7768])
		); 

/******************* CELL 7769 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7769 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7673]),
			.N(gen[7674]),
			.NE(gen[7675]),

			.O(gen[7768]),
			.E(gen[7770]),

			.SO(gen[7863]),
			.S(gen[7864]),
			.SE(gen[7865]),

			.SELF(gen[7769]),
			.cell_state(gen[7769])
		); 

/******************* CELL 7770 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7770 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7674]),
			.N(gen[7675]),
			.NE(gen[7676]),

			.O(gen[7769]),
			.E(gen[7771]),

			.SO(gen[7864]),
			.S(gen[7865]),
			.SE(gen[7866]),

			.SELF(gen[7770]),
			.cell_state(gen[7770])
		); 

/******************* CELL 7771 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7771 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7675]),
			.N(gen[7676]),
			.NE(gen[7677]),

			.O(gen[7770]),
			.E(gen[7772]),

			.SO(gen[7865]),
			.S(gen[7866]),
			.SE(gen[7867]),

			.SELF(gen[7771]),
			.cell_state(gen[7771])
		); 

/******************* CELL 7772 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7772 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7676]),
			.N(gen[7677]),
			.NE(gen[7678]),

			.O(gen[7771]),
			.E(gen[7773]),

			.SO(gen[7866]),
			.S(gen[7867]),
			.SE(gen[7868]),

			.SELF(gen[7772]),
			.cell_state(gen[7772])
		); 

/******************* CELL 7773 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7773 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7677]),
			.N(gen[7678]),
			.NE(gen[7679]),

			.O(gen[7772]),
			.E(gen[7774]),

			.SO(gen[7867]),
			.S(gen[7868]),
			.SE(gen[7869]),

			.SELF(gen[7773]),
			.cell_state(gen[7773])
		); 

/******************* CELL 7774 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7774 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7678]),
			.N(gen[7679]),
			.NE(gen[7680]),

			.O(gen[7773]),
			.E(gen[7775]),

			.SO(gen[7868]),
			.S(gen[7869]),
			.SE(gen[7870]),

			.SELF(gen[7774]),
			.cell_state(gen[7774])
		); 

/******************* CELL 7775 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7775 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7679]),
			.N(gen[7680]),
			.NE(gen[7681]),

			.O(gen[7774]),
			.E(gen[7776]),

			.SO(gen[7869]),
			.S(gen[7870]),
			.SE(gen[7871]),

			.SELF(gen[7775]),
			.cell_state(gen[7775])
		); 

/******************* CELL 7776 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7776 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7680]),
			.N(gen[7681]),
			.NE(gen[7682]),

			.O(gen[7775]),
			.E(gen[7777]),

			.SO(gen[7870]),
			.S(gen[7871]),
			.SE(gen[7872]),

			.SELF(gen[7776]),
			.cell_state(gen[7776])
		); 

/******************* CELL 7777 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7777 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7681]),
			.N(gen[7682]),
			.NE(gen[7683]),

			.O(gen[7776]),
			.E(gen[7778]),

			.SO(gen[7871]),
			.S(gen[7872]),
			.SE(gen[7873]),

			.SELF(gen[7777]),
			.cell_state(gen[7777])
		); 

/******************* CELL 7778 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7778 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7682]),
			.N(gen[7683]),
			.NE(gen[7684]),

			.O(gen[7777]),
			.E(gen[7779]),

			.SO(gen[7872]),
			.S(gen[7873]),
			.SE(gen[7874]),

			.SELF(gen[7778]),
			.cell_state(gen[7778])
		); 

/******************* CELL 7779 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7779 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7683]),
			.N(gen[7684]),
			.NE(gen[7685]),

			.O(gen[7778]),
			.E(gen[7780]),

			.SO(gen[7873]),
			.S(gen[7874]),
			.SE(gen[7875]),

			.SELF(gen[7779]),
			.cell_state(gen[7779])
		); 

/******************* CELL 7780 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7780 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7684]),
			.N(gen[7685]),
			.NE(gen[7686]),

			.O(gen[7779]),
			.E(gen[7781]),

			.SO(gen[7874]),
			.S(gen[7875]),
			.SE(gen[7876]),

			.SELF(gen[7780]),
			.cell_state(gen[7780])
		); 

/******************* CELL 7781 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7781 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7685]),
			.N(gen[7686]),
			.NE(gen[7687]),

			.O(gen[7780]),
			.E(gen[7782]),

			.SO(gen[7875]),
			.S(gen[7876]),
			.SE(gen[7877]),

			.SELF(gen[7781]),
			.cell_state(gen[7781])
		); 

/******************* CELL 7782 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7782 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7686]),
			.N(gen[7687]),
			.NE(gen[7688]),

			.O(gen[7781]),
			.E(gen[7783]),

			.SO(gen[7876]),
			.S(gen[7877]),
			.SE(gen[7878]),

			.SELF(gen[7782]),
			.cell_state(gen[7782])
		); 

/******************* CELL 7783 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7783 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7687]),
			.N(gen[7688]),
			.NE(gen[7689]),

			.O(gen[7782]),
			.E(gen[7784]),

			.SO(gen[7877]),
			.S(gen[7878]),
			.SE(gen[7879]),

			.SELF(gen[7783]),
			.cell_state(gen[7783])
		); 

/******************* CELL 7784 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7784 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7688]),
			.N(gen[7689]),
			.NE(gen[7690]),

			.O(gen[7783]),
			.E(gen[7785]),

			.SO(gen[7878]),
			.S(gen[7879]),
			.SE(gen[7880]),

			.SELF(gen[7784]),
			.cell_state(gen[7784])
		); 

/******************* CELL 7785 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7785 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7689]),
			.N(gen[7690]),
			.NE(gen[7691]),

			.O(gen[7784]),
			.E(gen[7786]),

			.SO(gen[7879]),
			.S(gen[7880]),
			.SE(gen[7881]),

			.SELF(gen[7785]),
			.cell_state(gen[7785])
		); 

/******************* CELL 7786 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7786 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7690]),
			.N(gen[7691]),
			.NE(gen[7692]),

			.O(gen[7785]),
			.E(gen[7787]),

			.SO(gen[7880]),
			.S(gen[7881]),
			.SE(gen[7882]),

			.SELF(gen[7786]),
			.cell_state(gen[7786])
		); 

/******************* CELL 7787 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7787 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7691]),
			.N(gen[7692]),
			.NE(gen[7693]),

			.O(gen[7786]),
			.E(gen[7788]),

			.SO(gen[7881]),
			.S(gen[7882]),
			.SE(gen[7883]),

			.SELF(gen[7787]),
			.cell_state(gen[7787])
		); 

/******************* CELL 7788 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7788 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7692]),
			.N(gen[7693]),
			.NE(gen[7694]),

			.O(gen[7787]),
			.E(gen[7789]),

			.SO(gen[7882]),
			.S(gen[7883]),
			.SE(gen[7884]),

			.SELF(gen[7788]),
			.cell_state(gen[7788])
		); 

/******************* CELL 7789 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7789 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7693]),
			.N(gen[7694]),
			.NE(gen[7693]),

			.O(gen[7788]),
			.E(gen[7788]),

			.SO(gen[7883]),
			.S(gen[7884]),
			.SE(gen[7883]),

			.SELF(gen[7789]),
			.cell_state(gen[7789])
		); 

/******************* CELL 7790 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7790 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7696]),
			.N(gen[7695]),
			.NE(gen[7696]),

			.O(gen[7791]),
			.E(gen[7791]),

			.SO(gen[7886]),
			.S(gen[7885]),
			.SE(gen[7886]),

			.SELF(gen[7790]),
			.cell_state(gen[7790])
		); 

/******************* CELL 7791 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7791 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7695]),
			.N(gen[7696]),
			.NE(gen[7697]),

			.O(gen[7790]),
			.E(gen[7792]),

			.SO(gen[7885]),
			.S(gen[7886]),
			.SE(gen[7887]),

			.SELF(gen[7791]),
			.cell_state(gen[7791])
		); 

/******************* CELL 7792 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7792 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7696]),
			.N(gen[7697]),
			.NE(gen[7698]),

			.O(gen[7791]),
			.E(gen[7793]),

			.SO(gen[7886]),
			.S(gen[7887]),
			.SE(gen[7888]),

			.SELF(gen[7792]),
			.cell_state(gen[7792])
		); 

/******************* CELL 7793 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7793 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7697]),
			.N(gen[7698]),
			.NE(gen[7699]),

			.O(gen[7792]),
			.E(gen[7794]),

			.SO(gen[7887]),
			.S(gen[7888]),
			.SE(gen[7889]),

			.SELF(gen[7793]),
			.cell_state(gen[7793])
		); 

/******************* CELL 7794 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7794 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7698]),
			.N(gen[7699]),
			.NE(gen[7700]),

			.O(gen[7793]),
			.E(gen[7795]),

			.SO(gen[7888]),
			.S(gen[7889]),
			.SE(gen[7890]),

			.SELF(gen[7794]),
			.cell_state(gen[7794])
		); 

/******************* CELL 7795 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7795 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7699]),
			.N(gen[7700]),
			.NE(gen[7701]),

			.O(gen[7794]),
			.E(gen[7796]),

			.SO(gen[7889]),
			.S(gen[7890]),
			.SE(gen[7891]),

			.SELF(gen[7795]),
			.cell_state(gen[7795])
		); 

/******************* CELL 7796 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7796 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7700]),
			.N(gen[7701]),
			.NE(gen[7702]),

			.O(gen[7795]),
			.E(gen[7797]),

			.SO(gen[7890]),
			.S(gen[7891]),
			.SE(gen[7892]),

			.SELF(gen[7796]),
			.cell_state(gen[7796])
		); 

/******************* CELL 7797 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7797 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7701]),
			.N(gen[7702]),
			.NE(gen[7703]),

			.O(gen[7796]),
			.E(gen[7798]),

			.SO(gen[7891]),
			.S(gen[7892]),
			.SE(gen[7893]),

			.SELF(gen[7797]),
			.cell_state(gen[7797])
		); 

/******************* CELL 7798 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7798 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7702]),
			.N(gen[7703]),
			.NE(gen[7704]),

			.O(gen[7797]),
			.E(gen[7799]),

			.SO(gen[7892]),
			.S(gen[7893]),
			.SE(gen[7894]),

			.SELF(gen[7798]),
			.cell_state(gen[7798])
		); 

/******************* CELL 7799 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7799 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7703]),
			.N(gen[7704]),
			.NE(gen[7705]),

			.O(gen[7798]),
			.E(gen[7800]),

			.SO(gen[7893]),
			.S(gen[7894]),
			.SE(gen[7895]),

			.SELF(gen[7799]),
			.cell_state(gen[7799])
		); 

/******************* CELL 7800 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7800 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7704]),
			.N(gen[7705]),
			.NE(gen[7706]),

			.O(gen[7799]),
			.E(gen[7801]),

			.SO(gen[7894]),
			.S(gen[7895]),
			.SE(gen[7896]),

			.SELF(gen[7800]),
			.cell_state(gen[7800])
		); 

/******************* CELL 7801 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7801 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7705]),
			.N(gen[7706]),
			.NE(gen[7707]),

			.O(gen[7800]),
			.E(gen[7802]),

			.SO(gen[7895]),
			.S(gen[7896]),
			.SE(gen[7897]),

			.SELF(gen[7801]),
			.cell_state(gen[7801])
		); 

/******************* CELL 7802 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7802 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7706]),
			.N(gen[7707]),
			.NE(gen[7708]),

			.O(gen[7801]),
			.E(gen[7803]),

			.SO(gen[7896]),
			.S(gen[7897]),
			.SE(gen[7898]),

			.SELF(gen[7802]),
			.cell_state(gen[7802])
		); 

/******************* CELL 7803 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7803 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7707]),
			.N(gen[7708]),
			.NE(gen[7709]),

			.O(gen[7802]),
			.E(gen[7804]),

			.SO(gen[7897]),
			.S(gen[7898]),
			.SE(gen[7899]),

			.SELF(gen[7803]),
			.cell_state(gen[7803])
		); 

/******************* CELL 7804 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7804 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7708]),
			.N(gen[7709]),
			.NE(gen[7710]),

			.O(gen[7803]),
			.E(gen[7805]),

			.SO(gen[7898]),
			.S(gen[7899]),
			.SE(gen[7900]),

			.SELF(gen[7804]),
			.cell_state(gen[7804])
		); 

/******************* CELL 7805 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7805 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7709]),
			.N(gen[7710]),
			.NE(gen[7711]),

			.O(gen[7804]),
			.E(gen[7806]),

			.SO(gen[7899]),
			.S(gen[7900]),
			.SE(gen[7901]),

			.SELF(gen[7805]),
			.cell_state(gen[7805])
		); 

/******************* CELL 7806 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7806 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7710]),
			.N(gen[7711]),
			.NE(gen[7712]),

			.O(gen[7805]),
			.E(gen[7807]),

			.SO(gen[7900]),
			.S(gen[7901]),
			.SE(gen[7902]),

			.SELF(gen[7806]),
			.cell_state(gen[7806])
		); 

/******************* CELL 7807 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7807 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7711]),
			.N(gen[7712]),
			.NE(gen[7713]),

			.O(gen[7806]),
			.E(gen[7808]),

			.SO(gen[7901]),
			.S(gen[7902]),
			.SE(gen[7903]),

			.SELF(gen[7807]),
			.cell_state(gen[7807])
		); 

/******************* CELL 7808 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7808 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7712]),
			.N(gen[7713]),
			.NE(gen[7714]),

			.O(gen[7807]),
			.E(gen[7809]),

			.SO(gen[7902]),
			.S(gen[7903]),
			.SE(gen[7904]),

			.SELF(gen[7808]),
			.cell_state(gen[7808])
		); 

/******************* CELL 7809 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7809 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7713]),
			.N(gen[7714]),
			.NE(gen[7715]),

			.O(gen[7808]),
			.E(gen[7810]),

			.SO(gen[7903]),
			.S(gen[7904]),
			.SE(gen[7905]),

			.SELF(gen[7809]),
			.cell_state(gen[7809])
		); 

/******************* CELL 7810 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7810 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7714]),
			.N(gen[7715]),
			.NE(gen[7716]),

			.O(gen[7809]),
			.E(gen[7811]),

			.SO(gen[7904]),
			.S(gen[7905]),
			.SE(gen[7906]),

			.SELF(gen[7810]),
			.cell_state(gen[7810])
		); 

/******************* CELL 7811 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7811 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7715]),
			.N(gen[7716]),
			.NE(gen[7717]),

			.O(gen[7810]),
			.E(gen[7812]),

			.SO(gen[7905]),
			.S(gen[7906]),
			.SE(gen[7907]),

			.SELF(gen[7811]),
			.cell_state(gen[7811])
		); 

/******************* CELL 7812 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7812 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7716]),
			.N(gen[7717]),
			.NE(gen[7718]),

			.O(gen[7811]),
			.E(gen[7813]),

			.SO(gen[7906]),
			.S(gen[7907]),
			.SE(gen[7908]),

			.SELF(gen[7812]),
			.cell_state(gen[7812])
		); 

/******************* CELL 7813 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7813 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7717]),
			.N(gen[7718]),
			.NE(gen[7719]),

			.O(gen[7812]),
			.E(gen[7814]),

			.SO(gen[7907]),
			.S(gen[7908]),
			.SE(gen[7909]),

			.SELF(gen[7813]),
			.cell_state(gen[7813])
		); 

/******************* CELL 7814 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7814 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7718]),
			.N(gen[7719]),
			.NE(gen[7720]),

			.O(gen[7813]),
			.E(gen[7815]),

			.SO(gen[7908]),
			.S(gen[7909]),
			.SE(gen[7910]),

			.SELF(gen[7814]),
			.cell_state(gen[7814])
		); 

/******************* CELL 7815 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7815 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7719]),
			.N(gen[7720]),
			.NE(gen[7721]),

			.O(gen[7814]),
			.E(gen[7816]),

			.SO(gen[7909]),
			.S(gen[7910]),
			.SE(gen[7911]),

			.SELF(gen[7815]),
			.cell_state(gen[7815])
		); 

/******************* CELL 7816 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7816 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7720]),
			.N(gen[7721]),
			.NE(gen[7722]),

			.O(gen[7815]),
			.E(gen[7817]),

			.SO(gen[7910]),
			.S(gen[7911]),
			.SE(gen[7912]),

			.SELF(gen[7816]),
			.cell_state(gen[7816])
		); 

/******************* CELL 7817 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7817 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7721]),
			.N(gen[7722]),
			.NE(gen[7723]),

			.O(gen[7816]),
			.E(gen[7818]),

			.SO(gen[7911]),
			.S(gen[7912]),
			.SE(gen[7913]),

			.SELF(gen[7817]),
			.cell_state(gen[7817])
		); 

/******************* CELL 7818 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7818 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7722]),
			.N(gen[7723]),
			.NE(gen[7724]),

			.O(gen[7817]),
			.E(gen[7819]),

			.SO(gen[7912]),
			.S(gen[7913]),
			.SE(gen[7914]),

			.SELF(gen[7818]),
			.cell_state(gen[7818])
		); 

/******************* CELL 7819 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7819 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7723]),
			.N(gen[7724]),
			.NE(gen[7725]),

			.O(gen[7818]),
			.E(gen[7820]),

			.SO(gen[7913]),
			.S(gen[7914]),
			.SE(gen[7915]),

			.SELF(gen[7819]),
			.cell_state(gen[7819])
		); 

/******************* CELL 7820 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7820 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7724]),
			.N(gen[7725]),
			.NE(gen[7726]),

			.O(gen[7819]),
			.E(gen[7821]),

			.SO(gen[7914]),
			.S(gen[7915]),
			.SE(gen[7916]),

			.SELF(gen[7820]),
			.cell_state(gen[7820])
		); 

/******************* CELL 7821 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7821 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7725]),
			.N(gen[7726]),
			.NE(gen[7727]),

			.O(gen[7820]),
			.E(gen[7822]),

			.SO(gen[7915]),
			.S(gen[7916]),
			.SE(gen[7917]),

			.SELF(gen[7821]),
			.cell_state(gen[7821])
		); 

/******************* CELL 7822 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7822 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7726]),
			.N(gen[7727]),
			.NE(gen[7728]),

			.O(gen[7821]),
			.E(gen[7823]),

			.SO(gen[7916]),
			.S(gen[7917]),
			.SE(gen[7918]),

			.SELF(gen[7822]),
			.cell_state(gen[7822])
		); 

/******************* CELL 7823 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7823 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7727]),
			.N(gen[7728]),
			.NE(gen[7729]),

			.O(gen[7822]),
			.E(gen[7824]),

			.SO(gen[7917]),
			.S(gen[7918]),
			.SE(gen[7919]),

			.SELF(gen[7823]),
			.cell_state(gen[7823])
		); 

/******************* CELL 7824 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7824 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7728]),
			.N(gen[7729]),
			.NE(gen[7730]),

			.O(gen[7823]),
			.E(gen[7825]),

			.SO(gen[7918]),
			.S(gen[7919]),
			.SE(gen[7920]),

			.SELF(gen[7824]),
			.cell_state(gen[7824])
		); 

/******************* CELL 7825 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7825 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7729]),
			.N(gen[7730]),
			.NE(gen[7731]),

			.O(gen[7824]),
			.E(gen[7826]),

			.SO(gen[7919]),
			.S(gen[7920]),
			.SE(gen[7921]),

			.SELF(gen[7825]),
			.cell_state(gen[7825])
		); 

/******************* CELL 7826 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7826 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7730]),
			.N(gen[7731]),
			.NE(gen[7732]),

			.O(gen[7825]),
			.E(gen[7827]),

			.SO(gen[7920]),
			.S(gen[7921]),
			.SE(gen[7922]),

			.SELF(gen[7826]),
			.cell_state(gen[7826])
		); 

/******************* CELL 7827 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7827 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7731]),
			.N(gen[7732]),
			.NE(gen[7733]),

			.O(gen[7826]),
			.E(gen[7828]),

			.SO(gen[7921]),
			.S(gen[7922]),
			.SE(gen[7923]),

			.SELF(gen[7827]),
			.cell_state(gen[7827])
		); 

/******************* CELL 7828 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7828 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7732]),
			.N(gen[7733]),
			.NE(gen[7734]),

			.O(gen[7827]),
			.E(gen[7829]),

			.SO(gen[7922]),
			.S(gen[7923]),
			.SE(gen[7924]),

			.SELF(gen[7828]),
			.cell_state(gen[7828])
		); 

/******************* CELL 7829 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7829 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7733]),
			.N(gen[7734]),
			.NE(gen[7735]),

			.O(gen[7828]),
			.E(gen[7830]),

			.SO(gen[7923]),
			.S(gen[7924]),
			.SE(gen[7925]),

			.SELF(gen[7829]),
			.cell_state(gen[7829])
		); 

/******************* CELL 7830 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7830 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7734]),
			.N(gen[7735]),
			.NE(gen[7736]),

			.O(gen[7829]),
			.E(gen[7831]),

			.SO(gen[7924]),
			.S(gen[7925]),
			.SE(gen[7926]),

			.SELF(gen[7830]),
			.cell_state(gen[7830])
		); 

/******************* CELL 7831 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7831 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7735]),
			.N(gen[7736]),
			.NE(gen[7737]),

			.O(gen[7830]),
			.E(gen[7832]),

			.SO(gen[7925]),
			.S(gen[7926]),
			.SE(gen[7927]),

			.SELF(gen[7831]),
			.cell_state(gen[7831])
		); 

/******************* CELL 7832 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7832 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7736]),
			.N(gen[7737]),
			.NE(gen[7738]),

			.O(gen[7831]),
			.E(gen[7833]),

			.SO(gen[7926]),
			.S(gen[7927]),
			.SE(gen[7928]),

			.SELF(gen[7832]),
			.cell_state(gen[7832])
		); 

/******************* CELL 7833 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7833 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7737]),
			.N(gen[7738]),
			.NE(gen[7739]),

			.O(gen[7832]),
			.E(gen[7834]),

			.SO(gen[7927]),
			.S(gen[7928]),
			.SE(gen[7929]),

			.SELF(gen[7833]),
			.cell_state(gen[7833])
		); 

/******************* CELL 7834 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7834 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7738]),
			.N(gen[7739]),
			.NE(gen[7740]),

			.O(gen[7833]),
			.E(gen[7835]),

			.SO(gen[7928]),
			.S(gen[7929]),
			.SE(gen[7930]),

			.SELF(gen[7834]),
			.cell_state(gen[7834])
		); 

/******************* CELL 7835 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7835 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7739]),
			.N(gen[7740]),
			.NE(gen[7741]),

			.O(gen[7834]),
			.E(gen[7836]),

			.SO(gen[7929]),
			.S(gen[7930]),
			.SE(gen[7931]),

			.SELF(gen[7835]),
			.cell_state(gen[7835])
		); 

/******************* CELL 7836 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7836 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7740]),
			.N(gen[7741]),
			.NE(gen[7742]),

			.O(gen[7835]),
			.E(gen[7837]),

			.SO(gen[7930]),
			.S(gen[7931]),
			.SE(gen[7932]),

			.SELF(gen[7836]),
			.cell_state(gen[7836])
		); 

/******************* CELL 7837 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7837 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7741]),
			.N(gen[7742]),
			.NE(gen[7743]),

			.O(gen[7836]),
			.E(gen[7838]),

			.SO(gen[7931]),
			.S(gen[7932]),
			.SE(gen[7933]),

			.SELF(gen[7837]),
			.cell_state(gen[7837])
		); 

/******************* CELL 7838 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7838 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7742]),
			.N(gen[7743]),
			.NE(gen[7744]),

			.O(gen[7837]),
			.E(gen[7839]),

			.SO(gen[7932]),
			.S(gen[7933]),
			.SE(gen[7934]),

			.SELF(gen[7838]),
			.cell_state(gen[7838])
		); 

/******************* CELL 7839 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7839 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7743]),
			.N(gen[7744]),
			.NE(gen[7745]),

			.O(gen[7838]),
			.E(gen[7840]),

			.SO(gen[7933]),
			.S(gen[7934]),
			.SE(gen[7935]),

			.SELF(gen[7839]),
			.cell_state(gen[7839])
		); 

/******************* CELL 7840 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7840 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7744]),
			.N(gen[7745]),
			.NE(gen[7746]),

			.O(gen[7839]),
			.E(gen[7841]),

			.SO(gen[7934]),
			.S(gen[7935]),
			.SE(gen[7936]),

			.SELF(gen[7840]),
			.cell_state(gen[7840])
		); 

/******************* CELL 7841 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7841 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7745]),
			.N(gen[7746]),
			.NE(gen[7747]),

			.O(gen[7840]),
			.E(gen[7842]),

			.SO(gen[7935]),
			.S(gen[7936]),
			.SE(gen[7937]),

			.SELF(gen[7841]),
			.cell_state(gen[7841])
		); 

/******************* CELL 7842 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7842 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7746]),
			.N(gen[7747]),
			.NE(gen[7748]),

			.O(gen[7841]),
			.E(gen[7843]),

			.SO(gen[7936]),
			.S(gen[7937]),
			.SE(gen[7938]),

			.SELF(gen[7842]),
			.cell_state(gen[7842])
		); 

/******************* CELL 7843 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7843 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7747]),
			.N(gen[7748]),
			.NE(gen[7749]),

			.O(gen[7842]),
			.E(gen[7844]),

			.SO(gen[7937]),
			.S(gen[7938]),
			.SE(gen[7939]),

			.SELF(gen[7843]),
			.cell_state(gen[7843])
		); 

/******************* CELL 7844 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7844 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7748]),
			.N(gen[7749]),
			.NE(gen[7750]),

			.O(gen[7843]),
			.E(gen[7845]),

			.SO(gen[7938]),
			.S(gen[7939]),
			.SE(gen[7940]),

			.SELF(gen[7844]),
			.cell_state(gen[7844])
		); 

/******************* CELL 7845 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7845 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7749]),
			.N(gen[7750]),
			.NE(gen[7751]),

			.O(gen[7844]),
			.E(gen[7846]),

			.SO(gen[7939]),
			.S(gen[7940]),
			.SE(gen[7941]),

			.SELF(gen[7845]),
			.cell_state(gen[7845])
		); 

/******************* CELL 7846 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7846 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7750]),
			.N(gen[7751]),
			.NE(gen[7752]),

			.O(gen[7845]),
			.E(gen[7847]),

			.SO(gen[7940]),
			.S(gen[7941]),
			.SE(gen[7942]),

			.SELF(gen[7846]),
			.cell_state(gen[7846])
		); 

/******************* CELL 7847 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7847 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7751]),
			.N(gen[7752]),
			.NE(gen[7753]),

			.O(gen[7846]),
			.E(gen[7848]),

			.SO(gen[7941]),
			.S(gen[7942]),
			.SE(gen[7943]),

			.SELF(gen[7847]),
			.cell_state(gen[7847])
		); 

/******************* CELL 7848 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7848 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7752]),
			.N(gen[7753]),
			.NE(gen[7754]),

			.O(gen[7847]),
			.E(gen[7849]),

			.SO(gen[7942]),
			.S(gen[7943]),
			.SE(gen[7944]),

			.SELF(gen[7848]),
			.cell_state(gen[7848])
		); 

/******************* CELL 7849 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7849 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7753]),
			.N(gen[7754]),
			.NE(gen[7755]),

			.O(gen[7848]),
			.E(gen[7850]),

			.SO(gen[7943]),
			.S(gen[7944]),
			.SE(gen[7945]),

			.SELF(gen[7849]),
			.cell_state(gen[7849])
		); 

/******************* CELL 7850 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7850 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7754]),
			.N(gen[7755]),
			.NE(gen[7756]),

			.O(gen[7849]),
			.E(gen[7851]),

			.SO(gen[7944]),
			.S(gen[7945]),
			.SE(gen[7946]),

			.SELF(gen[7850]),
			.cell_state(gen[7850])
		); 

/******************* CELL 7851 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7851 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7755]),
			.N(gen[7756]),
			.NE(gen[7757]),

			.O(gen[7850]),
			.E(gen[7852]),

			.SO(gen[7945]),
			.S(gen[7946]),
			.SE(gen[7947]),

			.SELF(gen[7851]),
			.cell_state(gen[7851])
		); 

/******************* CELL 7852 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7852 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7756]),
			.N(gen[7757]),
			.NE(gen[7758]),

			.O(gen[7851]),
			.E(gen[7853]),

			.SO(gen[7946]),
			.S(gen[7947]),
			.SE(gen[7948]),

			.SELF(gen[7852]),
			.cell_state(gen[7852])
		); 

/******************* CELL 7853 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7853 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7757]),
			.N(gen[7758]),
			.NE(gen[7759]),

			.O(gen[7852]),
			.E(gen[7854]),

			.SO(gen[7947]),
			.S(gen[7948]),
			.SE(gen[7949]),

			.SELF(gen[7853]),
			.cell_state(gen[7853])
		); 

/******************* CELL 7854 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7854 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7758]),
			.N(gen[7759]),
			.NE(gen[7760]),

			.O(gen[7853]),
			.E(gen[7855]),

			.SO(gen[7948]),
			.S(gen[7949]),
			.SE(gen[7950]),

			.SELF(gen[7854]),
			.cell_state(gen[7854])
		); 

/******************* CELL 7855 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7855 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7759]),
			.N(gen[7760]),
			.NE(gen[7761]),

			.O(gen[7854]),
			.E(gen[7856]),

			.SO(gen[7949]),
			.S(gen[7950]),
			.SE(gen[7951]),

			.SELF(gen[7855]),
			.cell_state(gen[7855])
		); 

/******************* CELL 7856 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7856 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7760]),
			.N(gen[7761]),
			.NE(gen[7762]),

			.O(gen[7855]),
			.E(gen[7857]),

			.SO(gen[7950]),
			.S(gen[7951]),
			.SE(gen[7952]),

			.SELF(gen[7856]),
			.cell_state(gen[7856])
		); 

/******************* CELL 7857 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7857 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7761]),
			.N(gen[7762]),
			.NE(gen[7763]),

			.O(gen[7856]),
			.E(gen[7858]),

			.SO(gen[7951]),
			.S(gen[7952]),
			.SE(gen[7953]),

			.SELF(gen[7857]),
			.cell_state(gen[7857])
		); 

/******************* CELL 7858 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7858 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7762]),
			.N(gen[7763]),
			.NE(gen[7764]),

			.O(gen[7857]),
			.E(gen[7859]),

			.SO(gen[7952]),
			.S(gen[7953]),
			.SE(gen[7954]),

			.SELF(gen[7858]),
			.cell_state(gen[7858])
		); 

/******************* CELL 7859 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7859 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7763]),
			.N(gen[7764]),
			.NE(gen[7765]),

			.O(gen[7858]),
			.E(gen[7860]),

			.SO(gen[7953]),
			.S(gen[7954]),
			.SE(gen[7955]),

			.SELF(gen[7859]),
			.cell_state(gen[7859])
		); 

/******************* CELL 7860 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7860 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7764]),
			.N(gen[7765]),
			.NE(gen[7766]),

			.O(gen[7859]),
			.E(gen[7861]),

			.SO(gen[7954]),
			.S(gen[7955]),
			.SE(gen[7956]),

			.SELF(gen[7860]),
			.cell_state(gen[7860])
		); 

/******************* CELL 7861 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7861 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7765]),
			.N(gen[7766]),
			.NE(gen[7767]),

			.O(gen[7860]),
			.E(gen[7862]),

			.SO(gen[7955]),
			.S(gen[7956]),
			.SE(gen[7957]),

			.SELF(gen[7861]),
			.cell_state(gen[7861])
		); 

/******************* CELL 7862 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7862 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7766]),
			.N(gen[7767]),
			.NE(gen[7768]),

			.O(gen[7861]),
			.E(gen[7863]),

			.SO(gen[7956]),
			.S(gen[7957]),
			.SE(gen[7958]),

			.SELF(gen[7862]),
			.cell_state(gen[7862])
		); 

/******************* CELL 7863 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7863 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7767]),
			.N(gen[7768]),
			.NE(gen[7769]),

			.O(gen[7862]),
			.E(gen[7864]),

			.SO(gen[7957]),
			.S(gen[7958]),
			.SE(gen[7959]),

			.SELF(gen[7863]),
			.cell_state(gen[7863])
		); 

/******************* CELL 7864 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7864 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7768]),
			.N(gen[7769]),
			.NE(gen[7770]),

			.O(gen[7863]),
			.E(gen[7865]),

			.SO(gen[7958]),
			.S(gen[7959]),
			.SE(gen[7960]),

			.SELF(gen[7864]),
			.cell_state(gen[7864])
		); 

/******************* CELL 7865 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7865 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7769]),
			.N(gen[7770]),
			.NE(gen[7771]),

			.O(gen[7864]),
			.E(gen[7866]),

			.SO(gen[7959]),
			.S(gen[7960]),
			.SE(gen[7961]),

			.SELF(gen[7865]),
			.cell_state(gen[7865])
		); 

/******************* CELL 7866 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7866 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7770]),
			.N(gen[7771]),
			.NE(gen[7772]),

			.O(gen[7865]),
			.E(gen[7867]),

			.SO(gen[7960]),
			.S(gen[7961]),
			.SE(gen[7962]),

			.SELF(gen[7866]),
			.cell_state(gen[7866])
		); 

/******************* CELL 7867 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7867 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7771]),
			.N(gen[7772]),
			.NE(gen[7773]),

			.O(gen[7866]),
			.E(gen[7868]),

			.SO(gen[7961]),
			.S(gen[7962]),
			.SE(gen[7963]),

			.SELF(gen[7867]),
			.cell_state(gen[7867])
		); 

/******************* CELL 7868 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7868 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7772]),
			.N(gen[7773]),
			.NE(gen[7774]),

			.O(gen[7867]),
			.E(gen[7869]),

			.SO(gen[7962]),
			.S(gen[7963]),
			.SE(gen[7964]),

			.SELF(gen[7868]),
			.cell_state(gen[7868])
		); 

/******************* CELL 7869 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7869 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7773]),
			.N(gen[7774]),
			.NE(gen[7775]),

			.O(gen[7868]),
			.E(gen[7870]),

			.SO(gen[7963]),
			.S(gen[7964]),
			.SE(gen[7965]),

			.SELF(gen[7869]),
			.cell_state(gen[7869])
		); 

/******************* CELL 7870 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7870 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7774]),
			.N(gen[7775]),
			.NE(gen[7776]),

			.O(gen[7869]),
			.E(gen[7871]),

			.SO(gen[7964]),
			.S(gen[7965]),
			.SE(gen[7966]),

			.SELF(gen[7870]),
			.cell_state(gen[7870])
		); 

/******************* CELL 7871 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7871 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7775]),
			.N(gen[7776]),
			.NE(gen[7777]),

			.O(gen[7870]),
			.E(gen[7872]),

			.SO(gen[7965]),
			.S(gen[7966]),
			.SE(gen[7967]),

			.SELF(gen[7871]),
			.cell_state(gen[7871])
		); 

/******************* CELL 7872 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7872 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7776]),
			.N(gen[7777]),
			.NE(gen[7778]),

			.O(gen[7871]),
			.E(gen[7873]),

			.SO(gen[7966]),
			.S(gen[7967]),
			.SE(gen[7968]),

			.SELF(gen[7872]),
			.cell_state(gen[7872])
		); 

/******************* CELL 7873 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7873 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7777]),
			.N(gen[7778]),
			.NE(gen[7779]),

			.O(gen[7872]),
			.E(gen[7874]),

			.SO(gen[7967]),
			.S(gen[7968]),
			.SE(gen[7969]),

			.SELF(gen[7873]),
			.cell_state(gen[7873])
		); 

/******************* CELL 7874 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7874 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7778]),
			.N(gen[7779]),
			.NE(gen[7780]),

			.O(gen[7873]),
			.E(gen[7875]),

			.SO(gen[7968]),
			.S(gen[7969]),
			.SE(gen[7970]),

			.SELF(gen[7874]),
			.cell_state(gen[7874])
		); 

/******************* CELL 7875 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7875 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7779]),
			.N(gen[7780]),
			.NE(gen[7781]),

			.O(gen[7874]),
			.E(gen[7876]),

			.SO(gen[7969]),
			.S(gen[7970]),
			.SE(gen[7971]),

			.SELF(gen[7875]),
			.cell_state(gen[7875])
		); 

/******************* CELL 7876 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7876 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7780]),
			.N(gen[7781]),
			.NE(gen[7782]),

			.O(gen[7875]),
			.E(gen[7877]),

			.SO(gen[7970]),
			.S(gen[7971]),
			.SE(gen[7972]),

			.SELF(gen[7876]),
			.cell_state(gen[7876])
		); 

/******************* CELL 7877 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7877 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7781]),
			.N(gen[7782]),
			.NE(gen[7783]),

			.O(gen[7876]),
			.E(gen[7878]),

			.SO(gen[7971]),
			.S(gen[7972]),
			.SE(gen[7973]),

			.SELF(gen[7877]),
			.cell_state(gen[7877])
		); 

/******************* CELL 7878 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7878 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7782]),
			.N(gen[7783]),
			.NE(gen[7784]),

			.O(gen[7877]),
			.E(gen[7879]),

			.SO(gen[7972]),
			.S(gen[7973]),
			.SE(gen[7974]),

			.SELF(gen[7878]),
			.cell_state(gen[7878])
		); 

/******************* CELL 7879 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7879 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7783]),
			.N(gen[7784]),
			.NE(gen[7785]),

			.O(gen[7878]),
			.E(gen[7880]),

			.SO(gen[7973]),
			.S(gen[7974]),
			.SE(gen[7975]),

			.SELF(gen[7879]),
			.cell_state(gen[7879])
		); 

/******************* CELL 7880 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7880 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7784]),
			.N(gen[7785]),
			.NE(gen[7786]),

			.O(gen[7879]),
			.E(gen[7881]),

			.SO(gen[7974]),
			.S(gen[7975]),
			.SE(gen[7976]),

			.SELF(gen[7880]),
			.cell_state(gen[7880])
		); 

/******************* CELL 7881 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7881 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7785]),
			.N(gen[7786]),
			.NE(gen[7787]),

			.O(gen[7880]),
			.E(gen[7882]),

			.SO(gen[7975]),
			.S(gen[7976]),
			.SE(gen[7977]),

			.SELF(gen[7881]),
			.cell_state(gen[7881])
		); 

/******************* CELL 7882 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7882 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7786]),
			.N(gen[7787]),
			.NE(gen[7788]),

			.O(gen[7881]),
			.E(gen[7883]),

			.SO(gen[7976]),
			.S(gen[7977]),
			.SE(gen[7978]),

			.SELF(gen[7882]),
			.cell_state(gen[7882])
		); 

/******************* CELL 7883 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7883 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7787]),
			.N(gen[7788]),
			.NE(gen[7789]),

			.O(gen[7882]),
			.E(gen[7884]),

			.SO(gen[7977]),
			.S(gen[7978]),
			.SE(gen[7979]),

			.SELF(gen[7883]),
			.cell_state(gen[7883])
		); 

/******************* CELL 7884 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7884 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7788]),
			.N(gen[7789]),
			.NE(gen[7788]),

			.O(gen[7883]),
			.E(gen[7883]),

			.SO(gen[7978]),
			.S(gen[7979]),
			.SE(gen[7978]),

			.SELF(gen[7884]),
			.cell_state(gen[7884])
		); 

/******************* CELL 7885 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7885 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7791]),
			.N(gen[7790]),
			.NE(gen[7791]),

			.O(gen[7886]),
			.E(gen[7886]),

			.SO(gen[7981]),
			.S(gen[7980]),
			.SE(gen[7981]),

			.SELF(gen[7885]),
			.cell_state(gen[7885])
		); 

/******************* CELL 7886 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7886 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7790]),
			.N(gen[7791]),
			.NE(gen[7792]),

			.O(gen[7885]),
			.E(gen[7887]),

			.SO(gen[7980]),
			.S(gen[7981]),
			.SE(gen[7982]),

			.SELF(gen[7886]),
			.cell_state(gen[7886])
		); 

/******************* CELL 7887 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7887 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7791]),
			.N(gen[7792]),
			.NE(gen[7793]),

			.O(gen[7886]),
			.E(gen[7888]),

			.SO(gen[7981]),
			.S(gen[7982]),
			.SE(gen[7983]),

			.SELF(gen[7887]),
			.cell_state(gen[7887])
		); 

/******************* CELL 7888 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7888 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7792]),
			.N(gen[7793]),
			.NE(gen[7794]),

			.O(gen[7887]),
			.E(gen[7889]),

			.SO(gen[7982]),
			.S(gen[7983]),
			.SE(gen[7984]),

			.SELF(gen[7888]),
			.cell_state(gen[7888])
		); 

/******************* CELL 7889 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7889 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7793]),
			.N(gen[7794]),
			.NE(gen[7795]),

			.O(gen[7888]),
			.E(gen[7890]),

			.SO(gen[7983]),
			.S(gen[7984]),
			.SE(gen[7985]),

			.SELF(gen[7889]),
			.cell_state(gen[7889])
		); 

/******************* CELL 7890 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7890 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7794]),
			.N(gen[7795]),
			.NE(gen[7796]),

			.O(gen[7889]),
			.E(gen[7891]),

			.SO(gen[7984]),
			.S(gen[7985]),
			.SE(gen[7986]),

			.SELF(gen[7890]),
			.cell_state(gen[7890])
		); 

/******************* CELL 7891 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7891 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7795]),
			.N(gen[7796]),
			.NE(gen[7797]),

			.O(gen[7890]),
			.E(gen[7892]),

			.SO(gen[7985]),
			.S(gen[7986]),
			.SE(gen[7987]),

			.SELF(gen[7891]),
			.cell_state(gen[7891])
		); 

/******************* CELL 7892 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7892 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7796]),
			.N(gen[7797]),
			.NE(gen[7798]),

			.O(gen[7891]),
			.E(gen[7893]),

			.SO(gen[7986]),
			.S(gen[7987]),
			.SE(gen[7988]),

			.SELF(gen[7892]),
			.cell_state(gen[7892])
		); 

/******************* CELL 7893 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7893 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7797]),
			.N(gen[7798]),
			.NE(gen[7799]),

			.O(gen[7892]),
			.E(gen[7894]),

			.SO(gen[7987]),
			.S(gen[7988]),
			.SE(gen[7989]),

			.SELF(gen[7893]),
			.cell_state(gen[7893])
		); 

/******************* CELL 7894 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7894 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7798]),
			.N(gen[7799]),
			.NE(gen[7800]),

			.O(gen[7893]),
			.E(gen[7895]),

			.SO(gen[7988]),
			.S(gen[7989]),
			.SE(gen[7990]),

			.SELF(gen[7894]),
			.cell_state(gen[7894])
		); 

/******************* CELL 7895 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7895 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7799]),
			.N(gen[7800]),
			.NE(gen[7801]),

			.O(gen[7894]),
			.E(gen[7896]),

			.SO(gen[7989]),
			.S(gen[7990]),
			.SE(gen[7991]),

			.SELF(gen[7895]),
			.cell_state(gen[7895])
		); 

/******************* CELL 7896 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7896 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7800]),
			.N(gen[7801]),
			.NE(gen[7802]),

			.O(gen[7895]),
			.E(gen[7897]),

			.SO(gen[7990]),
			.S(gen[7991]),
			.SE(gen[7992]),

			.SELF(gen[7896]),
			.cell_state(gen[7896])
		); 

/******************* CELL 7897 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7897 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7801]),
			.N(gen[7802]),
			.NE(gen[7803]),

			.O(gen[7896]),
			.E(gen[7898]),

			.SO(gen[7991]),
			.S(gen[7992]),
			.SE(gen[7993]),

			.SELF(gen[7897]),
			.cell_state(gen[7897])
		); 

/******************* CELL 7898 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7898 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7802]),
			.N(gen[7803]),
			.NE(gen[7804]),

			.O(gen[7897]),
			.E(gen[7899]),

			.SO(gen[7992]),
			.S(gen[7993]),
			.SE(gen[7994]),

			.SELF(gen[7898]),
			.cell_state(gen[7898])
		); 

/******************* CELL 7899 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7899 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7803]),
			.N(gen[7804]),
			.NE(gen[7805]),

			.O(gen[7898]),
			.E(gen[7900]),

			.SO(gen[7993]),
			.S(gen[7994]),
			.SE(gen[7995]),

			.SELF(gen[7899]),
			.cell_state(gen[7899])
		); 

/******************* CELL 7900 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7900 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7804]),
			.N(gen[7805]),
			.NE(gen[7806]),

			.O(gen[7899]),
			.E(gen[7901]),

			.SO(gen[7994]),
			.S(gen[7995]),
			.SE(gen[7996]),

			.SELF(gen[7900]),
			.cell_state(gen[7900])
		); 

/******************* CELL 7901 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7901 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7805]),
			.N(gen[7806]),
			.NE(gen[7807]),

			.O(gen[7900]),
			.E(gen[7902]),

			.SO(gen[7995]),
			.S(gen[7996]),
			.SE(gen[7997]),

			.SELF(gen[7901]),
			.cell_state(gen[7901])
		); 

/******************* CELL 7902 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7902 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7806]),
			.N(gen[7807]),
			.NE(gen[7808]),

			.O(gen[7901]),
			.E(gen[7903]),

			.SO(gen[7996]),
			.S(gen[7997]),
			.SE(gen[7998]),

			.SELF(gen[7902]),
			.cell_state(gen[7902])
		); 

/******************* CELL 7903 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7903 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7807]),
			.N(gen[7808]),
			.NE(gen[7809]),

			.O(gen[7902]),
			.E(gen[7904]),

			.SO(gen[7997]),
			.S(gen[7998]),
			.SE(gen[7999]),

			.SELF(gen[7903]),
			.cell_state(gen[7903])
		); 

/******************* CELL 7904 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7904 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7808]),
			.N(gen[7809]),
			.NE(gen[7810]),

			.O(gen[7903]),
			.E(gen[7905]),

			.SO(gen[7998]),
			.S(gen[7999]),
			.SE(gen[8000]),

			.SELF(gen[7904]),
			.cell_state(gen[7904])
		); 

/******************* CELL 7905 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7905 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7809]),
			.N(gen[7810]),
			.NE(gen[7811]),

			.O(gen[7904]),
			.E(gen[7906]),

			.SO(gen[7999]),
			.S(gen[8000]),
			.SE(gen[8001]),

			.SELF(gen[7905]),
			.cell_state(gen[7905])
		); 

/******************* CELL 7906 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7906 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7810]),
			.N(gen[7811]),
			.NE(gen[7812]),

			.O(gen[7905]),
			.E(gen[7907]),

			.SO(gen[8000]),
			.S(gen[8001]),
			.SE(gen[8002]),

			.SELF(gen[7906]),
			.cell_state(gen[7906])
		); 

/******************* CELL 7907 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7907 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7811]),
			.N(gen[7812]),
			.NE(gen[7813]),

			.O(gen[7906]),
			.E(gen[7908]),

			.SO(gen[8001]),
			.S(gen[8002]),
			.SE(gen[8003]),

			.SELF(gen[7907]),
			.cell_state(gen[7907])
		); 

/******************* CELL 7908 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7908 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7812]),
			.N(gen[7813]),
			.NE(gen[7814]),

			.O(gen[7907]),
			.E(gen[7909]),

			.SO(gen[8002]),
			.S(gen[8003]),
			.SE(gen[8004]),

			.SELF(gen[7908]),
			.cell_state(gen[7908])
		); 

/******************* CELL 7909 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7909 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7813]),
			.N(gen[7814]),
			.NE(gen[7815]),

			.O(gen[7908]),
			.E(gen[7910]),

			.SO(gen[8003]),
			.S(gen[8004]),
			.SE(gen[8005]),

			.SELF(gen[7909]),
			.cell_state(gen[7909])
		); 

/******************* CELL 7910 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7910 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7814]),
			.N(gen[7815]),
			.NE(gen[7816]),

			.O(gen[7909]),
			.E(gen[7911]),

			.SO(gen[8004]),
			.S(gen[8005]),
			.SE(gen[8006]),

			.SELF(gen[7910]),
			.cell_state(gen[7910])
		); 

/******************* CELL 7911 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7911 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7815]),
			.N(gen[7816]),
			.NE(gen[7817]),

			.O(gen[7910]),
			.E(gen[7912]),

			.SO(gen[8005]),
			.S(gen[8006]),
			.SE(gen[8007]),

			.SELF(gen[7911]),
			.cell_state(gen[7911])
		); 

/******************* CELL 7912 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7912 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7816]),
			.N(gen[7817]),
			.NE(gen[7818]),

			.O(gen[7911]),
			.E(gen[7913]),

			.SO(gen[8006]),
			.S(gen[8007]),
			.SE(gen[8008]),

			.SELF(gen[7912]),
			.cell_state(gen[7912])
		); 

/******************* CELL 7913 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7913 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7817]),
			.N(gen[7818]),
			.NE(gen[7819]),

			.O(gen[7912]),
			.E(gen[7914]),

			.SO(gen[8007]),
			.S(gen[8008]),
			.SE(gen[8009]),

			.SELF(gen[7913]),
			.cell_state(gen[7913])
		); 

/******************* CELL 7914 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7914 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7818]),
			.N(gen[7819]),
			.NE(gen[7820]),

			.O(gen[7913]),
			.E(gen[7915]),

			.SO(gen[8008]),
			.S(gen[8009]),
			.SE(gen[8010]),

			.SELF(gen[7914]),
			.cell_state(gen[7914])
		); 

/******************* CELL 7915 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7915 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7819]),
			.N(gen[7820]),
			.NE(gen[7821]),

			.O(gen[7914]),
			.E(gen[7916]),

			.SO(gen[8009]),
			.S(gen[8010]),
			.SE(gen[8011]),

			.SELF(gen[7915]),
			.cell_state(gen[7915])
		); 

/******************* CELL 7916 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7916 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7820]),
			.N(gen[7821]),
			.NE(gen[7822]),

			.O(gen[7915]),
			.E(gen[7917]),

			.SO(gen[8010]),
			.S(gen[8011]),
			.SE(gen[8012]),

			.SELF(gen[7916]),
			.cell_state(gen[7916])
		); 

/******************* CELL 7917 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7917 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7821]),
			.N(gen[7822]),
			.NE(gen[7823]),

			.O(gen[7916]),
			.E(gen[7918]),

			.SO(gen[8011]),
			.S(gen[8012]),
			.SE(gen[8013]),

			.SELF(gen[7917]),
			.cell_state(gen[7917])
		); 

/******************* CELL 7918 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7918 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7822]),
			.N(gen[7823]),
			.NE(gen[7824]),

			.O(gen[7917]),
			.E(gen[7919]),

			.SO(gen[8012]),
			.S(gen[8013]),
			.SE(gen[8014]),

			.SELF(gen[7918]),
			.cell_state(gen[7918])
		); 

/******************* CELL 7919 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7919 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7823]),
			.N(gen[7824]),
			.NE(gen[7825]),

			.O(gen[7918]),
			.E(gen[7920]),

			.SO(gen[8013]),
			.S(gen[8014]),
			.SE(gen[8015]),

			.SELF(gen[7919]),
			.cell_state(gen[7919])
		); 

/******************* CELL 7920 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7920 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7824]),
			.N(gen[7825]),
			.NE(gen[7826]),

			.O(gen[7919]),
			.E(gen[7921]),

			.SO(gen[8014]),
			.S(gen[8015]),
			.SE(gen[8016]),

			.SELF(gen[7920]),
			.cell_state(gen[7920])
		); 

/******************* CELL 7921 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7921 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7825]),
			.N(gen[7826]),
			.NE(gen[7827]),

			.O(gen[7920]),
			.E(gen[7922]),

			.SO(gen[8015]),
			.S(gen[8016]),
			.SE(gen[8017]),

			.SELF(gen[7921]),
			.cell_state(gen[7921])
		); 

/******************* CELL 7922 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7922 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7826]),
			.N(gen[7827]),
			.NE(gen[7828]),

			.O(gen[7921]),
			.E(gen[7923]),

			.SO(gen[8016]),
			.S(gen[8017]),
			.SE(gen[8018]),

			.SELF(gen[7922]),
			.cell_state(gen[7922])
		); 

/******************* CELL 7923 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7923 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7827]),
			.N(gen[7828]),
			.NE(gen[7829]),

			.O(gen[7922]),
			.E(gen[7924]),

			.SO(gen[8017]),
			.S(gen[8018]),
			.SE(gen[8019]),

			.SELF(gen[7923]),
			.cell_state(gen[7923])
		); 

/******************* CELL 7924 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7924 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7828]),
			.N(gen[7829]),
			.NE(gen[7830]),

			.O(gen[7923]),
			.E(gen[7925]),

			.SO(gen[8018]),
			.S(gen[8019]),
			.SE(gen[8020]),

			.SELF(gen[7924]),
			.cell_state(gen[7924])
		); 

/******************* CELL 7925 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7925 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7829]),
			.N(gen[7830]),
			.NE(gen[7831]),

			.O(gen[7924]),
			.E(gen[7926]),

			.SO(gen[8019]),
			.S(gen[8020]),
			.SE(gen[8021]),

			.SELF(gen[7925]),
			.cell_state(gen[7925])
		); 

/******************* CELL 7926 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7926 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7830]),
			.N(gen[7831]),
			.NE(gen[7832]),

			.O(gen[7925]),
			.E(gen[7927]),

			.SO(gen[8020]),
			.S(gen[8021]),
			.SE(gen[8022]),

			.SELF(gen[7926]),
			.cell_state(gen[7926])
		); 

/******************* CELL 7927 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7927 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7831]),
			.N(gen[7832]),
			.NE(gen[7833]),

			.O(gen[7926]),
			.E(gen[7928]),

			.SO(gen[8021]),
			.S(gen[8022]),
			.SE(gen[8023]),

			.SELF(gen[7927]),
			.cell_state(gen[7927])
		); 

/******************* CELL 7928 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7928 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7832]),
			.N(gen[7833]),
			.NE(gen[7834]),

			.O(gen[7927]),
			.E(gen[7929]),

			.SO(gen[8022]),
			.S(gen[8023]),
			.SE(gen[8024]),

			.SELF(gen[7928]),
			.cell_state(gen[7928])
		); 

/******************* CELL 7929 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7929 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7833]),
			.N(gen[7834]),
			.NE(gen[7835]),

			.O(gen[7928]),
			.E(gen[7930]),

			.SO(gen[8023]),
			.S(gen[8024]),
			.SE(gen[8025]),

			.SELF(gen[7929]),
			.cell_state(gen[7929])
		); 

/******************* CELL 7930 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7930 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7834]),
			.N(gen[7835]),
			.NE(gen[7836]),

			.O(gen[7929]),
			.E(gen[7931]),

			.SO(gen[8024]),
			.S(gen[8025]),
			.SE(gen[8026]),

			.SELF(gen[7930]),
			.cell_state(gen[7930])
		); 

/******************* CELL 7931 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7931 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7835]),
			.N(gen[7836]),
			.NE(gen[7837]),

			.O(gen[7930]),
			.E(gen[7932]),

			.SO(gen[8025]),
			.S(gen[8026]),
			.SE(gen[8027]),

			.SELF(gen[7931]),
			.cell_state(gen[7931])
		); 

/******************* CELL 7932 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7932 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7836]),
			.N(gen[7837]),
			.NE(gen[7838]),

			.O(gen[7931]),
			.E(gen[7933]),

			.SO(gen[8026]),
			.S(gen[8027]),
			.SE(gen[8028]),

			.SELF(gen[7932]),
			.cell_state(gen[7932])
		); 

/******************* CELL 7933 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7933 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7837]),
			.N(gen[7838]),
			.NE(gen[7839]),

			.O(gen[7932]),
			.E(gen[7934]),

			.SO(gen[8027]),
			.S(gen[8028]),
			.SE(gen[8029]),

			.SELF(gen[7933]),
			.cell_state(gen[7933])
		); 

/******************* CELL 7934 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7934 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7838]),
			.N(gen[7839]),
			.NE(gen[7840]),

			.O(gen[7933]),
			.E(gen[7935]),

			.SO(gen[8028]),
			.S(gen[8029]),
			.SE(gen[8030]),

			.SELF(gen[7934]),
			.cell_state(gen[7934])
		); 

/******************* CELL 7935 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7935 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7839]),
			.N(gen[7840]),
			.NE(gen[7841]),

			.O(gen[7934]),
			.E(gen[7936]),

			.SO(gen[8029]),
			.S(gen[8030]),
			.SE(gen[8031]),

			.SELF(gen[7935]),
			.cell_state(gen[7935])
		); 

/******************* CELL 7936 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7936 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7840]),
			.N(gen[7841]),
			.NE(gen[7842]),

			.O(gen[7935]),
			.E(gen[7937]),

			.SO(gen[8030]),
			.S(gen[8031]),
			.SE(gen[8032]),

			.SELF(gen[7936]),
			.cell_state(gen[7936])
		); 

/******************* CELL 7937 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7937 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7841]),
			.N(gen[7842]),
			.NE(gen[7843]),

			.O(gen[7936]),
			.E(gen[7938]),

			.SO(gen[8031]),
			.S(gen[8032]),
			.SE(gen[8033]),

			.SELF(gen[7937]),
			.cell_state(gen[7937])
		); 

/******************* CELL 7938 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7938 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7842]),
			.N(gen[7843]),
			.NE(gen[7844]),

			.O(gen[7937]),
			.E(gen[7939]),

			.SO(gen[8032]),
			.S(gen[8033]),
			.SE(gen[8034]),

			.SELF(gen[7938]),
			.cell_state(gen[7938])
		); 

/******************* CELL 7939 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7939 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7843]),
			.N(gen[7844]),
			.NE(gen[7845]),

			.O(gen[7938]),
			.E(gen[7940]),

			.SO(gen[8033]),
			.S(gen[8034]),
			.SE(gen[8035]),

			.SELF(gen[7939]),
			.cell_state(gen[7939])
		); 

/******************* CELL 7940 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7940 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7844]),
			.N(gen[7845]),
			.NE(gen[7846]),

			.O(gen[7939]),
			.E(gen[7941]),

			.SO(gen[8034]),
			.S(gen[8035]),
			.SE(gen[8036]),

			.SELF(gen[7940]),
			.cell_state(gen[7940])
		); 

/******************* CELL 7941 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7941 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7845]),
			.N(gen[7846]),
			.NE(gen[7847]),

			.O(gen[7940]),
			.E(gen[7942]),

			.SO(gen[8035]),
			.S(gen[8036]),
			.SE(gen[8037]),

			.SELF(gen[7941]),
			.cell_state(gen[7941])
		); 

/******************* CELL 7942 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7942 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7846]),
			.N(gen[7847]),
			.NE(gen[7848]),

			.O(gen[7941]),
			.E(gen[7943]),

			.SO(gen[8036]),
			.S(gen[8037]),
			.SE(gen[8038]),

			.SELF(gen[7942]),
			.cell_state(gen[7942])
		); 

/******************* CELL 7943 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7943 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7847]),
			.N(gen[7848]),
			.NE(gen[7849]),

			.O(gen[7942]),
			.E(gen[7944]),

			.SO(gen[8037]),
			.S(gen[8038]),
			.SE(gen[8039]),

			.SELF(gen[7943]),
			.cell_state(gen[7943])
		); 

/******************* CELL 7944 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7944 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7848]),
			.N(gen[7849]),
			.NE(gen[7850]),

			.O(gen[7943]),
			.E(gen[7945]),

			.SO(gen[8038]),
			.S(gen[8039]),
			.SE(gen[8040]),

			.SELF(gen[7944]),
			.cell_state(gen[7944])
		); 

/******************* CELL 7945 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7945 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7849]),
			.N(gen[7850]),
			.NE(gen[7851]),

			.O(gen[7944]),
			.E(gen[7946]),

			.SO(gen[8039]),
			.S(gen[8040]),
			.SE(gen[8041]),

			.SELF(gen[7945]),
			.cell_state(gen[7945])
		); 

/******************* CELL 7946 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7946 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7850]),
			.N(gen[7851]),
			.NE(gen[7852]),

			.O(gen[7945]),
			.E(gen[7947]),

			.SO(gen[8040]),
			.S(gen[8041]),
			.SE(gen[8042]),

			.SELF(gen[7946]),
			.cell_state(gen[7946])
		); 

/******************* CELL 7947 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7947 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7851]),
			.N(gen[7852]),
			.NE(gen[7853]),

			.O(gen[7946]),
			.E(gen[7948]),

			.SO(gen[8041]),
			.S(gen[8042]),
			.SE(gen[8043]),

			.SELF(gen[7947]),
			.cell_state(gen[7947])
		); 

/******************* CELL 7948 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7948 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7852]),
			.N(gen[7853]),
			.NE(gen[7854]),

			.O(gen[7947]),
			.E(gen[7949]),

			.SO(gen[8042]),
			.S(gen[8043]),
			.SE(gen[8044]),

			.SELF(gen[7948]),
			.cell_state(gen[7948])
		); 

/******************* CELL 7949 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7949 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7853]),
			.N(gen[7854]),
			.NE(gen[7855]),

			.O(gen[7948]),
			.E(gen[7950]),

			.SO(gen[8043]),
			.S(gen[8044]),
			.SE(gen[8045]),

			.SELF(gen[7949]),
			.cell_state(gen[7949])
		); 

/******************* CELL 7950 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7950 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7854]),
			.N(gen[7855]),
			.NE(gen[7856]),

			.O(gen[7949]),
			.E(gen[7951]),

			.SO(gen[8044]),
			.S(gen[8045]),
			.SE(gen[8046]),

			.SELF(gen[7950]),
			.cell_state(gen[7950])
		); 

/******************* CELL 7951 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7951 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7855]),
			.N(gen[7856]),
			.NE(gen[7857]),

			.O(gen[7950]),
			.E(gen[7952]),

			.SO(gen[8045]),
			.S(gen[8046]),
			.SE(gen[8047]),

			.SELF(gen[7951]),
			.cell_state(gen[7951])
		); 

/******************* CELL 7952 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7952 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7856]),
			.N(gen[7857]),
			.NE(gen[7858]),

			.O(gen[7951]),
			.E(gen[7953]),

			.SO(gen[8046]),
			.S(gen[8047]),
			.SE(gen[8048]),

			.SELF(gen[7952]),
			.cell_state(gen[7952])
		); 

/******************* CELL 7953 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7953 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7857]),
			.N(gen[7858]),
			.NE(gen[7859]),

			.O(gen[7952]),
			.E(gen[7954]),

			.SO(gen[8047]),
			.S(gen[8048]),
			.SE(gen[8049]),

			.SELF(gen[7953]),
			.cell_state(gen[7953])
		); 

/******************* CELL 7954 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7954 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7858]),
			.N(gen[7859]),
			.NE(gen[7860]),

			.O(gen[7953]),
			.E(gen[7955]),

			.SO(gen[8048]),
			.S(gen[8049]),
			.SE(gen[8050]),

			.SELF(gen[7954]),
			.cell_state(gen[7954])
		); 

/******************* CELL 7955 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7955 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7859]),
			.N(gen[7860]),
			.NE(gen[7861]),

			.O(gen[7954]),
			.E(gen[7956]),

			.SO(gen[8049]),
			.S(gen[8050]),
			.SE(gen[8051]),

			.SELF(gen[7955]),
			.cell_state(gen[7955])
		); 

/******************* CELL 7956 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7956 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7860]),
			.N(gen[7861]),
			.NE(gen[7862]),

			.O(gen[7955]),
			.E(gen[7957]),

			.SO(gen[8050]),
			.S(gen[8051]),
			.SE(gen[8052]),

			.SELF(gen[7956]),
			.cell_state(gen[7956])
		); 

/******************* CELL 7957 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7957 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7861]),
			.N(gen[7862]),
			.NE(gen[7863]),

			.O(gen[7956]),
			.E(gen[7958]),

			.SO(gen[8051]),
			.S(gen[8052]),
			.SE(gen[8053]),

			.SELF(gen[7957]),
			.cell_state(gen[7957])
		); 

/******************* CELL 7958 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7958 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7862]),
			.N(gen[7863]),
			.NE(gen[7864]),

			.O(gen[7957]),
			.E(gen[7959]),

			.SO(gen[8052]),
			.S(gen[8053]),
			.SE(gen[8054]),

			.SELF(gen[7958]),
			.cell_state(gen[7958])
		); 

/******************* CELL 7959 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7959 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7863]),
			.N(gen[7864]),
			.NE(gen[7865]),

			.O(gen[7958]),
			.E(gen[7960]),

			.SO(gen[8053]),
			.S(gen[8054]),
			.SE(gen[8055]),

			.SELF(gen[7959]),
			.cell_state(gen[7959])
		); 

/******************* CELL 7960 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7960 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7864]),
			.N(gen[7865]),
			.NE(gen[7866]),

			.O(gen[7959]),
			.E(gen[7961]),

			.SO(gen[8054]),
			.S(gen[8055]),
			.SE(gen[8056]),

			.SELF(gen[7960]),
			.cell_state(gen[7960])
		); 

/******************* CELL 7961 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7961 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7865]),
			.N(gen[7866]),
			.NE(gen[7867]),

			.O(gen[7960]),
			.E(gen[7962]),

			.SO(gen[8055]),
			.S(gen[8056]),
			.SE(gen[8057]),

			.SELF(gen[7961]),
			.cell_state(gen[7961])
		); 

/******************* CELL 7962 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7962 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7866]),
			.N(gen[7867]),
			.NE(gen[7868]),

			.O(gen[7961]),
			.E(gen[7963]),

			.SO(gen[8056]),
			.S(gen[8057]),
			.SE(gen[8058]),

			.SELF(gen[7962]),
			.cell_state(gen[7962])
		); 

/******************* CELL 7963 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7963 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7867]),
			.N(gen[7868]),
			.NE(gen[7869]),

			.O(gen[7962]),
			.E(gen[7964]),

			.SO(gen[8057]),
			.S(gen[8058]),
			.SE(gen[8059]),

			.SELF(gen[7963]),
			.cell_state(gen[7963])
		); 

/******************* CELL 7964 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7964 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7868]),
			.N(gen[7869]),
			.NE(gen[7870]),

			.O(gen[7963]),
			.E(gen[7965]),

			.SO(gen[8058]),
			.S(gen[8059]),
			.SE(gen[8060]),

			.SELF(gen[7964]),
			.cell_state(gen[7964])
		); 

/******************* CELL 7965 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7965 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7869]),
			.N(gen[7870]),
			.NE(gen[7871]),

			.O(gen[7964]),
			.E(gen[7966]),

			.SO(gen[8059]),
			.S(gen[8060]),
			.SE(gen[8061]),

			.SELF(gen[7965]),
			.cell_state(gen[7965])
		); 

/******************* CELL 7966 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7966 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7870]),
			.N(gen[7871]),
			.NE(gen[7872]),

			.O(gen[7965]),
			.E(gen[7967]),

			.SO(gen[8060]),
			.S(gen[8061]),
			.SE(gen[8062]),

			.SELF(gen[7966]),
			.cell_state(gen[7966])
		); 

/******************* CELL 7967 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7967 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7871]),
			.N(gen[7872]),
			.NE(gen[7873]),

			.O(gen[7966]),
			.E(gen[7968]),

			.SO(gen[8061]),
			.S(gen[8062]),
			.SE(gen[8063]),

			.SELF(gen[7967]),
			.cell_state(gen[7967])
		); 

/******************* CELL 7968 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7968 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7872]),
			.N(gen[7873]),
			.NE(gen[7874]),

			.O(gen[7967]),
			.E(gen[7969]),

			.SO(gen[8062]),
			.S(gen[8063]),
			.SE(gen[8064]),

			.SELF(gen[7968]),
			.cell_state(gen[7968])
		); 

/******************* CELL 7969 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7969 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7873]),
			.N(gen[7874]),
			.NE(gen[7875]),

			.O(gen[7968]),
			.E(gen[7970]),

			.SO(gen[8063]),
			.S(gen[8064]),
			.SE(gen[8065]),

			.SELF(gen[7969]),
			.cell_state(gen[7969])
		); 

/******************* CELL 7970 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7970 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7874]),
			.N(gen[7875]),
			.NE(gen[7876]),

			.O(gen[7969]),
			.E(gen[7971]),

			.SO(gen[8064]),
			.S(gen[8065]),
			.SE(gen[8066]),

			.SELF(gen[7970]),
			.cell_state(gen[7970])
		); 

/******************* CELL 7971 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7971 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7875]),
			.N(gen[7876]),
			.NE(gen[7877]),

			.O(gen[7970]),
			.E(gen[7972]),

			.SO(gen[8065]),
			.S(gen[8066]),
			.SE(gen[8067]),

			.SELF(gen[7971]),
			.cell_state(gen[7971])
		); 

/******************* CELL 7972 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7972 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7876]),
			.N(gen[7877]),
			.NE(gen[7878]),

			.O(gen[7971]),
			.E(gen[7973]),

			.SO(gen[8066]),
			.S(gen[8067]),
			.SE(gen[8068]),

			.SELF(gen[7972]),
			.cell_state(gen[7972])
		); 

/******************* CELL 7973 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7973 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7877]),
			.N(gen[7878]),
			.NE(gen[7879]),

			.O(gen[7972]),
			.E(gen[7974]),

			.SO(gen[8067]),
			.S(gen[8068]),
			.SE(gen[8069]),

			.SELF(gen[7973]),
			.cell_state(gen[7973])
		); 

/******************* CELL 7974 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7974 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7878]),
			.N(gen[7879]),
			.NE(gen[7880]),

			.O(gen[7973]),
			.E(gen[7975]),

			.SO(gen[8068]),
			.S(gen[8069]),
			.SE(gen[8070]),

			.SELF(gen[7974]),
			.cell_state(gen[7974])
		); 

/******************* CELL 7975 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7975 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7879]),
			.N(gen[7880]),
			.NE(gen[7881]),

			.O(gen[7974]),
			.E(gen[7976]),

			.SO(gen[8069]),
			.S(gen[8070]),
			.SE(gen[8071]),

			.SELF(gen[7975]),
			.cell_state(gen[7975])
		); 

/******************* CELL 7976 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7976 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7880]),
			.N(gen[7881]),
			.NE(gen[7882]),

			.O(gen[7975]),
			.E(gen[7977]),

			.SO(gen[8070]),
			.S(gen[8071]),
			.SE(gen[8072]),

			.SELF(gen[7976]),
			.cell_state(gen[7976])
		); 

/******************* CELL 7977 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7977 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7881]),
			.N(gen[7882]),
			.NE(gen[7883]),

			.O(gen[7976]),
			.E(gen[7978]),

			.SO(gen[8071]),
			.S(gen[8072]),
			.SE(gen[8073]),

			.SELF(gen[7977]),
			.cell_state(gen[7977])
		); 

/******************* CELL 7978 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7978 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7882]),
			.N(gen[7883]),
			.NE(gen[7884]),

			.O(gen[7977]),
			.E(gen[7979]),

			.SO(gen[8072]),
			.S(gen[8073]),
			.SE(gen[8074]),

			.SELF(gen[7978]),
			.cell_state(gen[7978])
		); 

/******************* CELL 7979 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7979 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7883]),
			.N(gen[7884]),
			.NE(gen[7883]),

			.O(gen[7978]),
			.E(gen[7978]),

			.SO(gen[8073]),
			.S(gen[8074]),
			.SE(gen[8073]),

			.SELF(gen[7979]),
			.cell_state(gen[7979])
		); 

/******************* CELL 7980 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7980 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7886]),
			.N(gen[7885]),
			.NE(gen[7886]),

			.O(gen[7981]),
			.E(gen[7981]),

			.SO(gen[8076]),
			.S(gen[8075]),
			.SE(gen[8076]),

			.SELF(gen[7980]),
			.cell_state(gen[7980])
		); 

/******************* CELL 7981 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7981 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7885]),
			.N(gen[7886]),
			.NE(gen[7887]),

			.O(gen[7980]),
			.E(gen[7982]),

			.SO(gen[8075]),
			.S(gen[8076]),
			.SE(gen[8077]),

			.SELF(gen[7981]),
			.cell_state(gen[7981])
		); 

/******************* CELL 7982 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7982 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7886]),
			.N(gen[7887]),
			.NE(gen[7888]),

			.O(gen[7981]),
			.E(gen[7983]),

			.SO(gen[8076]),
			.S(gen[8077]),
			.SE(gen[8078]),

			.SELF(gen[7982]),
			.cell_state(gen[7982])
		); 

/******************* CELL 7983 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7983 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7887]),
			.N(gen[7888]),
			.NE(gen[7889]),

			.O(gen[7982]),
			.E(gen[7984]),

			.SO(gen[8077]),
			.S(gen[8078]),
			.SE(gen[8079]),

			.SELF(gen[7983]),
			.cell_state(gen[7983])
		); 

/******************* CELL 7984 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7984 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7888]),
			.N(gen[7889]),
			.NE(gen[7890]),

			.O(gen[7983]),
			.E(gen[7985]),

			.SO(gen[8078]),
			.S(gen[8079]),
			.SE(gen[8080]),

			.SELF(gen[7984]),
			.cell_state(gen[7984])
		); 

/******************* CELL 7985 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7985 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7889]),
			.N(gen[7890]),
			.NE(gen[7891]),

			.O(gen[7984]),
			.E(gen[7986]),

			.SO(gen[8079]),
			.S(gen[8080]),
			.SE(gen[8081]),

			.SELF(gen[7985]),
			.cell_state(gen[7985])
		); 

/******************* CELL 7986 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7986 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7890]),
			.N(gen[7891]),
			.NE(gen[7892]),

			.O(gen[7985]),
			.E(gen[7987]),

			.SO(gen[8080]),
			.S(gen[8081]),
			.SE(gen[8082]),

			.SELF(gen[7986]),
			.cell_state(gen[7986])
		); 

/******************* CELL 7987 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7987 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7891]),
			.N(gen[7892]),
			.NE(gen[7893]),

			.O(gen[7986]),
			.E(gen[7988]),

			.SO(gen[8081]),
			.S(gen[8082]),
			.SE(gen[8083]),

			.SELF(gen[7987]),
			.cell_state(gen[7987])
		); 

/******************* CELL 7988 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7988 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7892]),
			.N(gen[7893]),
			.NE(gen[7894]),

			.O(gen[7987]),
			.E(gen[7989]),

			.SO(gen[8082]),
			.S(gen[8083]),
			.SE(gen[8084]),

			.SELF(gen[7988]),
			.cell_state(gen[7988])
		); 

/******************* CELL 7989 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7989 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7893]),
			.N(gen[7894]),
			.NE(gen[7895]),

			.O(gen[7988]),
			.E(gen[7990]),

			.SO(gen[8083]),
			.S(gen[8084]),
			.SE(gen[8085]),

			.SELF(gen[7989]),
			.cell_state(gen[7989])
		); 

/******************* CELL 7990 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7990 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7894]),
			.N(gen[7895]),
			.NE(gen[7896]),

			.O(gen[7989]),
			.E(gen[7991]),

			.SO(gen[8084]),
			.S(gen[8085]),
			.SE(gen[8086]),

			.SELF(gen[7990]),
			.cell_state(gen[7990])
		); 

/******************* CELL 7991 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7991 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7895]),
			.N(gen[7896]),
			.NE(gen[7897]),

			.O(gen[7990]),
			.E(gen[7992]),

			.SO(gen[8085]),
			.S(gen[8086]),
			.SE(gen[8087]),

			.SELF(gen[7991]),
			.cell_state(gen[7991])
		); 

/******************* CELL 7992 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7992 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7896]),
			.N(gen[7897]),
			.NE(gen[7898]),

			.O(gen[7991]),
			.E(gen[7993]),

			.SO(gen[8086]),
			.S(gen[8087]),
			.SE(gen[8088]),

			.SELF(gen[7992]),
			.cell_state(gen[7992])
		); 

/******************* CELL 7993 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7993 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7897]),
			.N(gen[7898]),
			.NE(gen[7899]),

			.O(gen[7992]),
			.E(gen[7994]),

			.SO(gen[8087]),
			.S(gen[8088]),
			.SE(gen[8089]),

			.SELF(gen[7993]),
			.cell_state(gen[7993])
		); 

/******************* CELL 7994 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7994 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7898]),
			.N(gen[7899]),
			.NE(gen[7900]),

			.O(gen[7993]),
			.E(gen[7995]),

			.SO(gen[8088]),
			.S(gen[8089]),
			.SE(gen[8090]),

			.SELF(gen[7994]),
			.cell_state(gen[7994])
		); 

/******************* CELL 7995 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7995 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7899]),
			.N(gen[7900]),
			.NE(gen[7901]),

			.O(gen[7994]),
			.E(gen[7996]),

			.SO(gen[8089]),
			.S(gen[8090]),
			.SE(gen[8091]),

			.SELF(gen[7995]),
			.cell_state(gen[7995])
		); 

/******************* CELL 7996 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7996 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7900]),
			.N(gen[7901]),
			.NE(gen[7902]),

			.O(gen[7995]),
			.E(gen[7997]),

			.SO(gen[8090]),
			.S(gen[8091]),
			.SE(gen[8092]),

			.SELF(gen[7996]),
			.cell_state(gen[7996])
		); 

/******************* CELL 7997 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7997 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7901]),
			.N(gen[7902]),
			.NE(gen[7903]),

			.O(gen[7996]),
			.E(gen[7998]),

			.SO(gen[8091]),
			.S(gen[8092]),
			.SE(gen[8093]),

			.SELF(gen[7997]),
			.cell_state(gen[7997])
		); 

/******************* CELL 7998 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7998 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7902]),
			.N(gen[7903]),
			.NE(gen[7904]),

			.O(gen[7997]),
			.E(gen[7999]),

			.SO(gen[8092]),
			.S(gen[8093]),
			.SE(gen[8094]),

			.SELF(gen[7998]),
			.cell_state(gen[7998])
		); 

/******************* CELL 7999 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell7999 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7903]),
			.N(gen[7904]),
			.NE(gen[7905]),

			.O(gen[7998]),
			.E(gen[8000]),

			.SO(gen[8093]),
			.S(gen[8094]),
			.SE(gen[8095]),

			.SELF(gen[7999]),
			.cell_state(gen[7999])
		); 

/******************* CELL 8000 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8000 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7904]),
			.N(gen[7905]),
			.NE(gen[7906]),

			.O(gen[7999]),
			.E(gen[8001]),

			.SO(gen[8094]),
			.S(gen[8095]),
			.SE(gen[8096]),

			.SELF(gen[8000]),
			.cell_state(gen[8000])
		); 

/******************* CELL 8001 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8001 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7905]),
			.N(gen[7906]),
			.NE(gen[7907]),

			.O(gen[8000]),
			.E(gen[8002]),

			.SO(gen[8095]),
			.S(gen[8096]),
			.SE(gen[8097]),

			.SELF(gen[8001]),
			.cell_state(gen[8001])
		); 

/******************* CELL 8002 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8002 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7906]),
			.N(gen[7907]),
			.NE(gen[7908]),

			.O(gen[8001]),
			.E(gen[8003]),

			.SO(gen[8096]),
			.S(gen[8097]),
			.SE(gen[8098]),

			.SELF(gen[8002]),
			.cell_state(gen[8002])
		); 

/******************* CELL 8003 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8003 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7907]),
			.N(gen[7908]),
			.NE(gen[7909]),

			.O(gen[8002]),
			.E(gen[8004]),

			.SO(gen[8097]),
			.S(gen[8098]),
			.SE(gen[8099]),

			.SELF(gen[8003]),
			.cell_state(gen[8003])
		); 

/******************* CELL 8004 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8004 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7908]),
			.N(gen[7909]),
			.NE(gen[7910]),

			.O(gen[8003]),
			.E(gen[8005]),

			.SO(gen[8098]),
			.S(gen[8099]),
			.SE(gen[8100]),

			.SELF(gen[8004]),
			.cell_state(gen[8004])
		); 

/******************* CELL 8005 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8005 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7909]),
			.N(gen[7910]),
			.NE(gen[7911]),

			.O(gen[8004]),
			.E(gen[8006]),

			.SO(gen[8099]),
			.S(gen[8100]),
			.SE(gen[8101]),

			.SELF(gen[8005]),
			.cell_state(gen[8005])
		); 

/******************* CELL 8006 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8006 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7910]),
			.N(gen[7911]),
			.NE(gen[7912]),

			.O(gen[8005]),
			.E(gen[8007]),

			.SO(gen[8100]),
			.S(gen[8101]),
			.SE(gen[8102]),

			.SELF(gen[8006]),
			.cell_state(gen[8006])
		); 

/******************* CELL 8007 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8007 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7911]),
			.N(gen[7912]),
			.NE(gen[7913]),

			.O(gen[8006]),
			.E(gen[8008]),

			.SO(gen[8101]),
			.S(gen[8102]),
			.SE(gen[8103]),

			.SELF(gen[8007]),
			.cell_state(gen[8007])
		); 

/******************* CELL 8008 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8008 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7912]),
			.N(gen[7913]),
			.NE(gen[7914]),

			.O(gen[8007]),
			.E(gen[8009]),

			.SO(gen[8102]),
			.S(gen[8103]),
			.SE(gen[8104]),

			.SELF(gen[8008]),
			.cell_state(gen[8008])
		); 

/******************* CELL 8009 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8009 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7913]),
			.N(gen[7914]),
			.NE(gen[7915]),

			.O(gen[8008]),
			.E(gen[8010]),

			.SO(gen[8103]),
			.S(gen[8104]),
			.SE(gen[8105]),

			.SELF(gen[8009]),
			.cell_state(gen[8009])
		); 

/******************* CELL 8010 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8010 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7914]),
			.N(gen[7915]),
			.NE(gen[7916]),

			.O(gen[8009]),
			.E(gen[8011]),

			.SO(gen[8104]),
			.S(gen[8105]),
			.SE(gen[8106]),

			.SELF(gen[8010]),
			.cell_state(gen[8010])
		); 

/******************* CELL 8011 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8011 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7915]),
			.N(gen[7916]),
			.NE(gen[7917]),

			.O(gen[8010]),
			.E(gen[8012]),

			.SO(gen[8105]),
			.S(gen[8106]),
			.SE(gen[8107]),

			.SELF(gen[8011]),
			.cell_state(gen[8011])
		); 

/******************* CELL 8012 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8012 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7916]),
			.N(gen[7917]),
			.NE(gen[7918]),

			.O(gen[8011]),
			.E(gen[8013]),

			.SO(gen[8106]),
			.S(gen[8107]),
			.SE(gen[8108]),

			.SELF(gen[8012]),
			.cell_state(gen[8012])
		); 

/******************* CELL 8013 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8013 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7917]),
			.N(gen[7918]),
			.NE(gen[7919]),

			.O(gen[8012]),
			.E(gen[8014]),

			.SO(gen[8107]),
			.S(gen[8108]),
			.SE(gen[8109]),

			.SELF(gen[8013]),
			.cell_state(gen[8013])
		); 

/******************* CELL 8014 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8014 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7918]),
			.N(gen[7919]),
			.NE(gen[7920]),

			.O(gen[8013]),
			.E(gen[8015]),

			.SO(gen[8108]),
			.S(gen[8109]),
			.SE(gen[8110]),

			.SELF(gen[8014]),
			.cell_state(gen[8014])
		); 

/******************* CELL 8015 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8015 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7919]),
			.N(gen[7920]),
			.NE(gen[7921]),

			.O(gen[8014]),
			.E(gen[8016]),

			.SO(gen[8109]),
			.S(gen[8110]),
			.SE(gen[8111]),

			.SELF(gen[8015]),
			.cell_state(gen[8015])
		); 

/******************* CELL 8016 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8016 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7920]),
			.N(gen[7921]),
			.NE(gen[7922]),

			.O(gen[8015]),
			.E(gen[8017]),

			.SO(gen[8110]),
			.S(gen[8111]),
			.SE(gen[8112]),

			.SELF(gen[8016]),
			.cell_state(gen[8016])
		); 

/******************* CELL 8017 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8017 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7921]),
			.N(gen[7922]),
			.NE(gen[7923]),

			.O(gen[8016]),
			.E(gen[8018]),

			.SO(gen[8111]),
			.S(gen[8112]),
			.SE(gen[8113]),

			.SELF(gen[8017]),
			.cell_state(gen[8017])
		); 

/******************* CELL 8018 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8018 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7922]),
			.N(gen[7923]),
			.NE(gen[7924]),

			.O(gen[8017]),
			.E(gen[8019]),

			.SO(gen[8112]),
			.S(gen[8113]),
			.SE(gen[8114]),

			.SELF(gen[8018]),
			.cell_state(gen[8018])
		); 

/******************* CELL 8019 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8019 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7923]),
			.N(gen[7924]),
			.NE(gen[7925]),

			.O(gen[8018]),
			.E(gen[8020]),

			.SO(gen[8113]),
			.S(gen[8114]),
			.SE(gen[8115]),

			.SELF(gen[8019]),
			.cell_state(gen[8019])
		); 

/******************* CELL 8020 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8020 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7924]),
			.N(gen[7925]),
			.NE(gen[7926]),

			.O(gen[8019]),
			.E(gen[8021]),

			.SO(gen[8114]),
			.S(gen[8115]),
			.SE(gen[8116]),

			.SELF(gen[8020]),
			.cell_state(gen[8020])
		); 

/******************* CELL 8021 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8021 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7925]),
			.N(gen[7926]),
			.NE(gen[7927]),

			.O(gen[8020]),
			.E(gen[8022]),

			.SO(gen[8115]),
			.S(gen[8116]),
			.SE(gen[8117]),

			.SELF(gen[8021]),
			.cell_state(gen[8021])
		); 

/******************* CELL 8022 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8022 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7926]),
			.N(gen[7927]),
			.NE(gen[7928]),

			.O(gen[8021]),
			.E(gen[8023]),

			.SO(gen[8116]),
			.S(gen[8117]),
			.SE(gen[8118]),

			.SELF(gen[8022]),
			.cell_state(gen[8022])
		); 

/******************* CELL 8023 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8023 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7927]),
			.N(gen[7928]),
			.NE(gen[7929]),

			.O(gen[8022]),
			.E(gen[8024]),

			.SO(gen[8117]),
			.S(gen[8118]),
			.SE(gen[8119]),

			.SELF(gen[8023]),
			.cell_state(gen[8023])
		); 

/******************* CELL 8024 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8024 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7928]),
			.N(gen[7929]),
			.NE(gen[7930]),

			.O(gen[8023]),
			.E(gen[8025]),

			.SO(gen[8118]),
			.S(gen[8119]),
			.SE(gen[8120]),

			.SELF(gen[8024]),
			.cell_state(gen[8024])
		); 

/******************* CELL 8025 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8025 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7929]),
			.N(gen[7930]),
			.NE(gen[7931]),

			.O(gen[8024]),
			.E(gen[8026]),

			.SO(gen[8119]),
			.S(gen[8120]),
			.SE(gen[8121]),

			.SELF(gen[8025]),
			.cell_state(gen[8025])
		); 

/******************* CELL 8026 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8026 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7930]),
			.N(gen[7931]),
			.NE(gen[7932]),

			.O(gen[8025]),
			.E(gen[8027]),

			.SO(gen[8120]),
			.S(gen[8121]),
			.SE(gen[8122]),

			.SELF(gen[8026]),
			.cell_state(gen[8026])
		); 

/******************* CELL 8027 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8027 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7931]),
			.N(gen[7932]),
			.NE(gen[7933]),

			.O(gen[8026]),
			.E(gen[8028]),

			.SO(gen[8121]),
			.S(gen[8122]),
			.SE(gen[8123]),

			.SELF(gen[8027]),
			.cell_state(gen[8027])
		); 

/******************* CELL 8028 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8028 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7932]),
			.N(gen[7933]),
			.NE(gen[7934]),

			.O(gen[8027]),
			.E(gen[8029]),

			.SO(gen[8122]),
			.S(gen[8123]),
			.SE(gen[8124]),

			.SELF(gen[8028]),
			.cell_state(gen[8028])
		); 

/******************* CELL 8029 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8029 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7933]),
			.N(gen[7934]),
			.NE(gen[7935]),

			.O(gen[8028]),
			.E(gen[8030]),

			.SO(gen[8123]),
			.S(gen[8124]),
			.SE(gen[8125]),

			.SELF(gen[8029]),
			.cell_state(gen[8029])
		); 

/******************* CELL 8030 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8030 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7934]),
			.N(gen[7935]),
			.NE(gen[7936]),

			.O(gen[8029]),
			.E(gen[8031]),

			.SO(gen[8124]),
			.S(gen[8125]),
			.SE(gen[8126]),

			.SELF(gen[8030]),
			.cell_state(gen[8030])
		); 

/******************* CELL 8031 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8031 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7935]),
			.N(gen[7936]),
			.NE(gen[7937]),

			.O(gen[8030]),
			.E(gen[8032]),

			.SO(gen[8125]),
			.S(gen[8126]),
			.SE(gen[8127]),

			.SELF(gen[8031]),
			.cell_state(gen[8031])
		); 

/******************* CELL 8032 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8032 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7936]),
			.N(gen[7937]),
			.NE(gen[7938]),

			.O(gen[8031]),
			.E(gen[8033]),

			.SO(gen[8126]),
			.S(gen[8127]),
			.SE(gen[8128]),

			.SELF(gen[8032]),
			.cell_state(gen[8032])
		); 

/******************* CELL 8033 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8033 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7937]),
			.N(gen[7938]),
			.NE(gen[7939]),

			.O(gen[8032]),
			.E(gen[8034]),

			.SO(gen[8127]),
			.S(gen[8128]),
			.SE(gen[8129]),

			.SELF(gen[8033]),
			.cell_state(gen[8033])
		); 

/******************* CELL 8034 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8034 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7938]),
			.N(gen[7939]),
			.NE(gen[7940]),

			.O(gen[8033]),
			.E(gen[8035]),

			.SO(gen[8128]),
			.S(gen[8129]),
			.SE(gen[8130]),

			.SELF(gen[8034]),
			.cell_state(gen[8034])
		); 

/******************* CELL 8035 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8035 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7939]),
			.N(gen[7940]),
			.NE(gen[7941]),

			.O(gen[8034]),
			.E(gen[8036]),

			.SO(gen[8129]),
			.S(gen[8130]),
			.SE(gen[8131]),

			.SELF(gen[8035]),
			.cell_state(gen[8035])
		); 

/******************* CELL 8036 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8036 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7940]),
			.N(gen[7941]),
			.NE(gen[7942]),

			.O(gen[8035]),
			.E(gen[8037]),

			.SO(gen[8130]),
			.S(gen[8131]),
			.SE(gen[8132]),

			.SELF(gen[8036]),
			.cell_state(gen[8036])
		); 

/******************* CELL 8037 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8037 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7941]),
			.N(gen[7942]),
			.NE(gen[7943]),

			.O(gen[8036]),
			.E(gen[8038]),

			.SO(gen[8131]),
			.S(gen[8132]),
			.SE(gen[8133]),

			.SELF(gen[8037]),
			.cell_state(gen[8037])
		); 

/******************* CELL 8038 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8038 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7942]),
			.N(gen[7943]),
			.NE(gen[7944]),

			.O(gen[8037]),
			.E(gen[8039]),

			.SO(gen[8132]),
			.S(gen[8133]),
			.SE(gen[8134]),

			.SELF(gen[8038]),
			.cell_state(gen[8038])
		); 

/******************* CELL 8039 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8039 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7943]),
			.N(gen[7944]),
			.NE(gen[7945]),

			.O(gen[8038]),
			.E(gen[8040]),

			.SO(gen[8133]),
			.S(gen[8134]),
			.SE(gen[8135]),

			.SELF(gen[8039]),
			.cell_state(gen[8039])
		); 

/******************* CELL 8040 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8040 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7944]),
			.N(gen[7945]),
			.NE(gen[7946]),

			.O(gen[8039]),
			.E(gen[8041]),

			.SO(gen[8134]),
			.S(gen[8135]),
			.SE(gen[8136]),

			.SELF(gen[8040]),
			.cell_state(gen[8040])
		); 

/******************* CELL 8041 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8041 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7945]),
			.N(gen[7946]),
			.NE(gen[7947]),

			.O(gen[8040]),
			.E(gen[8042]),

			.SO(gen[8135]),
			.S(gen[8136]),
			.SE(gen[8137]),

			.SELF(gen[8041]),
			.cell_state(gen[8041])
		); 

/******************* CELL 8042 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8042 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7946]),
			.N(gen[7947]),
			.NE(gen[7948]),

			.O(gen[8041]),
			.E(gen[8043]),

			.SO(gen[8136]),
			.S(gen[8137]),
			.SE(gen[8138]),

			.SELF(gen[8042]),
			.cell_state(gen[8042])
		); 

/******************* CELL 8043 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8043 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7947]),
			.N(gen[7948]),
			.NE(gen[7949]),

			.O(gen[8042]),
			.E(gen[8044]),

			.SO(gen[8137]),
			.S(gen[8138]),
			.SE(gen[8139]),

			.SELF(gen[8043]),
			.cell_state(gen[8043])
		); 

/******************* CELL 8044 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8044 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7948]),
			.N(gen[7949]),
			.NE(gen[7950]),

			.O(gen[8043]),
			.E(gen[8045]),

			.SO(gen[8138]),
			.S(gen[8139]),
			.SE(gen[8140]),

			.SELF(gen[8044]),
			.cell_state(gen[8044])
		); 

/******************* CELL 8045 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8045 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7949]),
			.N(gen[7950]),
			.NE(gen[7951]),

			.O(gen[8044]),
			.E(gen[8046]),

			.SO(gen[8139]),
			.S(gen[8140]),
			.SE(gen[8141]),

			.SELF(gen[8045]),
			.cell_state(gen[8045])
		); 

/******************* CELL 8046 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8046 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7950]),
			.N(gen[7951]),
			.NE(gen[7952]),

			.O(gen[8045]),
			.E(gen[8047]),

			.SO(gen[8140]),
			.S(gen[8141]),
			.SE(gen[8142]),

			.SELF(gen[8046]),
			.cell_state(gen[8046])
		); 

/******************* CELL 8047 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8047 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7951]),
			.N(gen[7952]),
			.NE(gen[7953]),

			.O(gen[8046]),
			.E(gen[8048]),

			.SO(gen[8141]),
			.S(gen[8142]),
			.SE(gen[8143]),

			.SELF(gen[8047]),
			.cell_state(gen[8047])
		); 

/******************* CELL 8048 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8048 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7952]),
			.N(gen[7953]),
			.NE(gen[7954]),

			.O(gen[8047]),
			.E(gen[8049]),

			.SO(gen[8142]),
			.S(gen[8143]),
			.SE(gen[8144]),

			.SELF(gen[8048]),
			.cell_state(gen[8048])
		); 

/******************* CELL 8049 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8049 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7953]),
			.N(gen[7954]),
			.NE(gen[7955]),

			.O(gen[8048]),
			.E(gen[8050]),

			.SO(gen[8143]),
			.S(gen[8144]),
			.SE(gen[8145]),

			.SELF(gen[8049]),
			.cell_state(gen[8049])
		); 

/******************* CELL 8050 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8050 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7954]),
			.N(gen[7955]),
			.NE(gen[7956]),

			.O(gen[8049]),
			.E(gen[8051]),

			.SO(gen[8144]),
			.S(gen[8145]),
			.SE(gen[8146]),

			.SELF(gen[8050]),
			.cell_state(gen[8050])
		); 

/******************* CELL 8051 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8051 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7955]),
			.N(gen[7956]),
			.NE(gen[7957]),

			.O(gen[8050]),
			.E(gen[8052]),

			.SO(gen[8145]),
			.S(gen[8146]),
			.SE(gen[8147]),

			.SELF(gen[8051]),
			.cell_state(gen[8051])
		); 

/******************* CELL 8052 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8052 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7956]),
			.N(gen[7957]),
			.NE(gen[7958]),

			.O(gen[8051]),
			.E(gen[8053]),

			.SO(gen[8146]),
			.S(gen[8147]),
			.SE(gen[8148]),

			.SELF(gen[8052]),
			.cell_state(gen[8052])
		); 

/******************* CELL 8053 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8053 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7957]),
			.N(gen[7958]),
			.NE(gen[7959]),

			.O(gen[8052]),
			.E(gen[8054]),

			.SO(gen[8147]),
			.S(gen[8148]),
			.SE(gen[8149]),

			.SELF(gen[8053]),
			.cell_state(gen[8053])
		); 

/******************* CELL 8054 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8054 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7958]),
			.N(gen[7959]),
			.NE(gen[7960]),

			.O(gen[8053]),
			.E(gen[8055]),

			.SO(gen[8148]),
			.S(gen[8149]),
			.SE(gen[8150]),

			.SELF(gen[8054]),
			.cell_state(gen[8054])
		); 

/******************* CELL 8055 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8055 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7959]),
			.N(gen[7960]),
			.NE(gen[7961]),

			.O(gen[8054]),
			.E(gen[8056]),

			.SO(gen[8149]),
			.S(gen[8150]),
			.SE(gen[8151]),

			.SELF(gen[8055]),
			.cell_state(gen[8055])
		); 

/******************* CELL 8056 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8056 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7960]),
			.N(gen[7961]),
			.NE(gen[7962]),

			.O(gen[8055]),
			.E(gen[8057]),

			.SO(gen[8150]),
			.S(gen[8151]),
			.SE(gen[8152]),

			.SELF(gen[8056]),
			.cell_state(gen[8056])
		); 

/******************* CELL 8057 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8057 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7961]),
			.N(gen[7962]),
			.NE(gen[7963]),

			.O(gen[8056]),
			.E(gen[8058]),

			.SO(gen[8151]),
			.S(gen[8152]),
			.SE(gen[8153]),

			.SELF(gen[8057]),
			.cell_state(gen[8057])
		); 

/******************* CELL 8058 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8058 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7962]),
			.N(gen[7963]),
			.NE(gen[7964]),

			.O(gen[8057]),
			.E(gen[8059]),

			.SO(gen[8152]),
			.S(gen[8153]),
			.SE(gen[8154]),

			.SELF(gen[8058]),
			.cell_state(gen[8058])
		); 

/******************* CELL 8059 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8059 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7963]),
			.N(gen[7964]),
			.NE(gen[7965]),

			.O(gen[8058]),
			.E(gen[8060]),

			.SO(gen[8153]),
			.S(gen[8154]),
			.SE(gen[8155]),

			.SELF(gen[8059]),
			.cell_state(gen[8059])
		); 

/******************* CELL 8060 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8060 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7964]),
			.N(gen[7965]),
			.NE(gen[7966]),

			.O(gen[8059]),
			.E(gen[8061]),

			.SO(gen[8154]),
			.S(gen[8155]),
			.SE(gen[8156]),

			.SELF(gen[8060]),
			.cell_state(gen[8060])
		); 

/******************* CELL 8061 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8061 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7965]),
			.N(gen[7966]),
			.NE(gen[7967]),

			.O(gen[8060]),
			.E(gen[8062]),

			.SO(gen[8155]),
			.S(gen[8156]),
			.SE(gen[8157]),

			.SELF(gen[8061]),
			.cell_state(gen[8061])
		); 

/******************* CELL 8062 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8062 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7966]),
			.N(gen[7967]),
			.NE(gen[7968]),

			.O(gen[8061]),
			.E(gen[8063]),

			.SO(gen[8156]),
			.S(gen[8157]),
			.SE(gen[8158]),

			.SELF(gen[8062]),
			.cell_state(gen[8062])
		); 

/******************* CELL 8063 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8063 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7967]),
			.N(gen[7968]),
			.NE(gen[7969]),

			.O(gen[8062]),
			.E(gen[8064]),

			.SO(gen[8157]),
			.S(gen[8158]),
			.SE(gen[8159]),

			.SELF(gen[8063]),
			.cell_state(gen[8063])
		); 

/******************* CELL 8064 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8064 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7968]),
			.N(gen[7969]),
			.NE(gen[7970]),

			.O(gen[8063]),
			.E(gen[8065]),

			.SO(gen[8158]),
			.S(gen[8159]),
			.SE(gen[8160]),

			.SELF(gen[8064]),
			.cell_state(gen[8064])
		); 

/******************* CELL 8065 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8065 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7969]),
			.N(gen[7970]),
			.NE(gen[7971]),

			.O(gen[8064]),
			.E(gen[8066]),

			.SO(gen[8159]),
			.S(gen[8160]),
			.SE(gen[8161]),

			.SELF(gen[8065]),
			.cell_state(gen[8065])
		); 

/******************* CELL 8066 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8066 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7970]),
			.N(gen[7971]),
			.NE(gen[7972]),

			.O(gen[8065]),
			.E(gen[8067]),

			.SO(gen[8160]),
			.S(gen[8161]),
			.SE(gen[8162]),

			.SELF(gen[8066]),
			.cell_state(gen[8066])
		); 

/******************* CELL 8067 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8067 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7971]),
			.N(gen[7972]),
			.NE(gen[7973]),

			.O(gen[8066]),
			.E(gen[8068]),

			.SO(gen[8161]),
			.S(gen[8162]),
			.SE(gen[8163]),

			.SELF(gen[8067]),
			.cell_state(gen[8067])
		); 

/******************* CELL 8068 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8068 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7972]),
			.N(gen[7973]),
			.NE(gen[7974]),

			.O(gen[8067]),
			.E(gen[8069]),

			.SO(gen[8162]),
			.S(gen[8163]),
			.SE(gen[8164]),

			.SELF(gen[8068]),
			.cell_state(gen[8068])
		); 

/******************* CELL 8069 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8069 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7973]),
			.N(gen[7974]),
			.NE(gen[7975]),

			.O(gen[8068]),
			.E(gen[8070]),

			.SO(gen[8163]),
			.S(gen[8164]),
			.SE(gen[8165]),

			.SELF(gen[8069]),
			.cell_state(gen[8069])
		); 

/******************* CELL 8070 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8070 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7974]),
			.N(gen[7975]),
			.NE(gen[7976]),

			.O(gen[8069]),
			.E(gen[8071]),

			.SO(gen[8164]),
			.S(gen[8165]),
			.SE(gen[8166]),

			.SELF(gen[8070]),
			.cell_state(gen[8070])
		); 

/******************* CELL 8071 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8071 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7975]),
			.N(gen[7976]),
			.NE(gen[7977]),

			.O(gen[8070]),
			.E(gen[8072]),

			.SO(gen[8165]),
			.S(gen[8166]),
			.SE(gen[8167]),

			.SELF(gen[8071]),
			.cell_state(gen[8071])
		); 

/******************* CELL 8072 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8072 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7976]),
			.N(gen[7977]),
			.NE(gen[7978]),

			.O(gen[8071]),
			.E(gen[8073]),

			.SO(gen[8166]),
			.S(gen[8167]),
			.SE(gen[8168]),

			.SELF(gen[8072]),
			.cell_state(gen[8072])
		); 

/******************* CELL 8073 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8073 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7977]),
			.N(gen[7978]),
			.NE(gen[7979]),

			.O(gen[8072]),
			.E(gen[8074]),

			.SO(gen[8167]),
			.S(gen[8168]),
			.SE(gen[8169]),

			.SELF(gen[8073]),
			.cell_state(gen[8073])
		); 

/******************* CELL 8074 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8074 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7978]),
			.N(gen[7979]),
			.NE(gen[7978]),

			.O(gen[8073]),
			.E(gen[8073]),

			.SO(gen[8168]),
			.S(gen[8169]),
			.SE(gen[8168]),

			.SELF(gen[8074]),
			.cell_state(gen[8074])
		); 

/******************* CELL 8075 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8075 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7981]),
			.N(gen[7980]),
			.NE(gen[7981]),

			.O(gen[8076]),
			.E(gen[8076]),

			.SO(gen[8171]),
			.S(gen[8170]),
			.SE(gen[8171]),

			.SELF(gen[8075]),
			.cell_state(gen[8075])
		); 

/******************* CELL 8076 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8076 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7980]),
			.N(gen[7981]),
			.NE(gen[7982]),

			.O(gen[8075]),
			.E(gen[8077]),

			.SO(gen[8170]),
			.S(gen[8171]),
			.SE(gen[8172]),

			.SELF(gen[8076]),
			.cell_state(gen[8076])
		); 

/******************* CELL 8077 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8077 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7981]),
			.N(gen[7982]),
			.NE(gen[7983]),

			.O(gen[8076]),
			.E(gen[8078]),

			.SO(gen[8171]),
			.S(gen[8172]),
			.SE(gen[8173]),

			.SELF(gen[8077]),
			.cell_state(gen[8077])
		); 

/******************* CELL 8078 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8078 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7982]),
			.N(gen[7983]),
			.NE(gen[7984]),

			.O(gen[8077]),
			.E(gen[8079]),

			.SO(gen[8172]),
			.S(gen[8173]),
			.SE(gen[8174]),

			.SELF(gen[8078]),
			.cell_state(gen[8078])
		); 

/******************* CELL 8079 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8079 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7983]),
			.N(gen[7984]),
			.NE(gen[7985]),

			.O(gen[8078]),
			.E(gen[8080]),

			.SO(gen[8173]),
			.S(gen[8174]),
			.SE(gen[8175]),

			.SELF(gen[8079]),
			.cell_state(gen[8079])
		); 

/******************* CELL 8080 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8080 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7984]),
			.N(gen[7985]),
			.NE(gen[7986]),

			.O(gen[8079]),
			.E(gen[8081]),

			.SO(gen[8174]),
			.S(gen[8175]),
			.SE(gen[8176]),

			.SELF(gen[8080]),
			.cell_state(gen[8080])
		); 

/******************* CELL 8081 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8081 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7985]),
			.N(gen[7986]),
			.NE(gen[7987]),

			.O(gen[8080]),
			.E(gen[8082]),

			.SO(gen[8175]),
			.S(gen[8176]),
			.SE(gen[8177]),

			.SELF(gen[8081]),
			.cell_state(gen[8081])
		); 

/******************* CELL 8082 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8082 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7986]),
			.N(gen[7987]),
			.NE(gen[7988]),

			.O(gen[8081]),
			.E(gen[8083]),

			.SO(gen[8176]),
			.S(gen[8177]),
			.SE(gen[8178]),

			.SELF(gen[8082]),
			.cell_state(gen[8082])
		); 

/******************* CELL 8083 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8083 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7987]),
			.N(gen[7988]),
			.NE(gen[7989]),

			.O(gen[8082]),
			.E(gen[8084]),

			.SO(gen[8177]),
			.S(gen[8178]),
			.SE(gen[8179]),

			.SELF(gen[8083]),
			.cell_state(gen[8083])
		); 

/******************* CELL 8084 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8084 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7988]),
			.N(gen[7989]),
			.NE(gen[7990]),

			.O(gen[8083]),
			.E(gen[8085]),

			.SO(gen[8178]),
			.S(gen[8179]),
			.SE(gen[8180]),

			.SELF(gen[8084]),
			.cell_state(gen[8084])
		); 

/******************* CELL 8085 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8085 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7989]),
			.N(gen[7990]),
			.NE(gen[7991]),

			.O(gen[8084]),
			.E(gen[8086]),

			.SO(gen[8179]),
			.S(gen[8180]),
			.SE(gen[8181]),

			.SELF(gen[8085]),
			.cell_state(gen[8085])
		); 

/******************* CELL 8086 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8086 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7990]),
			.N(gen[7991]),
			.NE(gen[7992]),

			.O(gen[8085]),
			.E(gen[8087]),

			.SO(gen[8180]),
			.S(gen[8181]),
			.SE(gen[8182]),

			.SELF(gen[8086]),
			.cell_state(gen[8086])
		); 

/******************* CELL 8087 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8087 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7991]),
			.N(gen[7992]),
			.NE(gen[7993]),

			.O(gen[8086]),
			.E(gen[8088]),

			.SO(gen[8181]),
			.S(gen[8182]),
			.SE(gen[8183]),

			.SELF(gen[8087]),
			.cell_state(gen[8087])
		); 

/******************* CELL 8088 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8088 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7992]),
			.N(gen[7993]),
			.NE(gen[7994]),

			.O(gen[8087]),
			.E(gen[8089]),

			.SO(gen[8182]),
			.S(gen[8183]),
			.SE(gen[8184]),

			.SELF(gen[8088]),
			.cell_state(gen[8088])
		); 

/******************* CELL 8089 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8089 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7993]),
			.N(gen[7994]),
			.NE(gen[7995]),

			.O(gen[8088]),
			.E(gen[8090]),

			.SO(gen[8183]),
			.S(gen[8184]),
			.SE(gen[8185]),

			.SELF(gen[8089]),
			.cell_state(gen[8089])
		); 

/******************* CELL 8090 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8090 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7994]),
			.N(gen[7995]),
			.NE(gen[7996]),

			.O(gen[8089]),
			.E(gen[8091]),

			.SO(gen[8184]),
			.S(gen[8185]),
			.SE(gen[8186]),

			.SELF(gen[8090]),
			.cell_state(gen[8090])
		); 

/******************* CELL 8091 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8091 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7995]),
			.N(gen[7996]),
			.NE(gen[7997]),

			.O(gen[8090]),
			.E(gen[8092]),

			.SO(gen[8185]),
			.S(gen[8186]),
			.SE(gen[8187]),

			.SELF(gen[8091]),
			.cell_state(gen[8091])
		); 

/******************* CELL 8092 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8092 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7996]),
			.N(gen[7997]),
			.NE(gen[7998]),

			.O(gen[8091]),
			.E(gen[8093]),

			.SO(gen[8186]),
			.S(gen[8187]),
			.SE(gen[8188]),

			.SELF(gen[8092]),
			.cell_state(gen[8092])
		); 

/******************* CELL 8093 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8093 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7997]),
			.N(gen[7998]),
			.NE(gen[7999]),

			.O(gen[8092]),
			.E(gen[8094]),

			.SO(gen[8187]),
			.S(gen[8188]),
			.SE(gen[8189]),

			.SELF(gen[8093]),
			.cell_state(gen[8093])
		); 

/******************* CELL 8094 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8094 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7998]),
			.N(gen[7999]),
			.NE(gen[8000]),

			.O(gen[8093]),
			.E(gen[8095]),

			.SO(gen[8188]),
			.S(gen[8189]),
			.SE(gen[8190]),

			.SELF(gen[8094]),
			.cell_state(gen[8094])
		); 

/******************* CELL 8095 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8095 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7999]),
			.N(gen[8000]),
			.NE(gen[8001]),

			.O(gen[8094]),
			.E(gen[8096]),

			.SO(gen[8189]),
			.S(gen[8190]),
			.SE(gen[8191]),

			.SELF(gen[8095]),
			.cell_state(gen[8095])
		); 

/******************* CELL 8096 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8096 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8000]),
			.N(gen[8001]),
			.NE(gen[8002]),

			.O(gen[8095]),
			.E(gen[8097]),

			.SO(gen[8190]),
			.S(gen[8191]),
			.SE(gen[8192]),

			.SELF(gen[8096]),
			.cell_state(gen[8096])
		); 

/******************* CELL 8097 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8097 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8001]),
			.N(gen[8002]),
			.NE(gen[8003]),

			.O(gen[8096]),
			.E(gen[8098]),

			.SO(gen[8191]),
			.S(gen[8192]),
			.SE(gen[8193]),

			.SELF(gen[8097]),
			.cell_state(gen[8097])
		); 

/******************* CELL 8098 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8098 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8002]),
			.N(gen[8003]),
			.NE(gen[8004]),

			.O(gen[8097]),
			.E(gen[8099]),

			.SO(gen[8192]),
			.S(gen[8193]),
			.SE(gen[8194]),

			.SELF(gen[8098]),
			.cell_state(gen[8098])
		); 

/******************* CELL 8099 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8099 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8003]),
			.N(gen[8004]),
			.NE(gen[8005]),

			.O(gen[8098]),
			.E(gen[8100]),

			.SO(gen[8193]),
			.S(gen[8194]),
			.SE(gen[8195]),

			.SELF(gen[8099]),
			.cell_state(gen[8099])
		); 

/******************* CELL 8100 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8100 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8004]),
			.N(gen[8005]),
			.NE(gen[8006]),

			.O(gen[8099]),
			.E(gen[8101]),

			.SO(gen[8194]),
			.S(gen[8195]),
			.SE(gen[8196]),

			.SELF(gen[8100]),
			.cell_state(gen[8100])
		); 

/******************* CELL 8101 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8101 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8005]),
			.N(gen[8006]),
			.NE(gen[8007]),

			.O(gen[8100]),
			.E(gen[8102]),

			.SO(gen[8195]),
			.S(gen[8196]),
			.SE(gen[8197]),

			.SELF(gen[8101]),
			.cell_state(gen[8101])
		); 

/******************* CELL 8102 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8102 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8006]),
			.N(gen[8007]),
			.NE(gen[8008]),

			.O(gen[8101]),
			.E(gen[8103]),

			.SO(gen[8196]),
			.S(gen[8197]),
			.SE(gen[8198]),

			.SELF(gen[8102]),
			.cell_state(gen[8102])
		); 

/******************* CELL 8103 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8103 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8007]),
			.N(gen[8008]),
			.NE(gen[8009]),

			.O(gen[8102]),
			.E(gen[8104]),

			.SO(gen[8197]),
			.S(gen[8198]),
			.SE(gen[8199]),

			.SELF(gen[8103]),
			.cell_state(gen[8103])
		); 

/******************* CELL 8104 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8104 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8008]),
			.N(gen[8009]),
			.NE(gen[8010]),

			.O(gen[8103]),
			.E(gen[8105]),

			.SO(gen[8198]),
			.S(gen[8199]),
			.SE(gen[8200]),

			.SELF(gen[8104]),
			.cell_state(gen[8104])
		); 

/******************* CELL 8105 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8105 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8009]),
			.N(gen[8010]),
			.NE(gen[8011]),

			.O(gen[8104]),
			.E(gen[8106]),

			.SO(gen[8199]),
			.S(gen[8200]),
			.SE(gen[8201]),

			.SELF(gen[8105]),
			.cell_state(gen[8105])
		); 

/******************* CELL 8106 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8106 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8010]),
			.N(gen[8011]),
			.NE(gen[8012]),

			.O(gen[8105]),
			.E(gen[8107]),

			.SO(gen[8200]),
			.S(gen[8201]),
			.SE(gen[8202]),

			.SELF(gen[8106]),
			.cell_state(gen[8106])
		); 

/******************* CELL 8107 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8107 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8011]),
			.N(gen[8012]),
			.NE(gen[8013]),

			.O(gen[8106]),
			.E(gen[8108]),

			.SO(gen[8201]),
			.S(gen[8202]),
			.SE(gen[8203]),

			.SELF(gen[8107]),
			.cell_state(gen[8107])
		); 

/******************* CELL 8108 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8108 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8012]),
			.N(gen[8013]),
			.NE(gen[8014]),

			.O(gen[8107]),
			.E(gen[8109]),

			.SO(gen[8202]),
			.S(gen[8203]),
			.SE(gen[8204]),

			.SELF(gen[8108]),
			.cell_state(gen[8108])
		); 

/******************* CELL 8109 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8109 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8013]),
			.N(gen[8014]),
			.NE(gen[8015]),

			.O(gen[8108]),
			.E(gen[8110]),

			.SO(gen[8203]),
			.S(gen[8204]),
			.SE(gen[8205]),

			.SELF(gen[8109]),
			.cell_state(gen[8109])
		); 

/******************* CELL 8110 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8110 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8014]),
			.N(gen[8015]),
			.NE(gen[8016]),

			.O(gen[8109]),
			.E(gen[8111]),

			.SO(gen[8204]),
			.S(gen[8205]),
			.SE(gen[8206]),

			.SELF(gen[8110]),
			.cell_state(gen[8110])
		); 

/******************* CELL 8111 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8111 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8015]),
			.N(gen[8016]),
			.NE(gen[8017]),

			.O(gen[8110]),
			.E(gen[8112]),

			.SO(gen[8205]),
			.S(gen[8206]),
			.SE(gen[8207]),

			.SELF(gen[8111]),
			.cell_state(gen[8111])
		); 

/******************* CELL 8112 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8112 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8016]),
			.N(gen[8017]),
			.NE(gen[8018]),

			.O(gen[8111]),
			.E(gen[8113]),

			.SO(gen[8206]),
			.S(gen[8207]),
			.SE(gen[8208]),

			.SELF(gen[8112]),
			.cell_state(gen[8112])
		); 

/******************* CELL 8113 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8113 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8017]),
			.N(gen[8018]),
			.NE(gen[8019]),

			.O(gen[8112]),
			.E(gen[8114]),

			.SO(gen[8207]),
			.S(gen[8208]),
			.SE(gen[8209]),

			.SELF(gen[8113]),
			.cell_state(gen[8113])
		); 

/******************* CELL 8114 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8114 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8018]),
			.N(gen[8019]),
			.NE(gen[8020]),

			.O(gen[8113]),
			.E(gen[8115]),

			.SO(gen[8208]),
			.S(gen[8209]),
			.SE(gen[8210]),

			.SELF(gen[8114]),
			.cell_state(gen[8114])
		); 

/******************* CELL 8115 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8115 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8019]),
			.N(gen[8020]),
			.NE(gen[8021]),

			.O(gen[8114]),
			.E(gen[8116]),

			.SO(gen[8209]),
			.S(gen[8210]),
			.SE(gen[8211]),

			.SELF(gen[8115]),
			.cell_state(gen[8115])
		); 

/******************* CELL 8116 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8116 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8020]),
			.N(gen[8021]),
			.NE(gen[8022]),

			.O(gen[8115]),
			.E(gen[8117]),

			.SO(gen[8210]),
			.S(gen[8211]),
			.SE(gen[8212]),

			.SELF(gen[8116]),
			.cell_state(gen[8116])
		); 

/******************* CELL 8117 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8117 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8021]),
			.N(gen[8022]),
			.NE(gen[8023]),

			.O(gen[8116]),
			.E(gen[8118]),

			.SO(gen[8211]),
			.S(gen[8212]),
			.SE(gen[8213]),

			.SELF(gen[8117]),
			.cell_state(gen[8117])
		); 

/******************* CELL 8118 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8118 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8022]),
			.N(gen[8023]),
			.NE(gen[8024]),

			.O(gen[8117]),
			.E(gen[8119]),

			.SO(gen[8212]),
			.S(gen[8213]),
			.SE(gen[8214]),

			.SELF(gen[8118]),
			.cell_state(gen[8118])
		); 

/******************* CELL 8119 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8119 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8023]),
			.N(gen[8024]),
			.NE(gen[8025]),

			.O(gen[8118]),
			.E(gen[8120]),

			.SO(gen[8213]),
			.S(gen[8214]),
			.SE(gen[8215]),

			.SELF(gen[8119]),
			.cell_state(gen[8119])
		); 

/******************* CELL 8120 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8120 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8024]),
			.N(gen[8025]),
			.NE(gen[8026]),

			.O(gen[8119]),
			.E(gen[8121]),

			.SO(gen[8214]),
			.S(gen[8215]),
			.SE(gen[8216]),

			.SELF(gen[8120]),
			.cell_state(gen[8120])
		); 

/******************* CELL 8121 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8121 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8025]),
			.N(gen[8026]),
			.NE(gen[8027]),

			.O(gen[8120]),
			.E(gen[8122]),

			.SO(gen[8215]),
			.S(gen[8216]),
			.SE(gen[8217]),

			.SELF(gen[8121]),
			.cell_state(gen[8121])
		); 

/******************* CELL 8122 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8122 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8026]),
			.N(gen[8027]),
			.NE(gen[8028]),

			.O(gen[8121]),
			.E(gen[8123]),

			.SO(gen[8216]),
			.S(gen[8217]),
			.SE(gen[8218]),

			.SELF(gen[8122]),
			.cell_state(gen[8122])
		); 

/******************* CELL 8123 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8123 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8027]),
			.N(gen[8028]),
			.NE(gen[8029]),

			.O(gen[8122]),
			.E(gen[8124]),

			.SO(gen[8217]),
			.S(gen[8218]),
			.SE(gen[8219]),

			.SELF(gen[8123]),
			.cell_state(gen[8123])
		); 

/******************* CELL 8124 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8124 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8028]),
			.N(gen[8029]),
			.NE(gen[8030]),

			.O(gen[8123]),
			.E(gen[8125]),

			.SO(gen[8218]),
			.S(gen[8219]),
			.SE(gen[8220]),

			.SELF(gen[8124]),
			.cell_state(gen[8124])
		); 

/******************* CELL 8125 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8125 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8029]),
			.N(gen[8030]),
			.NE(gen[8031]),

			.O(gen[8124]),
			.E(gen[8126]),

			.SO(gen[8219]),
			.S(gen[8220]),
			.SE(gen[8221]),

			.SELF(gen[8125]),
			.cell_state(gen[8125])
		); 

/******************* CELL 8126 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8126 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8030]),
			.N(gen[8031]),
			.NE(gen[8032]),

			.O(gen[8125]),
			.E(gen[8127]),

			.SO(gen[8220]),
			.S(gen[8221]),
			.SE(gen[8222]),

			.SELF(gen[8126]),
			.cell_state(gen[8126])
		); 

/******************* CELL 8127 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8127 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8031]),
			.N(gen[8032]),
			.NE(gen[8033]),

			.O(gen[8126]),
			.E(gen[8128]),

			.SO(gen[8221]),
			.S(gen[8222]),
			.SE(gen[8223]),

			.SELF(gen[8127]),
			.cell_state(gen[8127])
		); 

/******************* CELL 8128 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8128 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8032]),
			.N(gen[8033]),
			.NE(gen[8034]),

			.O(gen[8127]),
			.E(gen[8129]),

			.SO(gen[8222]),
			.S(gen[8223]),
			.SE(gen[8224]),

			.SELF(gen[8128]),
			.cell_state(gen[8128])
		); 

/******************* CELL 8129 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8129 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8033]),
			.N(gen[8034]),
			.NE(gen[8035]),

			.O(gen[8128]),
			.E(gen[8130]),

			.SO(gen[8223]),
			.S(gen[8224]),
			.SE(gen[8225]),

			.SELF(gen[8129]),
			.cell_state(gen[8129])
		); 

/******************* CELL 8130 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8130 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8034]),
			.N(gen[8035]),
			.NE(gen[8036]),

			.O(gen[8129]),
			.E(gen[8131]),

			.SO(gen[8224]),
			.S(gen[8225]),
			.SE(gen[8226]),

			.SELF(gen[8130]),
			.cell_state(gen[8130])
		); 

/******************* CELL 8131 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8131 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8035]),
			.N(gen[8036]),
			.NE(gen[8037]),

			.O(gen[8130]),
			.E(gen[8132]),

			.SO(gen[8225]),
			.S(gen[8226]),
			.SE(gen[8227]),

			.SELF(gen[8131]),
			.cell_state(gen[8131])
		); 

/******************* CELL 8132 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8132 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8036]),
			.N(gen[8037]),
			.NE(gen[8038]),

			.O(gen[8131]),
			.E(gen[8133]),

			.SO(gen[8226]),
			.S(gen[8227]),
			.SE(gen[8228]),

			.SELF(gen[8132]),
			.cell_state(gen[8132])
		); 

/******************* CELL 8133 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8133 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8037]),
			.N(gen[8038]),
			.NE(gen[8039]),

			.O(gen[8132]),
			.E(gen[8134]),

			.SO(gen[8227]),
			.S(gen[8228]),
			.SE(gen[8229]),

			.SELF(gen[8133]),
			.cell_state(gen[8133])
		); 

/******************* CELL 8134 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8134 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8038]),
			.N(gen[8039]),
			.NE(gen[8040]),

			.O(gen[8133]),
			.E(gen[8135]),

			.SO(gen[8228]),
			.S(gen[8229]),
			.SE(gen[8230]),

			.SELF(gen[8134]),
			.cell_state(gen[8134])
		); 

/******************* CELL 8135 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8135 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8039]),
			.N(gen[8040]),
			.NE(gen[8041]),

			.O(gen[8134]),
			.E(gen[8136]),

			.SO(gen[8229]),
			.S(gen[8230]),
			.SE(gen[8231]),

			.SELF(gen[8135]),
			.cell_state(gen[8135])
		); 

/******************* CELL 8136 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8136 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8040]),
			.N(gen[8041]),
			.NE(gen[8042]),

			.O(gen[8135]),
			.E(gen[8137]),

			.SO(gen[8230]),
			.S(gen[8231]),
			.SE(gen[8232]),

			.SELF(gen[8136]),
			.cell_state(gen[8136])
		); 

/******************* CELL 8137 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8137 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8041]),
			.N(gen[8042]),
			.NE(gen[8043]),

			.O(gen[8136]),
			.E(gen[8138]),

			.SO(gen[8231]),
			.S(gen[8232]),
			.SE(gen[8233]),

			.SELF(gen[8137]),
			.cell_state(gen[8137])
		); 

/******************* CELL 8138 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8138 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8042]),
			.N(gen[8043]),
			.NE(gen[8044]),

			.O(gen[8137]),
			.E(gen[8139]),

			.SO(gen[8232]),
			.S(gen[8233]),
			.SE(gen[8234]),

			.SELF(gen[8138]),
			.cell_state(gen[8138])
		); 

/******************* CELL 8139 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8139 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8043]),
			.N(gen[8044]),
			.NE(gen[8045]),

			.O(gen[8138]),
			.E(gen[8140]),

			.SO(gen[8233]),
			.S(gen[8234]),
			.SE(gen[8235]),

			.SELF(gen[8139]),
			.cell_state(gen[8139])
		); 

/******************* CELL 8140 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8140 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8044]),
			.N(gen[8045]),
			.NE(gen[8046]),

			.O(gen[8139]),
			.E(gen[8141]),

			.SO(gen[8234]),
			.S(gen[8235]),
			.SE(gen[8236]),

			.SELF(gen[8140]),
			.cell_state(gen[8140])
		); 

/******************* CELL 8141 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8141 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8045]),
			.N(gen[8046]),
			.NE(gen[8047]),

			.O(gen[8140]),
			.E(gen[8142]),

			.SO(gen[8235]),
			.S(gen[8236]),
			.SE(gen[8237]),

			.SELF(gen[8141]),
			.cell_state(gen[8141])
		); 

/******************* CELL 8142 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8142 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8046]),
			.N(gen[8047]),
			.NE(gen[8048]),

			.O(gen[8141]),
			.E(gen[8143]),

			.SO(gen[8236]),
			.S(gen[8237]),
			.SE(gen[8238]),

			.SELF(gen[8142]),
			.cell_state(gen[8142])
		); 

/******************* CELL 8143 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8143 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8047]),
			.N(gen[8048]),
			.NE(gen[8049]),

			.O(gen[8142]),
			.E(gen[8144]),

			.SO(gen[8237]),
			.S(gen[8238]),
			.SE(gen[8239]),

			.SELF(gen[8143]),
			.cell_state(gen[8143])
		); 

/******************* CELL 8144 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8144 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8048]),
			.N(gen[8049]),
			.NE(gen[8050]),

			.O(gen[8143]),
			.E(gen[8145]),

			.SO(gen[8238]),
			.S(gen[8239]),
			.SE(gen[8240]),

			.SELF(gen[8144]),
			.cell_state(gen[8144])
		); 

/******************* CELL 8145 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8145 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8049]),
			.N(gen[8050]),
			.NE(gen[8051]),

			.O(gen[8144]),
			.E(gen[8146]),

			.SO(gen[8239]),
			.S(gen[8240]),
			.SE(gen[8241]),

			.SELF(gen[8145]),
			.cell_state(gen[8145])
		); 

/******************* CELL 8146 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8146 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8050]),
			.N(gen[8051]),
			.NE(gen[8052]),

			.O(gen[8145]),
			.E(gen[8147]),

			.SO(gen[8240]),
			.S(gen[8241]),
			.SE(gen[8242]),

			.SELF(gen[8146]),
			.cell_state(gen[8146])
		); 

/******************* CELL 8147 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8147 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8051]),
			.N(gen[8052]),
			.NE(gen[8053]),

			.O(gen[8146]),
			.E(gen[8148]),

			.SO(gen[8241]),
			.S(gen[8242]),
			.SE(gen[8243]),

			.SELF(gen[8147]),
			.cell_state(gen[8147])
		); 

/******************* CELL 8148 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8148 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8052]),
			.N(gen[8053]),
			.NE(gen[8054]),

			.O(gen[8147]),
			.E(gen[8149]),

			.SO(gen[8242]),
			.S(gen[8243]),
			.SE(gen[8244]),

			.SELF(gen[8148]),
			.cell_state(gen[8148])
		); 

/******************* CELL 8149 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8149 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8053]),
			.N(gen[8054]),
			.NE(gen[8055]),

			.O(gen[8148]),
			.E(gen[8150]),

			.SO(gen[8243]),
			.S(gen[8244]),
			.SE(gen[8245]),

			.SELF(gen[8149]),
			.cell_state(gen[8149])
		); 

/******************* CELL 8150 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8150 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8054]),
			.N(gen[8055]),
			.NE(gen[8056]),

			.O(gen[8149]),
			.E(gen[8151]),

			.SO(gen[8244]),
			.S(gen[8245]),
			.SE(gen[8246]),

			.SELF(gen[8150]),
			.cell_state(gen[8150])
		); 

/******************* CELL 8151 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8151 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8055]),
			.N(gen[8056]),
			.NE(gen[8057]),

			.O(gen[8150]),
			.E(gen[8152]),

			.SO(gen[8245]),
			.S(gen[8246]),
			.SE(gen[8247]),

			.SELF(gen[8151]),
			.cell_state(gen[8151])
		); 

/******************* CELL 8152 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8152 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8056]),
			.N(gen[8057]),
			.NE(gen[8058]),

			.O(gen[8151]),
			.E(gen[8153]),

			.SO(gen[8246]),
			.S(gen[8247]),
			.SE(gen[8248]),

			.SELF(gen[8152]),
			.cell_state(gen[8152])
		); 

/******************* CELL 8153 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8153 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8057]),
			.N(gen[8058]),
			.NE(gen[8059]),

			.O(gen[8152]),
			.E(gen[8154]),

			.SO(gen[8247]),
			.S(gen[8248]),
			.SE(gen[8249]),

			.SELF(gen[8153]),
			.cell_state(gen[8153])
		); 

/******************* CELL 8154 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8154 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8058]),
			.N(gen[8059]),
			.NE(gen[8060]),

			.O(gen[8153]),
			.E(gen[8155]),

			.SO(gen[8248]),
			.S(gen[8249]),
			.SE(gen[8250]),

			.SELF(gen[8154]),
			.cell_state(gen[8154])
		); 

/******************* CELL 8155 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8155 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8059]),
			.N(gen[8060]),
			.NE(gen[8061]),

			.O(gen[8154]),
			.E(gen[8156]),

			.SO(gen[8249]),
			.S(gen[8250]),
			.SE(gen[8251]),

			.SELF(gen[8155]),
			.cell_state(gen[8155])
		); 

/******************* CELL 8156 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8156 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8060]),
			.N(gen[8061]),
			.NE(gen[8062]),

			.O(gen[8155]),
			.E(gen[8157]),

			.SO(gen[8250]),
			.S(gen[8251]),
			.SE(gen[8252]),

			.SELF(gen[8156]),
			.cell_state(gen[8156])
		); 

/******************* CELL 8157 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8157 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8061]),
			.N(gen[8062]),
			.NE(gen[8063]),

			.O(gen[8156]),
			.E(gen[8158]),

			.SO(gen[8251]),
			.S(gen[8252]),
			.SE(gen[8253]),

			.SELF(gen[8157]),
			.cell_state(gen[8157])
		); 

/******************* CELL 8158 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8158 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8062]),
			.N(gen[8063]),
			.NE(gen[8064]),

			.O(gen[8157]),
			.E(gen[8159]),

			.SO(gen[8252]),
			.S(gen[8253]),
			.SE(gen[8254]),

			.SELF(gen[8158]),
			.cell_state(gen[8158])
		); 

/******************* CELL 8159 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8159 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8063]),
			.N(gen[8064]),
			.NE(gen[8065]),

			.O(gen[8158]),
			.E(gen[8160]),

			.SO(gen[8253]),
			.S(gen[8254]),
			.SE(gen[8255]),

			.SELF(gen[8159]),
			.cell_state(gen[8159])
		); 

/******************* CELL 8160 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8160 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8064]),
			.N(gen[8065]),
			.NE(gen[8066]),

			.O(gen[8159]),
			.E(gen[8161]),

			.SO(gen[8254]),
			.S(gen[8255]),
			.SE(gen[8256]),

			.SELF(gen[8160]),
			.cell_state(gen[8160])
		); 

/******************* CELL 8161 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8161 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8065]),
			.N(gen[8066]),
			.NE(gen[8067]),

			.O(gen[8160]),
			.E(gen[8162]),

			.SO(gen[8255]),
			.S(gen[8256]),
			.SE(gen[8257]),

			.SELF(gen[8161]),
			.cell_state(gen[8161])
		); 

/******************* CELL 8162 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8162 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8066]),
			.N(gen[8067]),
			.NE(gen[8068]),

			.O(gen[8161]),
			.E(gen[8163]),

			.SO(gen[8256]),
			.S(gen[8257]),
			.SE(gen[8258]),

			.SELF(gen[8162]),
			.cell_state(gen[8162])
		); 

/******************* CELL 8163 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8163 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8067]),
			.N(gen[8068]),
			.NE(gen[8069]),

			.O(gen[8162]),
			.E(gen[8164]),

			.SO(gen[8257]),
			.S(gen[8258]),
			.SE(gen[8259]),

			.SELF(gen[8163]),
			.cell_state(gen[8163])
		); 

/******************* CELL 8164 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8164 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8068]),
			.N(gen[8069]),
			.NE(gen[8070]),

			.O(gen[8163]),
			.E(gen[8165]),

			.SO(gen[8258]),
			.S(gen[8259]),
			.SE(gen[8260]),

			.SELF(gen[8164]),
			.cell_state(gen[8164])
		); 

/******************* CELL 8165 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8165 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8069]),
			.N(gen[8070]),
			.NE(gen[8071]),

			.O(gen[8164]),
			.E(gen[8166]),

			.SO(gen[8259]),
			.S(gen[8260]),
			.SE(gen[8261]),

			.SELF(gen[8165]),
			.cell_state(gen[8165])
		); 

/******************* CELL 8166 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8166 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8070]),
			.N(gen[8071]),
			.NE(gen[8072]),

			.O(gen[8165]),
			.E(gen[8167]),

			.SO(gen[8260]),
			.S(gen[8261]),
			.SE(gen[8262]),

			.SELF(gen[8166]),
			.cell_state(gen[8166])
		); 

/******************* CELL 8167 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8167 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8071]),
			.N(gen[8072]),
			.NE(gen[8073]),

			.O(gen[8166]),
			.E(gen[8168]),

			.SO(gen[8261]),
			.S(gen[8262]),
			.SE(gen[8263]),

			.SELF(gen[8167]),
			.cell_state(gen[8167])
		); 

/******************* CELL 8168 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8168 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8072]),
			.N(gen[8073]),
			.NE(gen[8074]),

			.O(gen[8167]),
			.E(gen[8169]),

			.SO(gen[8262]),
			.S(gen[8263]),
			.SE(gen[8264]),

			.SELF(gen[8168]),
			.cell_state(gen[8168])
		); 

/******************* CELL 8169 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8169 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8073]),
			.N(gen[8074]),
			.NE(gen[8073]),

			.O(gen[8168]),
			.E(gen[8168]),

			.SO(gen[8263]),
			.S(gen[8264]),
			.SE(gen[8263]),

			.SELF(gen[8169]),
			.cell_state(gen[8169])
		); 

/******************* CELL 8170 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8170 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8076]),
			.N(gen[8075]),
			.NE(gen[8076]),

			.O(gen[8171]),
			.E(gen[8171]),

			.SO(gen[8266]),
			.S(gen[8265]),
			.SE(gen[8266]),

			.SELF(gen[8170]),
			.cell_state(gen[8170])
		); 

/******************* CELL 8171 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8171 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8075]),
			.N(gen[8076]),
			.NE(gen[8077]),

			.O(gen[8170]),
			.E(gen[8172]),

			.SO(gen[8265]),
			.S(gen[8266]),
			.SE(gen[8267]),

			.SELF(gen[8171]),
			.cell_state(gen[8171])
		); 

/******************* CELL 8172 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8172 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8076]),
			.N(gen[8077]),
			.NE(gen[8078]),

			.O(gen[8171]),
			.E(gen[8173]),

			.SO(gen[8266]),
			.S(gen[8267]),
			.SE(gen[8268]),

			.SELF(gen[8172]),
			.cell_state(gen[8172])
		); 

/******************* CELL 8173 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8173 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8077]),
			.N(gen[8078]),
			.NE(gen[8079]),

			.O(gen[8172]),
			.E(gen[8174]),

			.SO(gen[8267]),
			.S(gen[8268]),
			.SE(gen[8269]),

			.SELF(gen[8173]),
			.cell_state(gen[8173])
		); 

/******************* CELL 8174 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8174 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8078]),
			.N(gen[8079]),
			.NE(gen[8080]),

			.O(gen[8173]),
			.E(gen[8175]),

			.SO(gen[8268]),
			.S(gen[8269]),
			.SE(gen[8270]),

			.SELF(gen[8174]),
			.cell_state(gen[8174])
		); 

/******************* CELL 8175 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8175 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8079]),
			.N(gen[8080]),
			.NE(gen[8081]),

			.O(gen[8174]),
			.E(gen[8176]),

			.SO(gen[8269]),
			.S(gen[8270]),
			.SE(gen[8271]),

			.SELF(gen[8175]),
			.cell_state(gen[8175])
		); 

/******************* CELL 8176 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8176 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8080]),
			.N(gen[8081]),
			.NE(gen[8082]),

			.O(gen[8175]),
			.E(gen[8177]),

			.SO(gen[8270]),
			.S(gen[8271]),
			.SE(gen[8272]),

			.SELF(gen[8176]),
			.cell_state(gen[8176])
		); 

/******************* CELL 8177 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8177 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8081]),
			.N(gen[8082]),
			.NE(gen[8083]),

			.O(gen[8176]),
			.E(gen[8178]),

			.SO(gen[8271]),
			.S(gen[8272]),
			.SE(gen[8273]),

			.SELF(gen[8177]),
			.cell_state(gen[8177])
		); 

/******************* CELL 8178 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8178 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8082]),
			.N(gen[8083]),
			.NE(gen[8084]),

			.O(gen[8177]),
			.E(gen[8179]),

			.SO(gen[8272]),
			.S(gen[8273]),
			.SE(gen[8274]),

			.SELF(gen[8178]),
			.cell_state(gen[8178])
		); 

/******************* CELL 8179 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8179 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8083]),
			.N(gen[8084]),
			.NE(gen[8085]),

			.O(gen[8178]),
			.E(gen[8180]),

			.SO(gen[8273]),
			.S(gen[8274]),
			.SE(gen[8275]),

			.SELF(gen[8179]),
			.cell_state(gen[8179])
		); 

/******************* CELL 8180 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8180 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8084]),
			.N(gen[8085]),
			.NE(gen[8086]),

			.O(gen[8179]),
			.E(gen[8181]),

			.SO(gen[8274]),
			.S(gen[8275]),
			.SE(gen[8276]),

			.SELF(gen[8180]),
			.cell_state(gen[8180])
		); 

/******************* CELL 8181 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8181 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8085]),
			.N(gen[8086]),
			.NE(gen[8087]),

			.O(gen[8180]),
			.E(gen[8182]),

			.SO(gen[8275]),
			.S(gen[8276]),
			.SE(gen[8277]),

			.SELF(gen[8181]),
			.cell_state(gen[8181])
		); 

/******************* CELL 8182 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8182 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8086]),
			.N(gen[8087]),
			.NE(gen[8088]),

			.O(gen[8181]),
			.E(gen[8183]),

			.SO(gen[8276]),
			.S(gen[8277]),
			.SE(gen[8278]),

			.SELF(gen[8182]),
			.cell_state(gen[8182])
		); 

/******************* CELL 8183 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8183 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8087]),
			.N(gen[8088]),
			.NE(gen[8089]),

			.O(gen[8182]),
			.E(gen[8184]),

			.SO(gen[8277]),
			.S(gen[8278]),
			.SE(gen[8279]),

			.SELF(gen[8183]),
			.cell_state(gen[8183])
		); 

/******************* CELL 8184 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8184 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8088]),
			.N(gen[8089]),
			.NE(gen[8090]),

			.O(gen[8183]),
			.E(gen[8185]),

			.SO(gen[8278]),
			.S(gen[8279]),
			.SE(gen[8280]),

			.SELF(gen[8184]),
			.cell_state(gen[8184])
		); 

/******************* CELL 8185 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8185 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8089]),
			.N(gen[8090]),
			.NE(gen[8091]),

			.O(gen[8184]),
			.E(gen[8186]),

			.SO(gen[8279]),
			.S(gen[8280]),
			.SE(gen[8281]),

			.SELF(gen[8185]),
			.cell_state(gen[8185])
		); 

/******************* CELL 8186 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8186 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8090]),
			.N(gen[8091]),
			.NE(gen[8092]),

			.O(gen[8185]),
			.E(gen[8187]),

			.SO(gen[8280]),
			.S(gen[8281]),
			.SE(gen[8282]),

			.SELF(gen[8186]),
			.cell_state(gen[8186])
		); 

/******************* CELL 8187 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8187 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8091]),
			.N(gen[8092]),
			.NE(gen[8093]),

			.O(gen[8186]),
			.E(gen[8188]),

			.SO(gen[8281]),
			.S(gen[8282]),
			.SE(gen[8283]),

			.SELF(gen[8187]),
			.cell_state(gen[8187])
		); 

/******************* CELL 8188 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8188 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8092]),
			.N(gen[8093]),
			.NE(gen[8094]),

			.O(gen[8187]),
			.E(gen[8189]),

			.SO(gen[8282]),
			.S(gen[8283]),
			.SE(gen[8284]),

			.SELF(gen[8188]),
			.cell_state(gen[8188])
		); 

/******************* CELL 8189 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8189 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8093]),
			.N(gen[8094]),
			.NE(gen[8095]),

			.O(gen[8188]),
			.E(gen[8190]),

			.SO(gen[8283]),
			.S(gen[8284]),
			.SE(gen[8285]),

			.SELF(gen[8189]),
			.cell_state(gen[8189])
		); 

/******************* CELL 8190 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8190 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8094]),
			.N(gen[8095]),
			.NE(gen[8096]),

			.O(gen[8189]),
			.E(gen[8191]),

			.SO(gen[8284]),
			.S(gen[8285]),
			.SE(gen[8286]),

			.SELF(gen[8190]),
			.cell_state(gen[8190])
		); 

/******************* CELL 8191 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8191 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8095]),
			.N(gen[8096]),
			.NE(gen[8097]),

			.O(gen[8190]),
			.E(gen[8192]),

			.SO(gen[8285]),
			.S(gen[8286]),
			.SE(gen[8287]),

			.SELF(gen[8191]),
			.cell_state(gen[8191])
		); 

/******************* CELL 8192 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8192 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8096]),
			.N(gen[8097]),
			.NE(gen[8098]),

			.O(gen[8191]),
			.E(gen[8193]),

			.SO(gen[8286]),
			.S(gen[8287]),
			.SE(gen[8288]),

			.SELF(gen[8192]),
			.cell_state(gen[8192])
		); 

/******************* CELL 8193 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8193 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8097]),
			.N(gen[8098]),
			.NE(gen[8099]),

			.O(gen[8192]),
			.E(gen[8194]),

			.SO(gen[8287]),
			.S(gen[8288]),
			.SE(gen[8289]),

			.SELF(gen[8193]),
			.cell_state(gen[8193])
		); 

/******************* CELL 8194 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8194 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8098]),
			.N(gen[8099]),
			.NE(gen[8100]),

			.O(gen[8193]),
			.E(gen[8195]),

			.SO(gen[8288]),
			.S(gen[8289]),
			.SE(gen[8290]),

			.SELF(gen[8194]),
			.cell_state(gen[8194])
		); 

/******************* CELL 8195 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8195 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8099]),
			.N(gen[8100]),
			.NE(gen[8101]),

			.O(gen[8194]),
			.E(gen[8196]),

			.SO(gen[8289]),
			.S(gen[8290]),
			.SE(gen[8291]),

			.SELF(gen[8195]),
			.cell_state(gen[8195])
		); 

/******************* CELL 8196 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8196 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8100]),
			.N(gen[8101]),
			.NE(gen[8102]),

			.O(gen[8195]),
			.E(gen[8197]),

			.SO(gen[8290]),
			.S(gen[8291]),
			.SE(gen[8292]),

			.SELF(gen[8196]),
			.cell_state(gen[8196])
		); 

/******************* CELL 8197 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8197 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8101]),
			.N(gen[8102]),
			.NE(gen[8103]),

			.O(gen[8196]),
			.E(gen[8198]),

			.SO(gen[8291]),
			.S(gen[8292]),
			.SE(gen[8293]),

			.SELF(gen[8197]),
			.cell_state(gen[8197])
		); 

/******************* CELL 8198 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8198 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8102]),
			.N(gen[8103]),
			.NE(gen[8104]),

			.O(gen[8197]),
			.E(gen[8199]),

			.SO(gen[8292]),
			.S(gen[8293]),
			.SE(gen[8294]),

			.SELF(gen[8198]),
			.cell_state(gen[8198])
		); 

/******************* CELL 8199 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8199 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8103]),
			.N(gen[8104]),
			.NE(gen[8105]),

			.O(gen[8198]),
			.E(gen[8200]),

			.SO(gen[8293]),
			.S(gen[8294]),
			.SE(gen[8295]),

			.SELF(gen[8199]),
			.cell_state(gen[8199])
		); 

/******************* CELL 8200 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8200 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8104]),
			.N(gen[8105]),
			.NE(gen[8106]),

			.O(gen[8199]),
			.E(gen[8201]),

			.SO(gen[8294]),
			.S(gen[8295]),
			.SE(gen[8296]),

			.SELF(gen[8200]),
			.cell_state(gen[8200])
		); 

/******************* CELL 8201 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8201 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8105]),
			.N(gen[8106]),
			.NE(gen[8107]),

			.O(gen[8200]),
			.E(gen[8202]),

			.SO(gen[8295]),
			.S(gen[8296]),
			.SE(gen[8297]),

			.SELF(gen[8201]),
			.cell_state(gen[8201])
		); 

/******************* CELL 8202 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8202 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8106]),
			.N(gen[8107]),
			.NE(gen[8108]),

			.O(gen[8201]),
			.E(gen[8203]),

			.SO(gen[8296]),
			.S(gen[8297]),
			.SE(gen[8298]),

			.SELF(gen[8202]),
			.cell_state(gen[8202])
		); 

/******************* CELL 8203 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8203 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8107]),
			.N(gen[8108]),
			.NE(gen[8109]),

			.O(gen[8202]),
			.E(gen[8204]),

			.SO(gen[8297]),
			.S(gen[8298]),
			.SE(gen[8299]),

			.SELF(gen[8203]),
			.cell_state(gen[8203])
		); 

/******************* CELL 8204 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8204 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8108]),
			.N(gen[8109]),
			.NE(gen[8110]),

			.O(gen[8203]),
			.E(gen[8205]),

			.SO(gen[8298]),
			.S(gen[8299]),
			.SE(gen[8300]),

			.SELF(gen[8204]),
			.cell_state(gen[8204])
		); 

/******************* CELL 8205 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8205 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8109]),
			.N(gen[8110]),
			.NE(gen[8111]),

			.O(gen[8204]),
			.E(gen[8206]),

			.SO(gen[8299]),
			.S(gen[8300]),
			.SE(gen[8301]),

			.SELF(gen[8205]),
			.cell_state(gen[8205])
		); 

/******************* CELL 8206 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8206 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8110]),
			.N(gen[8111]),
			.NE(gen[8112]),

			.O(gen[8205]),
			.E(gen[8207]),

			.SO(gen[8300]),
			.S(gen[8301]),
			.SE(gen[8302]),

			.SELF(gen[8206]),
			.cell_state(gen[8206])
		); 

/******************* CELL 8207 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8207 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8111]),
			.N(gen[8112]),
			.NE(gen[8113]),

			.O(gen[8206]),
			.E(gen[8208]),

			.SO(gen[8301]),
			.S(gen[8302]),
			.SE(gen[8303]),

			.SELF(gen[8207]),
			.cell_state(gen[8207])
		); 

/******************* CELL 8208 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8208 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8112]),
			.N(gen[8113]),
			.NE(gen[8114]),

			.O(gen[8207]),
			.E(gen[8209]),

			.SO(gen[8302]),
			.S(gen[8303]),
			.SE(gen[8304]),

			.SELF(gen[8208]),
			.cell_state(gen[8208])
		); 

/******************* CELL 8209 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8209 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8113]),
			.N(gen[8114]),
			.NE(gen[8115]),

			.O(gen[8208]),
			.E(gen[8210]),

			.SO(gen[8303]),
			.S(gen[8304]),
			.SE(gen[8305]),

			.SELF(gen[8209]),
			.cell_state(gen[8209])
		); 

/******************* CELL 8210 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8210 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8114]),
			.N(gen[8115]),
			.NE(gen[8116]),

			.O(gen[8209]),
			.E(gen[8211]),

			.SO(gen[8304]),
			.S(gen[8305]),
			.SE(gen[8306]),

			.SELF(gen[8210]),
			.cell_state(gen[8210])
		); 

/******************* CELL 8211 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8211 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8115]),
			.N(gen[8116]),
			.NE(gen[8117]),

			.O(gen[8210]),
			.E(gen[8212]),

			.SO(gen[8305]),
			.S(gen[8306]),
			.SE(gen[8307]),

			.SELF(gen[8211]),
			.cell_state(gen[8211])
		); 

/******************* CELL 8212 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8212 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8116]),
			.N(gen[8117]),
			.NE(gen[8118]),

			.O(gen[8211]),
			.E(gen[8213]),

			.SO(gen[8306]),
			.S(gen[8307]),
			.SE(gen[8308]),

			.SELF(gen[8212]),
			.cell_state(gen[8212])
		); 

/******************* CELL 8213 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8213 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8117]),
			.N(gen[8118]),
			.NE(gen[8119]),

			.O(gen[8212]),
			.E(gen[8214]),

			.SO(gen[8307]),
			.S(gen[8308]),
			.SE(gen[8309]),

			.SELF(gen[8213]),
			.cell_state(gen[8213])
		); 

/******************* CELL 8214 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8214 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8118]),
			.N(gen[8119]),
			.NE(gen[8120]),

			.O(gen[8213]),
			.E(gen[8215]),

			.SO(gen[8308]),
			.S(gen[8309]),
			.SE(gen[8310]),

			.SELF(gen[8214]),
			.cell_state(gen[8214])
		); 

/******************* CELL 8215 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8215 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8119]),
			.N(gen[8120]),
			.NE(gen[8121]),

			.O(gen[8214]),
			.E(gen[8216]),

			.SO(gen[8309]),
			.S(gen[8310]),
			.SE(gen[8311]),

			.SELF(gen[8215]),
			.cell_state(gen[8215])
		); 

/******************* CELL 8216 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8216 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8120]),
			.N(gen[8121]),
			.NE(gen[8122]),

			.O(gen[8215]),
			.E(gen[8217]),

			.SO(gen[8310]),
			.S(gen[8311]),
			.SE(gen[8312]),

			.SELF(gen[8216]),
			.cell_state(gen[8216])
		); 

/******************* CELL 8217 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8217 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8121]),
			.N(gen[8122]),
			.NE(gen[8123]),

			.O(gen[8216]),
			.E(gen[8218]),

			.SO(gen[8311]),
			.S(gen[8312]),
			.SE(gen[8313]),

			.SELF(gen[8217]),
			.cell_state(gen[8217])
		); 

/******************* CELL 8218 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8218 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8122]),
			.N(gen[8123]),
			.NE(gen[8124]),

			.O(gen[8217]),
			.E(gen[8219]),

			.SO(gen[8312]),
			.S(gen[8313]),
			.SE(gen[8314]),

			.SELF(gen[8218]),
			.cell_state(gen[8218])
		); 

/******************* CELL 8219 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8219 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8123]),
			.N(gen[8124]),
			.NE(gen[8125]),

			.O(gen[8218]),
			.E(gen[8220]),

			.SO(gen[8313]),
			.S(gen[8314]),
			.SE(gen[8315]),

			.SELF(gen[8219]),
			.cell_state(gen[8219])
		); 

/******************* CELL 8220 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8220 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8124]),
			.N(gen[8125]),
			.NE(gen[8126]),

			.O(gen[8219]),
			.E(gen[8221]),

			.SO(gen[8314]),
			.S(gen[8315]),
			.SE(gen[8316]),

			.SELF(gen[8220]),
			.cell_state(gen[8220])
		); 

/******************* CELL 8221 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8221 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8125]),
			.N(gen[8126]),
			.NE(gen[8127]),

			.O(gen[8220]),
			.E(gen[8222]),

			.SO(gen[8315]),
			.S(gen[8316]),
			.SE(gen[8317]),

			.SELF(gen[8221]),
			.cell_state(gen[8221])
		); 

/******************* CELL 8222 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8222 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8126]),
			.N(gen[8127]),
			.NE(gen[8128]),

			.O(gen[8221]),
			.E(gen[8223]),

			.SO(gen[8316]),
			.S(gen[8317]),
			.SE(gen[8318]),

			.SELF(gen[8222]),
			.cell_state(gen[8222])
		); 

/******************* CELL 8223 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8223 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8127]),
			.N(gen[8128]),
			.NE(gen[8129]),

			.O(gen[8222]),
			.E(gen[8224]),

			.SO(gen[8317]),
			.S(gen[8318]),
			.SE(gen[8319]),

			.SELF(gen[8223]),
			.cell_state(gen[8223])
		); 

/******************* CELL 8224 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8224 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8128]),
			.N(gen[8129]),
			.NE(gen[8130]),

			.O(gen[8223]),
			.E(gen[8225]),

			.SO(gen[8318]),
			.S(gen[8319]),
			.SE(gen[8320]),

			.SELF(gen[8224]),
			.cell_state(gen[8224])
		); 

/******************* CELL 8225 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8225 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8129]),
			.N(gen[8130]),
			.NE(gen[8131]),

			.O(gen[8224]),
			.E(gen[8226]),

			.SO(gen[8319]),
			.S(gen[8320]),
			.SE(gen[8321]),

			.SELF(gen[8225]),
			.cell_state(gen[8225])
		); 

/******************* CELL 8226 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8226 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8130]),
			.N(gen[8131]),
			.NE(gen[8132]),

			.O(gen[8225]),
			.E(gen[8227]),

			.SO(gen[8320]),
			.S(gen[8321]),
			.SE(gen[8322]),

			.SELF(gen[8226]),
			.cell_state(gen[8226])
		); 

/******************* CELL 8227 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8227 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8131]),
			.N(gen[8132]),
			.NE(gen[8133]),

			.O(gen[8226]),
			.E(gen[8228]),

			.SO(gen[8321]),
			.S(gen[8322]),
			.SE(gen[8323]),

			.SELF(gen[8227]),
			.cell_state(gen[8227])
		); 

/******************* CELL 8228 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8228 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8132]),
			.N(gen[8133]),
			.NE(gen[8134]),

			.O(gen[8227]),
			.E(gen[8229]),

			.SO(gen[8322]),
			.S(gen[8323]),
			.SE(gen[8324]),

			.SELF(gen[8228]),
			.cell_state(gen[8228])
		); 

/******************* CELL 8229 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8229 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8133]),
			.N(gen[8134]),
			.NE(gen[8135]),

			.O(gen[8228]),
			.E(gen[8230]),

			.SO(gen[8323]),
			.S(gen[8324]),
			.SE(gen[8325]),

			.SELF(gen[8229]),
			.cell_state(gen[8229])
		); 

/******************* CELL 8230 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8230 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8134]),
			.N(gen[8135]),
			.NE(gen[8136]),

			.O(gen[8229]),
			.E(gen[8231]),

			.SO(gen[8324]),
			.S(gen[8325]),
			.SE(gen[8326]),

			.SELF(gen[8230]),
			.cell_state(gen[8230])
		); 

/******************* CELL 8231 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8231 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8135]),
			.N(gen[8136]),
			.NE(gen[8137]),

			.O(gen[8230]),
			.E(gen[8232]),

			.SO(gen[8325]),
			.S(gen[8326]),
			.SE(gen[8327]),

			.SELF(gen[8231]),
			.cell_state(gen[8231])
		); 

/******************* CELL 8232 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8232 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8136]),
			.N(gen[8137]),
			.NE(gen[8138]),

			.O(gen[8231]),
			.E(gen[8233]),

			.SO(gen[8326]),
			.S(gen[8327]),
			.SE(gen[8328]),

			.SELF(gen[8232]),
			.cell_state(gen[8232])
		); 

/******************* CELL 8233 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8233 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8137]),
			.N(gen[8138]),
			.NE(gen[8139]),

			.O(gen[8232]),
			.E(gen[8234]),

			.SO(gen[8327]),
			.S(gen[8328]),
			.SE(gen[8329]),

			.SELF(gen[8233]),
			.cell_state(gen[8233])
		); 

/******************* CELL 8234 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8234 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8138]),
			.N(gen[8139]),
			.NE(gen[8140]),

			.O(gen[8233]),
			.E(gen[8235]),

			.SO(gen[8328]),
			.S(gen[8329]),
			.SE(gen[8330]),

			.SELF(gen[8234]),
			.cell_state(gen[8234])
		); 

/******************* CELL 8235 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8235 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8139]),
			.N(gen[8140]),
			.NE(gen[8141]),

			.O(gen[8234]),
			.E(gen[8236]),

			.SO(gen[8329]),
			.S(gen[8330]),
			.SE(gen[8331]),

			.SELF(gen[8235]),
			.cell_state(gen[8235])
		); 

/******************* CELL 8236 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8236 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8140]),
			.N(gen[8141]),
			.NE(gen[8142]),

			.O(gen[8235]),
			.E(gen[8237]),

			.SO(gen[8330]),
			.S(gen[8331]),
			.SE(gen[8332]),

			.SELF(gen[8236]),
			.cell_state(gen[8236])
		); 

/******************* CELL 8237 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8237 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8141]),
			.N(gen[8142]),
			.NE(gen[8143]),

			.O(gen[8236]),
			.E(gen[8238]),

			.SO(gen[8331]),
			.S(gen[8332]),
			.SE(gen[8333]),

			.SELF(gen[8237]),
			.cell_state(gen[8237])
		); 

/******************* CELL 8238 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8238 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8142]),
			.N(gen[8143]),
			.NE(gen[8144]),

			.O(gen[8237]),
			.E(gen[8239]),

			.SO(gen[8332]),
			.S(gen[8333]),
			.SE(gen[8334]),

			.SELF(gen[8238]),
			.cell_state(gen[8238])
		); 

/******************* CELL 8239 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8239 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8143]),
			.N(gen[8144]),
			.NE(gen[8145]),

			.O(gen[8238]),
			.E(gen[8240]),

			.SO(gen[8333]),
			.S(gen[8334]),
			.SE(gen[8335]),

			.SELF(gen[8239]),
			.cell_state(gen[8239])
		); 

/******************* CELL 8240 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8240 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8144]),
			.N(gen[8145]),
			.NE(gen[8146]),

			.O(gen[8239]),
			.E(gen[8241]),

			.SO(gen[8334]),
			.S(gen[8335]),
			.SE(gen[8336]),

			.SELF(gen[8240]),
			.cell_state(gen[8240])
		); 

/******************* CELL 8241 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8241 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8145]),
			.N(gen[8146]),
			.NE(gen[8147]),

			.O(gen[8240]),
			.E(gen[8242]),

			.SO(gen[8335]),
			.S(gen[8336]),
			.SE(gen[8337]),

			.SELF(gen[8241]),
			.cell_state(gen[8241])
		); 

/******************* CELL 8242 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8242 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8146]),
			.N(gen[8147]),
			.NE(gen[8148]),

			.O(gen[8241]),
			.E(gen[8243]),

			.SO(gen[8336]),
			.S(gen[8337]),
			.SE(gen[8338]),

			.SELF(gen[8242]),
			.cell_state(gen[8242])
		); 

/******************* CELL 8243 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8243 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8147]),
			.N(gen[8148]),
			.NE(gen[8149]),

			.O(gen[8242]),
			.E(gen[8244]),

			.SO(gen[8337]),
			.S(gen[8338]),
			.SE(gen[8339]),

			.SELF(gen[8243]),
			.cell_state(gen[8243])
		); 

/******************* CELL 8244 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8244 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8148]),
			.N(gen[8149]),
			.NE(gen[8150]),

			.O(gen[8243]),
			.E(gen[8245]),

			.SO(gen[8338]),
			.S(gen[8339]),
			.SE(gen[8340]),

			.SELF(gen[8244]),
			.cell_state(gen[8244])
		); 

/******************* CELL 8245 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8245 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8149]),
			.N(gen[8150]),
			.NE(gen[8151]),

			.O(gen[8244]),
			.E(gen[8246]),

			.SO(gen[8339]),
			.S(gen[8340]),
			.SE(gen[8341]),

			.SELF(gen[8245]),
			.cell_state(gen[8245])
		); 

/******************* CELL 8246 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8246 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8150]),
			.N(gen[8151]),
			.NE(gen[8152]),

			.O(gen[8245]),
			.E(gen[8247]),

			.SO(gen[8340]),
			.S(gen[8341]),
			.SE(gen[8342]),

			.SELF(gen[8246]),
			.cell_state(gen[8246])
		); 

/******************* CELL 8247 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8247 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8151]),
			.N(gen[8152]),
			.NE(gen[8153]),

			.O(gen[8246]),
			.E(gen[8248]),

			.SO(gen[8341]),
			.S(gen[8342]),
			.SE(gen[8343]),

			.SELF(gen[8247]),
			.cell_state(gen[8247])
		); 

/******************* CELL 8248 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8248 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8152]),
			.N(gen[8153]),
			.NE(gen[8154]),

			.O(gen[8247]),
			.E(gen[8249]),

			.SO(gen[8342]),
			.S(gen[8343]),
			.SE(gen[8344]),

			.SELF(gen[8248]),
			.cell_state(gen[8248])
		); 

/******************* CELL 8249 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8249 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8153]),
			.N(gen[8154]),
			.NE(gen[8155]),

			.O(gen[8248]),
			.E(gen[8250]),

			.SO(gen[8343]),
			.S(gen[8344]),
			.SE(gen[8345]),

			.SELF(gen[8249]),
			.cell_state(gen[8249])
		); 

/******************* CELL 8250 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8250 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8154]),
			.N(gen[8155]),
			.NE(gen[8156]),

			.O(gen[8249]),
			.E(gen[8251]),

			.SO(gen[8344]),
			.S(gen[8345]),
			.SE(gen[8346]),

			.SELF(gen[8250]),
			.cell_state(gen[8250])
		); 

/******************* CELL 8251 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8251 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8155]),
			.N(gen[8156]),
			.NE(gen[8157]),

			.O(gen[8250]),
			.E(gen[8252]),

			.SO(gen[8345]),
			.S(gen[8346]),
			.SE(gen[8347]),

			.SELF(gen[8251]),
			.cell_state(gen[8251])
		); 

/******************* CELL 8252 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8252 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8156]),
			.N(gen[8157]),
			.NE(gen[8158]),

			.O(gen[8251]),
			.E(gen[8253]),

			.SO(gen[8346]),
			.S(gen[8347]),
			.SE(gen[8348]),

			.SELF(gen[8252]),
			.cell_state(gen[8252])
		); 

/******************* CELL 8253 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8253 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8157]),
			.N(gen[8158]),
			.NE(gen[8159]),

			.O(gen[8252]),
			.E(gen[8254]),

			.SO(gen[8347]),
			.S(gen[8348]),
			.SE(gen[8349]),

			.SELF(gen[8253]),
			.cell_state(gen[8253])
		); 

/******************* CELL 8254 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8254 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8158]),
			.N(gen[8159]),
			.NE(gen[8160]),

			.O(gen[8253]),
			.E(gen[8255]),

			.SO(gen[8348]),
			.S(gen[8349]),
			.SE(gen[8350]),

			.SELF(gen[8254]),
			.cell_state(gen[8254])
		); 

/******************* CELL 8255 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8255 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8159]),
			.N(gen[8160]),
			.NE(gen[8161]),

			.O(gen[8254]),
			.E(gen[8256]),

			.SO(gen[8349]),
			.S(gen[8350]),
			.SE(gen[8351]),

			.SELF(gen[8255]),
			.cell_state(gen[8255])
		); 

/******************* CELL 8256 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8256 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8160]),
			.N(gen[8161]),
			.NE(gen[8162]),

			.O(gen[8255]),
			.E(gen[8257]),

			.SO(gen[8350]),
			.S(gen[8351]),
			.SE(gen[8352]),

			.SELF(gen[8256]),
			.cell_state(gen[8256])
		); 

/******************* CELL 8257 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8257 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8161]),
			.N(gen[8162]),
			.NE(gen[8163]),

			.O(gen[8256]),
			.E(gen[8258]),

			.SO(gen[8351]),
			.S(gen[8352]),
			.SE(gen[8353]),

			.SELF(gen[8257]),
			.cell_state(gen[8257])
		); 

/******************* CELL 8258 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8258 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8162]),
			.N(gen[8163]),
			.NE(gen[8164]),

			.O(gen[8257]),
			.E(gen[8259]),

			.SO(gen[8352]),
			.S(gen[8353]),
			.SE(gen[8354]),

			.SELF(gen[8258]),
			.cell_state(gen[8258])
		); 

/******************* CELL 8259 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8259 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8163]),
			.N(gen[8164]),
			.NE(gen[8165]),

			.O(gen[8258]),
			.E(gen[8260]),

			.SO(gen[8353]),
			.S(gen[8354]),
			.SE(gen[8355]),

			.SELF(gen[8259]),
			.cell_state(gen[8259])
		); 

/******************* CELL 8260 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8260 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8164]),
			.N(gen[8165]),
			.NE(gen[8166]),

			.O(gen[8259]),
			.E(gen[8261]),

			.SO(gen[8354]),
			.S(gen[8355]),
			.SE(gen[8356]),

			.SELF(gen[8260]),
			.cell_state(gen[8260])
		); 

/******************* CELL 8261 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8261 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8165]),
			.N(gen[8166]),
			.NE(gen[8167]),

			.O(gen[8260]),
			.E(gen[8262]),

			.SO(gen[8355]),
			.S(gen[8356]),
			.SE(gen[8357]),

			.SELF(gen[8261]),
			.cell_state(gen[8261])
		); 

/******************* CELL 8262 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8262 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8166]),
			.N(gen[8167]),
			.NE(gen[8168]),

			.O(gen[8261]),
			.E(gen[8263]),

			.SO(gen[8356]),
			.S(gen[8357]),
			.SE(gen[8358]),

			.SELF(gen[8262]),
			.cell_state(gen[8262])
		); 

/******************* CELL 8263 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8263 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8167]),
			.N(gen[8168]),
			.NE(gen[8169]),

			.O(gen[8262]),
			.E(gen[8264]),

			.SO(gen[8357]),
			.S(gen[8358]),
			.SE(gen[8359]),

			.SELF(gen[8263]),
			.cell_state(gen[8263])
		); 

/******************* CELL 8264 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8264 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8168]),
			.N(gen[8169]),
			.NE(gen[8168]),

			.O(gen[8263]),
			.E(gen[8263]),

			.SO(gen[8358]),
			.S(gen[8359]),
			.SE(gen[8358]),

			.SELF(gen[8264]),
			.cell_state(gen[8264])
		); 

/******************* CELL 8265 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8265 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8171]),
			.N(gen[8170]),
			.NE(gen[8171]),

			.O(gen[8266]),
			.E(gen[8266]),

			.SO(gen[8361]),
			.S(gen[8360]),
			.SE(gen[8361]),

			.SELF(gen[8265]),
			.cell_state(gen[8265])
		); 

/******************* CELL 8266 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8266 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8170]),
			.N(gen[8171]),
			.NE(gen[8172]),

			.O(gen[8265]),
			.E(gen[8267]),

			.SO(gen[8360]),
			.S(gen[8361]),
			.SE(gen[8362]),

			.SELF(gen[8266]),
			.cell_state(gen[8266])
		); 

/******************* CELL 8267 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8267 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8171]),
			.N(gen[8172]),
			.NE(gen[8173]),

			.O(gen[8266]),
			.E(gen[8268]),

			.SO(gen[8361]),
			.S(gen[8362]),
			.SE(gen[8363]),

			.SELF(gen[8267]),
			.cell_state(gen[8267])
		); 

/******************* CELL 8268 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8268 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8172]),
			.N(gen[8173]),
			.NE(gen[8174]),

			.O(gen[8267]),
			.E(gen[8269]),

			.SO(gen[8362]),
			.S(gen[8363]),
			.SE(gen[8364]),

			.SELF(gen[8268]),
			.cell_state(gen[8268])
		); 

/******************* CELL 8269 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8269 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8173]),
			.N(gen[8174]),
			.NE(gen[8175]),

			.O(gen[8268]),
			.E(gen[8270]),

			.SO(gen[8363]),
			.S(gen[8364]),
			.SE(gen[8365]),

			.SELF(gen[8269]),
			.cell_state(gen[8269])
		); 

/******************* CELL 8270 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8270 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8174]),
			.N(gen[8175]),
			.NE(gen[8176]),

			.O(gen[8269]),
			.E(gen[8271]),

			.SO(gen[8364]),
			.S(gen[8365]),
			.SE(gen[8366]),

			.SELF(gen[8270]),
			.cell_state(gen[8270])
		); 

/******************* CELL 8271 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8271 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8175]),
			.N(gen[8176]),
			.NE(gen[8177]),

			.O(gen[8270]),
			.E(gen[8272]),

			.SO(gen[8365]),
			.S(gen[8366]),
			.SE(gen[8367]),

			.SELF(gen[8271]),
			.cell_state(gen[8271])
		); 

/******************* CELL 8272 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8272 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8176]),
			.N(gen[8177]),
			.NE(gen[8178]),

			.O(gen[8271]),
			.E(gen[8273]),

			.SO(gen[8366]),
			.S(gen[8367]),
			.SE(gen[8368]),

			.SELF(gen[8272]),
			.cell_state(gen[8272])
		); 

/******************* CELL 8273 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8273 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8177]),
			.N(gen[8178]),
			.NE(gen[8179]),

			.O(gen[8272]),
			.E(gen[8274]),

			.SO(gen[8367]),
			.S(gen[8368]),
			.SE(gen[8369]),

			.SELF(gen[8273]),
			.cell_state(gen[8273])
		); 

/******************* CELL 8274 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8274 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8178]),
			.N(gen[8179]),
			.NE(gen[8180]),

			.O(gen[8273]),
			.E(gen[8275]),

			.SO(gen[8368]),
			.S(gen[8369]),
			.SE(gen[8370]),

			.SELF(gen[8274]),
			.cell_state(gen[8274])
		); 

/******************* CELL 8275 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8275 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8179]),
			.N(gen[8180]),
			.NE(gen[8181]),

			.O(gen[8274]),
			.E(gen[8276]),

			.SO(gen[8369]),
			.S(gen[8370]),
			.SE(gen[8371]),

			.SELF(gen[8275]),
			.cell_state(gen[8275])
		); 

/******************* CELL 8276 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8276 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8180]),
			.N(gen[8181]),
			.NE(gen[8182]),

			.O(gen[8275]),
			.E(gen[8277]),

			.SO(gen[8370]),
			.S(gen[8371]),
			.SE(gen[8372]),

			.SELF(gen[8276]),
			.cell_state(gen[8276])
		); 

/******************* CELL 8277 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8277 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8181]),
			.N(gen[8182]),
			.NE(gen[8183]),

			.O(gen[8276]),
			.E(gen[8278]),

			.SO(gen[8371]),
			.S(gen[8372]),
			.SE(gen[8373]),

			.SELF(gen[8277]),
			.cell_state(gen[8277])
		); 

/******************* CELL 8278 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8278 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8182]),
			.N(gen[8183]),
			.NE(gen[8184]),

			.O(gen[8277]),
			.E(gen[8279]),

			.SO(gen[8372]),
			.S(gen[8373]),
			.SE(gen[8374]),

			.SELF(gen[8278]),
			.cell_state(gen[8278])
		); 

/******************* CELL 8279 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8279 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8183]),
			.N(gen[8184]),
			.NE(gen[8185]),

			.O(gen[8278]),
			.E(gen[8280]),

			.SO(gen[8373]),
			.S(gen[8374]),
			.SE(gen[8375]),

			.SELF(gen[8279]),
			.cell_state(gen[8279])
		); 

/******************* CELL 8280 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8280 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8184]),
			.N(gen[8185]),
			.NE(gen[8186]),

			.O(gen[8279]),
			.E(gen[8281]),

			.SO(gen[8374]),
			.S(gen[8375]),
			.SE(gen[8376]),

			.SELF(gen[8280]),
			.cell_state(gen[8280])
		); 

/******************* CELL 8281 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8281 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8185]),
			.N(gen[8186]),
			.NE(gen[8187]),

			.O(gen[8280]),
			.E(gen[8282]),

			.SO(gen[8375]),
			.S(gen[8376]),
			.SE(gen[8377]),

			.SELF(gen[8281]),
			.cell_state(gen[8281])
		); 

/******************* CELL 8282 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8282 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8186]),
			.N(gen[8187]),
			.NE(gen[8188]),

			.O(gen[8281]),
			.E(gen[8283]),

			.SO(gen[8376]),
			.S(gen[8377]),
			.SE(gen[8378]),

			.SELF(gen[8282]),
			.cell_state(gen[8282])
		); 

/******************* CELL 8283 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8283 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8187]),
			.N(gen[8188]),
			.NE(gen[8189]),

			.O(gen[8282]),
			.E(gen[8284]),

			.SO(gen[8377]),
			.S(gen[8378]),
			.SE(gen[8379]),

			.SELF(gen[8283]),
			.cell_state(gen[8283])
		); 

/******************* CELL 8284 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8284 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8188]),
			.N(gen[8189]),
			.NE(gen[8190]),

			.O(gen[8283]),
			.E(gen[8285]),

			.SO(gen[8378]),
			.S(gen[8379]),
			.SE(gen[8380]),

			.SELF(gen[8284]),
			.cell_state(gen[8284])
		); 

/******************* CELL 8285 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8285 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8189]),
			.N(gen[8190]),
			.NE(gen[8191]),

			.O(gen[8284]),
			.E(gen[8286]),

			.SO(gen[8379]),
			.S(gen[8380]),
			.SE(gen[8381]),

			.SELF(gen[8285]),
			.cell_state(gen[8285])
		); 

/******************* CELL 8286 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8286 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8190]),
			.N(gen[8191]),
			.NE(gen[8192]),

			.O(gen[8285]),
			.E(gen[8287]),

			.SO(gen[8380]),
			.S(gen[8381]),
			.SE(gen[8382]),

			.SELF(gen[8286]),
			.cell_state(gen[8286])
		); 

/******************* CELL 8287 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8287 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8191]),
			.N(gen[8192]),
			.NE(gen[8193]),

			.O(gen[8286]),
			.E(gen[8288]),

			.SO(gen[8381]),
			.S(gen[8382]),
			.SE(gen[8383]),

			.SELF(gen[8287]),
			.cell_state(gen[8287])
		); 

/******************* CELL 8288 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8288 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8192]),
			.N(gen[8193]),
			.NE(gen[8194]),

			.O(gen[8287]),
			.E(gen[8289]),

			.SO(gen[8382]),
			.S(gen[8383]),
			.SE(gen[8384]),

			.SELF(gen[8288]),
			.cell_state(gen[8288])
		); 

/******************* CELL 8289 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8289 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8193]),
			.N(gen[8194]),
			.NE(gen[8195]),

			.O(gen[8288]),
			.E(gen[8290]),

			.SO(gen[8383]),
			.S(gen[8384]),
			.SE(gen[8385]),

			.SELF(gen[8289]),
			.cell_state(gen[8289])
		); 

/******************* CELL 8290 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8290 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8194]),
			.N(gen[8195]),
			.NE(gen[8196]),

			.O(gen[8289]),
			.E(gen[8291]),

			.SO(gen[8384]),
			.S(gen[8385]),
			.SE(gen[8386]),

			.SELF(gen[8290]),
			.cell_state(gen[8290])
		); 

/******************* CELL 8291 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8291 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8195]),
			.N(gen[8196]),
			.NE(gen[8197]),

			.O(gen[8290]),
			.E(gen[8292]),

			.SO(gen[8385]),
			.S(gen[8386]),
			.SE(gen[8387]),

			.SELF(gen[8291]),
			.cell_state(gen[8291])
		); 

/******************* CELL 8292 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8292 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8196]),
			.N(gen[8197]),
			.NE(gen[8198]),

			.O(gen[8291]),
			.E(gen[8293]),

			.SO(gen[8386]),
			.S(gen[8387]),
			.SE(gen[8388]),

			.SELF(gen[8292]),
			.cell_state(gen[8292])
		); 

/******************* CELL 8293 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8293 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8197]),
			.N(gen[8198]),
			.NE(gen[8199]),

			.O(gen[8292]),
			.E(gen[8294]),

			.SO(gen[8387]),
			.S(gen[8388]),
			.SE(gen[8389]),

			.SELF(gen[8293]),
			.cell_state(gen[8293])
		); 

/******************* CELL 8294 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8294 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8198]),
			.N(gen[8199]),
			.NE(gen[8200]),

			.O(gen[8293]),
			.E(gen[8295]),

			.SO(gen[8388]),
			.S(gen[8389]),
			.SE(gen[8390]),

			.SELF(gen[8294]),
			.cell_state(gen[8294])
		); 

/******************* CELL 8295 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8295 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8199]),
			.N(gen[8200]),
			.NE(gen[8201]),

			.O(gen[8294]),
			.E(gen[8296]),

			.SO(gen[8389]),
			.S(gen[8390]),
			.SE(gen[8391]),

			.SELF(gen[8295]),
			.cell_state(gen[8295])
		); 

/******************* CELL 8296 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8296 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8200]),
			.N(gen[8201]),
			.NE(gen[8202]),

			.O(gen[8295]),
			.E(gen[8297]),

			.SO(gen[8390]),
			.S(gen[8391]),
			.SE(gen[8392]),

			.SELF(gen[8296]),
			.cell_state(gen[8296])
		); 

/******************* CELL 8297 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8297 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8201]),
			.N(gen[8202]),
			.NE(gen[8203]),

			.O(gen[8296]),
			.E(gen[8298]),

			.SO(gen[8391]),
			.S(gen[8392]),
			.SE(gen[8393]),

			.SELF(gen[8297]),
			.cell_state(gen[8297])
		); 

/******************* CELL 8298 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8298 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8202]),
			.N(gen[8203]),
			.NE(gen[8204]),

			.O(gen[8297]),
			.E(gen[8299]),

			.SO(gen[8392]),
			.S(gen[8393]),
			.SE(gen[8394]),

			.SELF(gen[8298]),
			.cell_state(gen[8298])
		); 

/******************* CELL 8299 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8299 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8203]),
			.N(gen[8204]),
			.NE(gen[8205]),

			.O(gen[8298]),
			.E(gen[8300]),

			.SO(gen[8393]),
			.S(gen[8394]),
			.SE(gen[8395]),

			.SELF(gen[8299]),
			.cell_state(gen[8299])
		); 

/******************* CELL 8300 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8300 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8204]),
			.N(gen[8205]),
			.NE(gen[8206]),

			.O(gen[8299]),
			.E(gen[8301]),

			.SO(gen[8394]),
			.S(gen[8395]),
			.SE(gen[8396]),

			.SELF(gen[8300]),
			.cell_state(gen[8300])
		); 

/******************* CELL 8301 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8301 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8205]),
			.N(gen[8206]),
			.NE(gen[8207]),

			.O(gen[8300]),
			.E(gen[8302]),

			.SO(gen[8395]),
			.S(gen[8396]),
			.SE(gen[8397]),

			.SELF(gen[8301]),
			.cell_state(gen[8301])
		); 

/******************* CELL 8302 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8302 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8206]),
			.N(gen[8207]),
			.NE(gen[8208]),

			.O(gen[8301]),
			.E(gen[8303]),

			.SO(gen[8396]),
			.S(gen[8397]),
			.SE(gen[8398]),

			.SELF(gen[8302]),
			.cell_state(gen[8302])
		); 

/******************* CELL 8303 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8303 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8207]),
			.N(gen[8208]),
			.NE(gen[8209]),

			.O(gen[8302]),
			.E(gen[8304]),

			.SO(gen[8397]),
			.S(gen[8398]),
			.SE(gen[8399]),

			.SELF(gen[8303]),
			.cell_state(gen[8303])
		); 

/******************* CELL 8304 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8304 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8208]),
			.N(gen[8209]),
			.NE(gen[8210]),

			.O(gen[8303]),
			.E(gen[8305]),

			.SO(gen[8398]),
			.S(gen[8399]),
			.SE(gen[8400]),

			.SELF(gen[8304]),
			.cell_state(gen[8304])
		); 

/******************* CELL 8305 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8305 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8209]),
			.N(gen[8210]),
			.NE(gen[8211]),

			.O(gen[8304]),
			.E(gen[8306]),

			.SO(gen[8399]),
			.S(gen[8400]),
			.SE(gen[8401]),

			.SELF(gen[8305]),
			.cell_state(gen[8305])
		); 

/******************* CELL 8306 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8306 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8210]),
			.N(gen[8211]),
			.NE(gen[8212]),

			.O(gen[8305]),
			.E(gen[8307]),

			.SO(gen[8400]),
			.S(gen[8401]),
			.SE(gen[8402]),

			.SELF(gen[8306]),
			.cell_state(gen[8306])
		); 

/******************* CELL 8307 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8307 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8211]),
			.N(gen[8212]),
			.NE(gen[8213]),

			.O(gen[8306]),
			.E(gen[8308]),

			.SO(gen[8401]),
			.S(gen[8402]),
			.SE(gen[8403]),

			.SELF(gen[8307]),
			.cell_state(gen[8307])
		); 

/******************* CELL 8308 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8308 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8212]),
			.N(gen[8213]),
			.NE(gen[8214]),

			.O(gen[8307]),
			.E(gen[8309]),

			.SO(gen[8402]),
			.S(gen[8403]),
			.SE(gen[8404]),

			.SELF(gen[8308]),
			.cell_state(gen[8308])
		); 

/******************* CELL 8309 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8309 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8213]),
			.N(gen[8214]),
			.NE(gen[8215]),

			.O(gen[8308]),
			.E(gen[8310]),

			.SO(gen[8403]),
			.S(gen[8404]),
			.SE(gen[8405]),

			.SELF(gen[8309]),
			.cell_state(gen[8309])
		); 

/******************* CELL 8310 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8310 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8214]),
			.N(gen[8215]),
			.NE(gen[8216]),

			.O(gen[8309]),
			.E(gen[8311]),

			.SO(gen[8404]),
			.S(gen[8405]),
			.SE(gen[8406]),

			.SELF(gen[8310]),
			.cell_state(gen[8310])
		); 

/******************* CELL 8311 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8311 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8215]),
			.N(gen[8216]),
			.NE(gen[8217]),

			.O(gen[8310]),
			.E(gen[8312]),

			.SO(gen[8405]),
			.S(gen[8406]),
			.SE(gen[8407]),

			.SELF(gen[8311]),
			.cell_state(gen[8311])
		); 

/******************* CELL 8312 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8312 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8216]),
			.N(gen[8217]),
			.NE(gen[8218]),

			.O(gen[8311]),
			.E(gen[8313]),

			.SO(gen[8406]),
			.S(gen[8407]),
			.SE(gen[8408]),

			.SELF(gen[8312]),
			.cell_state(gen[8312])
		); 

/******************* CELL 8313 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8313 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8217]),
			.N(gen[8218]),
			.NE(gen[8219]),

			.O(gen[8312]),
			.E(gen[8314]),

			.SO(gen[8407]),
			.S(gen[8408]),
			.SE(gen[8409]),

			.SELF(gen[8313]),
			.cell_state(gen[8313])
		); 

/******************* CELL 8314 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8314 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8218]),
			.N(gen[8219]),
			.NE(gen[8220]),

			.O(gen[8313]),
			.E(gen[8315]),

			.SO(gen[8408]),
			.S(gen[8409]),
			.SE(gen[8410]),

			.SELF(gen[8314]),
			.cell_state(gen[8314])
		); 

/******************* CELL 8315 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8315 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8219]),
			.N(gen[8220]),
			.NE(gen[8221]),

			.O(gen[8314]),
			.E(gen[8316]),

			.SO(gen[8409]),
			.S(gen[8410]),
			.SE(gen[8411]),

			.SELF(gen[8315]),
			.cell_state(gen[8315])
		); 

/******************* CELL 8316 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8316 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8220]),
			.N(gen[8221]),
			.NE(gen[8222]),

			.O(gen[8315]),
			.E(gen[8317]),

			.SO(gen[8410]),
			.S(gen[8411]),
			.SE(gen[8412]),

			.SELF(gen[8316]),
			.cell_state(gen[8316])
		); 

/******************* CELL 8317 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8317 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8221]),
			.N(gen[8222]),
			.NE(gen[8223]),

			.O(gen[8316]),
			.E(gen[8318]),

			.SO(gen[8411]),
			.S(gen[8412]),
			.SE(gen[8413]),

			.SELF(gen[8317]),
			.cell_state(gen[8317])
		); 

/******************* CELL 8318 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8318 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8222]),
			.N(gen[8223]),
			.NE(gen[8224]),

			.O(gen[8317]),
			.E(gen[8319]),

			.SO(gen[8412]),
			.S(gen[8413]),
			.SE(gen[8414]),

			.SELF(gen[8318]),
			.cell_state(gen[8318])
		); 

/******************* CELL 8319 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8319 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8223]),
			.N(gen[8224]),
			.NE(gen[8225]),

			.O(gen[8318]),
			.E(gen[8320]),

			.SO(gen[8413]),
			.S(gen[8414]),
			.SE(gen[8415]),

			.SELF(gen[8319]),
			.cell_state(gen[8319])
		); 

/******************* CELL 8320 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8320 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8224]),
			.N(gen[8225]),
			.NE(gen[8226]),

			.O(gen[8319]),
			.E(gen[8321]),

			.SO(gen[8414]),
			.S(gen[8415]),
			.SE(gen[8416]),

			.SELF(gen[8320]),
			.cell_state(gen[8320])
		); 

/******************* CELL 8321 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8321 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8225]),
			.N(gen[8226]),
			.NE(gen[8227]),

			.O(gen[8320]),
			.E(gen[8322]),

			.SO(gen[8415]),
			.S(gen[8416]),
			.SE(gen[8417]),

			.SELF(gen[8321]),
			.cell_state(gen[8321])
		); 

/******************* CELL 8322 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8322 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8226]),
			.N(gen[8227]),
			.NE(gen[8228]),

			.O(gen[8321]),
			.E(gen[8323]),

			.SO(gen[8416]),
			.S(gen[8417]),
			.SE(gen[8418]),

			.SELF(gen[8322]),
			.cell_state(gen[8322])
		); 

/******************* CELL 8323 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8323 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8227]),
			.N(gen[8228]),
			.NE(gen[8229]),

			.O(gen[8322]),
			.E(gen[8324]),

			.SO(gen[8417]),
			.S(gen[8418]),
			.SE(gen[8419]),

			.SELF(gen[8323]),
			.cell_state(gen[8323])
		); 

/******************* CELL 8324 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8324 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8228]),
			.N(gen[8229]),
			.NE(gen[8230]),

			.O(gen[8323]),
			.E(gen[8325]),

			.SO(gen[8418]),
			.S(gen[8419]),
			.SE(gen[8420]),

			.SELF(gen[8324]),
			.cell_state(gen[8324])
		); 

/******************* CELL 8325 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8325 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8229]),
			.N(gen[8230]),
			.NE(gen[8231]),

			.O(gen[8324]),
			.E(gen[8326]),

			.SO(gen[8419]),
			.S(gen[8420]),
			.SE(gen[8421]),

			.SELF(gen[8325]),
			.cell_state(gen[8325])
		); 

/******************* CELL 8326 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8326 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8230]),
			.N(gen[8231]),
			.NE(gen[8232]),

			.O(gen[8325]),
			.E(gen[8327]),

			.SO(gen[8420]),
			.S(gen[8421]),
			.SE(gen[8422]),

			.SELF(gen[8326]),
			.cell_state(gen[8326])
		); 

/******************* CELL 8327 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8327 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8231]),
			.N(gen[8232]),
			.NE(gen[8233]),

			.O(gen[8326]),
			.E(gen[8328]),

			.SO(gen[8421]),
			.S(gen[8422]),
			.SE(gen[8423]),

			.SELF(gen[8327]),
			.cell_state(gen[8327])
		); 

/******************* CELL 8328 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8328 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8232]),
			.N(gen[8233]),
			.NE(gen[8234]),

			.O(gen[8327]),
			.E(gen[8329]),

			.SO(gen[8422]),
			.S(gen[8423]),
			.SE(gen[8424]),

			.SELF(gen[8328]),
			.cell_state(gen[8328])
		); 

/******************* CELL 8329 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8329 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8233]),
			.N(gen[8234]),
			.NE(gen[8235]),

			.O(gen[8328]),
			.E(gen[8330]),

			.SO(gen[8423]),
			.S(gen[8424]),
			.SE(gen[8425]),

			.SELF(gen[8329]),
			.cell_state(gen[8329])
		); 

/******************* CELL 8330 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8330 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8234]),
			.N(gen[8235]),
			.NE(gen[8236]),

			.O(gen[8329]),
			.E(gen[8331]),

			.SO(gen[8424]),
			.S(gen[8425]),
			.SE(gen[8426]),

			.SELF(gen[8330]),
			.cell_state(gen[8330])
		); 

/******************* CELL 8331 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8331 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8235]),
			.N(gen[8236]),
			.NE(gen[8237]),

			.O(gen[8330]),
			.E(gen[8332]),

			.SO(gen[8425]),
			.S(gen[8426]),
			.SE(gen[8427]),

			.SELF(gen[8331]),
			.cell_state(gen[8331])
		); 

/******************* CELL 8332 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8332 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8236]),
			.N(gen[8237]),
			.NE(gen[8238]),

			.O(gen[8331]),
			.E(gen[8333]),

			.SO(gen[8426]),
			.S(gen[8427]),
			.SE(gen[8428]),

			.SELF(gen[8332]),
			.cell_state(gen[8332])
		); 

/******************* CELL 8333 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8333 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8237]),
			.N(gen[8238]),
			.NE(gen[8239]),

			.O(gen[8332]),
			.E(gen[8334]),

			.SO(gen[8427]),
			.S(gen[8428]),
			.SE(gen[8429]),

			.SELF(gen[8333]),
			.cell_state(gen[8333])
		); 

/******************* CELL 8334 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8334 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8238]),
			.N(gen[8239]),
			.NE(gen[8240]),

			.O(gen[8333]),
			.E(gen[8335]),

			.SO(gen[8428]),
			.S(gen[8429]),
			.SE(gen[8430]),

			.SELF(gen[8334]),
			.cell_state(gen[8334])
		); 

/******************* CELL 8335 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8335 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8239]),
			.N(gen[8240]),
			.NE(gen[8241]),

			.O(gen[8334]),
			.E(gen[8336]),

			.SO(gen[8429]),
			.S(gen[8430]),
			.SE(gen[8431]),

			.SELF(gen[8335]),
			.cell_state(gen[8335])
		); 

/******************* CELL 8336 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8336 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8240]),
			.N(gen[8241]),
			.NE(gen[8242]),

			.O(gen[8335]),
			.E(gen[8337]),

			.SO(gen[8430]),
			.S(gen[8431]),
			.SE(gen[8432]),

			.SELF(gen[8336]),
			.cell_state(gen[8336])
		); 

/******************* CELL 8337 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8337 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8241]),
			.N(gen[8242]),
			.NE(gen[8243]),

			.O(gen[8336]),
			.E(gen[8338]),

			.SO(gen[8431]),
			.S(gen[8432]),
			.SE(gen[8433]),

			.SELF(gen[8337]),
			.cell_state(gen[8337])
		); 

/******************* CELL 8338 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8338 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8242]),
			.N(gen[8243]),
			.NE(gen[8244]),

			.O(gen[8337]),
			.E(gen[8339]),

			.SO(gen[8432]),
			.S(gen[8433]),
			.SE(gen[8434]),

			.SELF(gen[8338]),
			.cell_state(gen[8338])
		); 

/******************* CELL 8339 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8339 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8243]),
			.N(gen[8244]),
			.NE(gen[8245]),

			.O(gen[8338]),
			.E(gen[8340]),

			.SO(gen[8433]),
			.S(gen[8434]),
			.SE(gen[8435]),

			.SELF(gen[8339]),
			.cell_state(gen[8339])
		); 

/******************* CELL 8340 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8340 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8244]),
			.N(gen[8245]),
			.NE(gen[8246]),

			.O(gen[8339]),
			.E(gen[8341]),

			.SO(gen[8434]),
			.S(gen[8435]),
			.SE(gen[8436]),

			.SELF(gen[8340]),
			.cell_state(gen[8340])
		); 

/******************* CELL 8341 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8341 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8245]),
			.N(gen[8246]),
			.NE(gen[8247]),

			.O(gen[8340]),
			.E(gen[8342]),

			.SO(gen[8435]),
			.S(gen[8436]),
			.SE(gen[8437]),

			.SELF(gen[8341]),
			.cell_state(gen[8341])
		); 

/******************* CELL 8342 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8342 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8246]),
			.N(gen[8247]),
			.NE(gen[8248]),

			.O(gen[8341]),
			.E(gen[8343]),

			.SO(gen[8436]),
			.S(gen[8437]),
			.SE(gen[8438]),

			.SELF(gen[8342]),
			.cell_state(gen[8342])
		); 

/******************* CELL 8343 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8343 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8247]),
			.N(gen[8248]),
			.NE(gen[8249]),

			.O(gen[8342]),
			.E(gen[8344]),

			.SO(gen[8437]),
			.S(gen[8438]),
			.SE(gen[8439]),

			.SELF(gen[8343]),
			.cell_state(gen[8343])
		); 

/******************* CELL 8344 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8344 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8248]),
			.N(gen[8249]),
			.NE(gen[8250]),

			.O(gen[8343]),
			.E(gen[8345]),

			.SO(gen[8438]),
			.S(gen[8439]),
			.SE(gen[8440]),

			.SELF(gen[8344]),
			.cell_state(gen[8344])
		); 

/******************* CELL 8345 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8345 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8249]),
			.N(gen[8250]),
			.NE(gen[8251]),

			.O(gen[8344]),
			.E(gen[8346]),

			.SO(gen[8439]),
			.S(gen[8440]),
			.SE(gen[8441]),

			.SELF(gen[8345]),
			.cell_state(gen[8345])
		); 

/******************* CELL 8346 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8346 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8250]),
			.N(gen[8251]),
			.NE(gen[8252]),

			.O(gen[8345]),
			.E(gen[8347]),

			.SO(gen[8440]),
			.S(gen[8441]),
			.SE(gen[8442]),

			.SELF(gen[8346]),
			.cell_state(gen[8346])
		); 

/******************* CELL 8347 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8347 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8251]),
			.N(gen[8252]),
			.NE(gen[8253]),

			.O(gen[8346]),
			.E(gen[8348]),

			.SO(gen[8441]),
			.S(gen[8442]),
			.SE(gen[8443]),

			.SELF(gen[8347]),
			.cell_state(gen[8347])
		); 

/******************* CELL 8348 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8348 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8252]),
			.N(gen[8253]),
			.NE(gen[8254]),

			.O(gen[8347]),
			.E(gen[8349]),

			.SO(gen[8442]),
			.S(gen[8443]),
			.SE(gen[8444]),

			.SELF(gen[8348]),
			.cell_state(gen[8348])
		); 

/******************* CELL 8349 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8349 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8253]),
			.N(gen[8254]),
			.NE(gen[8255]),

			.O(gen[8348]),
			.E(gen[8350]),

			.SO(gen[8443]),
			.S(gen[8444]),
			.SE(gen[8445]),

			.SELF(gen[8349]),
			.cell_state(gen[8349])
		); 

/******************* CELL 8350 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8350 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8254]),
			.N(gen[8255]),
			.NE(gen[8256]),

			.O(gen[8349]),
			.E(gen[8351]),

			.SO(gen[8444]),
			.S(gen[8445]),
			.SE(gen[8446]),

			.SELF(gen[8350]),
			.cell_state(gen[8350])
		); 

/******************* CELL 8351 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8351 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8255]),
			.N(gen[8256]),
			.NE(gen[8257]),

			.O(gen[8350]),
			.E(gen[8352]),

			.SO(gen[8445]),
			.S(gen[8446]),
			.SE(gen[8447]),

			.SELF(gen[8351]),
			.cell_state(gen[8351])
		); 

/******************* CELL 8352 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8352 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8256]),
			.N(gen[8257]),
			.NE(gen[8258]),

			.O(gen[8351]),
			.E(gen[8353]),

			.SO(gen[8446]),
			.S(gen[8447]),
			.SE(gen[8448]),

			.SELF(gen[8352]),
			.cell_state(gen[8352])
		); 

/******************* CELL 8353 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8353 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8257]),
			.N(gen[8258]),
			.NE(gen[8259]),

			.O(gen[8352]),
			.E(gen[8354]),

			.SO(gen[8447]),
			.S(gen[8448]),
			.SE(gen[8449]),

			.SELF(gen[8353]),
			.cell_state(gen[8353])
		); 

/******************* CELL 8354 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8354 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8258]),
			.N(gen[8259]),
			.NE(gen[8260]),

			.O(gen[8353]),
			.E(gen[8355]),

			.SO(gen[8448]),
			.S(gen[8449]),
			.SE(gen[8450]),

			.SELF(gen[8354]),
			.cell_state(gen[8354])
		); 

/******************* CELL 8355 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8355 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8259]),
			.N(gen[8260]),
			.NE(gen[8261]),

			.O(gen[8354]),
			.E(gen[8356]),

			.SO(gen[8449]),
			.S(gen[8450]),
			.SE(gen[8451]),

			.SELF(gen[8355]),
			.cell_state(gen[8355])
		); 

/******************* CELL 8356 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8356 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8260]),
			.N(gen[8261]),
			.NE(gen[8262]),

			.O(gen[8355]),
			.E(gen[8357]),

			.SO(gen[8450]),
			.S(gen[8451]),
			.SE(gen[8452]),

			.SELF(gen[8356]),
			.cell_state(gen[8356])
		); 

/******************* CELL 8357 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8357 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8261]),
			.N(gen[8262]),
			.NE(gen[8263]),

			.O(gen[8356]),
			.E(gen[8358]),

			.SO(gen[8451]),
			.S(gen[8452]),
			.SE(gen[8453]),

			.SELF(gen[8357]),
			.cell_state(gen[8357])
		); 

/******************* CELL 8358 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8358 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8262]),
			.N(gen[8263]),
			.NE(gen[8264]),

			.O(gen[8357]),
			.E(gen[8359]),

			.SO(gen[8452]),
			.S(gen[8453]),
			.SE(gen[8454]),

			.SELF(gen[8358]),
			.cell_state(gen[8358])
		); 

/******************* CELL 8359 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8359 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8263]),
			.N(gen[8264]),
			.NE(gen[8263]),

			.O(gen[8358]),
			.E(gen[8358]),

			.SO(gen[8453]),
			.S(gen[8454]),
			.SE(gen[8453]),

			.SELF(gen[8359]),
			.cell_state(gen[8359])
		); 

/******************* CELL 8360 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8360 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8266]),
			.N(gen[8265]),
			.NE(gen[8266]),

			.O(gen[8361]),
			.E(gen[8361]),

			.SO(gen[8456]),
			.S(gen[8455]),
			.SE(gen[8456]),

			.SELF(gen[8360]),
			.cell_state(gen[8360])
		); 

/******************* CELL 8361 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8361 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8265]),
			.N(gen[8266]),
			.NE(gen[8267]),

			.O(gen[8360]),
			.E(gen[8362]),

			.SO(gen[8455]),
			.S(gen[8456]),
			.SE(gen[8457]),

			.SELF(gen[8361]),
			.cell_state(gen[8361])
		); 

/******************* CELL 8362 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8362 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8266]),
			.N(gen[8267]),
			.NE(gen[8268]),

			.O(gen[8361]),
			.E(gen[8363]),

			.SO(gen[8456]),
			.S(gen[8457]),
			.SE(gen[8458]),

			.SELF(gen[8362]),
			.cell_state(gen[8362])
		); 

/******************* CELL 8363 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8363 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8267]),
			.N(gen[8268]),
			.NE(gen[8269]),

			.O(gen[8362]),
			.E(gen[8364]),

			.SO(gen[8457]),
			.S(gen[8458]),
			.SE(gen[8459]),

			.SELF(gen[8363]),
			.cell_state(gen[8363])
		); 

/******************* CELL 8364 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8364 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8268]),
			.N(gen[8269]),
			.NE(gen[8270]),

			.O(gen[8363]),
			.E(gen[8365]),

			.SO(gen[8458]),
			.S(gen[8459]),
			.SE(gen[8460]),

			.SELF(gen[8364]),
			.cell_state(gen[8364])
		); 

/******************* CELL 8365 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8365 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8269]),
			.N(gen[8270]),
			.NE(gen[8271]),

			.O(gen[8364]),
			.E(gen[8366]),

			.SO(gen[8459]),
			.S(gen[8460]),
			.SE(gen[8461]),

			.SELF(gen[8365]),
			.cell_state(gen[8365])
		); 

/******************* CELL 8366 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8366 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8270]),
			.N(gen[8271]),
			.NE(gen[8272]),

			.O(gen[8365]),
			.E(gen[8367]),

			.SO(gen[8460]),
			.S(gen[8461]),
			.SE(gen[8462]),

			.SELF(gen[8366]),
			.cell_state(gen[8366])
		); 

/******************* CELL 8367 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8367 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8271]),
			.N(gen[8272]),
			.NE(gen[8273]),

			.O(gen[8366]),
			.E(gen[8368]),

			.SO(gen[8461]),
			.S(gen[8462]),
			.SE(gen[8463]),

			.SELF(gen[8367]),
			.cell_state(gen[8367])
		); 

/******************* CELL 8368 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8368 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8272]),
			.N(gen[8273]),
			.NE(gen[8274]),

			.O(gen[8367]),
			.E(gen[8369]),

			.SO(gen[8462]),
			.S(gen[8463]),
			.SE(gen[8464]),

			.SELF(gen[8368]),
			.cell_state(gen[8368])
		); 

/******************* CELL 8369 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8369 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8273]),
			.N(gen[8274]),
			.NE(gen[8275]),

			.O(gen[8368]),
			.E(gen[8370]),

			.SO(gen[8463]),
			.S(gen[8464]),
			.SE(gen[8465]),

			.SELF(gen[8369]),
			.cell_state(gen[8369])
		); 

/******************* CELL 8370 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8370 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8274]),
			.N(gen[8275]),
			.NE(gen[8276]),

			.O(gen[8369]),
			.E(gen[8371]),

			.SO(gen[8464]),
			.S(gen[8465]),
			.SE(gen[8466]),

			.SELF(gen[8370]),
			.cell_state(gen[8370])
		); 

/******************* CELL 8371 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8371 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8275]),
			.N(gen[8276]),
			.NE(gen[8277]),

			.O(gen[8370]),
			.E(gen[8372]),

			.SO(gen[8465]),
			.S(gen[8466]),
			.SE(gen[8467]),

			.SELF(gen[8371]),
			.cell_state(gen[8371])
		); 

/******************* CELL 8372 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8372 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8276]),
			.N(gen[8277]),
			.NE(gen[8278]),

			.O(gen[8371]),
			.E(gen[8373]),

			.SO(gen[8466]),
			.S(gen[8467]),
			.SE(gen[8468]),

			.SELF(gen[8372]),
			.cell_state(gen[8372])
		); 

/******************* CELL 8373 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8373 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8277]),
			.N(gen[8278]),
			.NE(gen[8279]),

			.O(gen[8372]),
			.E(gen[8374]),

			.SO(gen[8467]),
			.S(gen[8468]),
			.SE(gen[8469]),

			.SELF(gen[8373]),
			.cell_state(gen[8373])
		); 

/******************* CELL 8374 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8374 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8278]),
			.N(gen[8279]),
			.NE(gen[8280]),

			.O(gen[8373]),
			.E(gen[8375]),

			.SO(gen[8468]),
			.S(gen[8469]),
			.SE(gen[8470]),

			.SELF(gen[8374]),
			.cell_state(gen[8374])
		); 

/******************* CELL 8375 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8375 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8279]),
			.N(gen[8280]),
			.NE(gen[8281]),

			.O(gen[8374]),
			.E(gen[8376]),

			.SO(gen[8469]),
			.S(gen[8470]),
			.SE(gen[8471]),

			.SELF(gen[8375]),
			.cell_state(gen[8375])
		); 

/******************* CELL 8376 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8376 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8280]),
			.N(gen[8281]),
			.NE(gen[8282]),

			.O(gen[8375]),
			.E(gen[8377]),

			.SO(gen[8470]),
			.S(gen[8471]),
			.SE(gen[8472]),

			.SELF(gen[8376]),
			.cell_state(gen[8376])
		); 

/******************* CELL 8377 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8377 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8281]),
			.N(gen[8282]),
			.NE(gen[8283]),

			.O(gen[8376]),
			.E(gen[8378]),

			.SO(gen[8471]),
			.S(gen[8472]),
			.SE(gen[8473]),

			.SELF(gen[8377]),
			.cell_state(gen[8377])
		); 

/******************* CELL 8378 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8378 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8282]),
			.N(gen[8283]),
			.NE(gen[8284]),

			.O(gen[8377]),
			.E(gen[8379]),

			.SO(gen[8472]),
			.S(gen[8473]),
			.SE(gen[8474]),

			.SELF(gen[8378]),
			.cell_state(gen[8378])
		); 

/******************* CELL 8379 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8379 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8283]),
			.N(gen[8284]),
			.NE(gen[8285]),

			.O(gen[8378]),
			.E(gen[8380]),

			.SO(gen[8473]),
			.S(gen[8474]),
			.SE(gen[8475]),

			.SELF(gen[8379]),
			.cell_state(gen[8379])
		); 

/******************* CELL 8380 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8380 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8284]),
			.N(gen[8285]),
			.NE(gen[8286]),

			.O(gen[8379]),
			.E(gen[8381]),

			.SO(gen[8474]),
			.S(gen[8475]),
			.SE(gen[8476]),

			.SELF(gen[8380]),
			.cell_state(gen[8380])
		); 

/******************* CELL 8381 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8381 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8285]),
			.N(gen[8286]),
			.NE(gen[8287]),

			.O(gen[8380]),
			.E(gen[8382]),

			.SO(gen[8475]),
			.S(gen[8476]),
			.SE(gen[8477]),

			.SELF(gen[8381]),
			.cell_state(gen[8381])
		); 

/******************* CELL 8382 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8382 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8286]),
			.N(gen[8287]),
			.NE(gen[8288]),

			.O(gen[8381]),
			.E(gen[8383]),

			.SO(gen[8476]),
			.S(gen[8477]),
			.SE(gen[8478]),

			.SELF(gen[8382]),
			.cell_state(gen[8382])
		); 

/******************* CELL 8383 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8383 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8287]),
			.N(gen[8288]),
			.NE(gen[8289]),

			.O(gen[8382]),
			.E(gen[8384]),

			.SO(gen[8477]),
			.S(gen[8478]),
			.SE(gen[8479]),

			.SELF(gen[8383]),
			.cell_state(gen[8383])
		); 

/******************* CELL 8384 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8384 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8288]),
			.N(gen[8289]),
			.NE(gen[8290]),

			.O(gen[8383]),
			.E(gen[8385]),

			.SO(gen[8478]),
			.S(gen[8479]),
			.SE(gen[8480]),

			.SELF(gen[8384]),
			.cell_state(gen[8384])
		); 

/******************* CELL 8385 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8385 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8289]),
			.N(gen[8290]),
			.NE(gen[8291]),

			.O(gen[8384]),
			.E(gen[8386]),

			.SO(gen[8479]),
			.S(gen[8480]),
			.SE(gen[8481]),

			.SELF(gen[8385]),
			.cell_state(gen[8385])
		); 

/******************* CELL 8386 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8386 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8290]),
			.N(gen[8291]),
			.NE(gen[8292]),

			.O(gen[8385]),
			.E(gen[8387]),

			.SO(gen[8480]),
			.S(gen[8481]),
			.SE(gen[8482]),

			.SELF(gen[8386]),
			.cell_state(gen[8386])
		); 

/******************* CELL 8387 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8387 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8291]),
			.N(gen[8292]),
			.NE(gen[8293]),

			.O(gen[8386]),
			.E(gen[8388]),

			.SO(gen[8481]),
			.S(gen[8482]),
			.SE(gen[8483]),

			.SELF(gen[8387]),
			.cell_state(gen[8387])
		); 

/******************* CELL 8388 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8388 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8292]),
			.N(gen[8293]),
			.NE(gen[8294]),

			.O(gen[8387]),
			.E(gen[8389]),

			.SO(gen[8482]),
			.S(gen[8483]),
			.SE(gen[8484]),

			.SELF(gen[8388]),
			.cell_state(gen[8388])
		); 

/******************* CELL 8389 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8389 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8293]),
			.N(gen[8294]),
			.NE(gen[8295]),

			.O(gen[8388]),
			.E(gen[8390]),

			.SO(gen[8483]),
			.S(gen[8484]),
			.SE(gen[8485]),

			.SELF(gen[8389]),
			.cell_state(gen[8389])
		); 

/******************* CELL 8390 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8390 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8294]),
			.N(gen[8295]),
			.NE(gen[8296]),

			.O(gen[8389]),
			.E(gen[8391]),

			.SO(gen[8484]),
			.S(gen[8485]),
			.SE(gen[8486]),

			.SELF(gen[8390]),
			.cell_state(gen[8390])
		); 

/******************* CELL 8391 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8391 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8295]),
			.N(gen[8296]),
			.NE(gen[8297]),

			.O(gen[8390]),
			.E(gen[8392]),

			.SO(gen[8485]),
			.S(gen[8486]),
			.SE(gen[8487]),

			.SELF(gen[8391]),
			.cell_state(gen[8391])
		); 

/******************* CELL 8392 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8392 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8296]),
			.N(gen[8297]),
			.NE(gen[8298]),

			.O(gen[8391]),
			.E(gen[8393]),

			.SO(gen[8486]),
			.S(gen[8487]),
			.SE(gen[8488]),

			.SELF(gen[8392]),
			.cell_state(gen[8392])
		); 

/******************* CELL 8393 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8393 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8297]),
			.N(gen[8298]),
			.NE(gen[8299]),

			.O(gen[8392]),
			.E(gen[8394]),

			.SO(gen[8487]),
			.S(gen[8488]),
			.SE(gen[8489]),

			.SELF(gen[8393]),
			.cell_state(gen[8393])
		); 

/******************* CELL 8394 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8394 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8298]),
			.N(gen[8299]),
			.NE(gen[8300]),

			.O(gen[8393]),
			.E(gen[8395]),

			.SO(gen[8488]),
			.S(gen[8489]),
			.SE(gen[8490]),

			.SELF(gen[8394]),
			.cell_state(gen[8394])
		); 

/******************* CELL 8395 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8395 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8299]),
			.N(gen[8300]),
			.NE(gen[8301]),

			.O(gen[8394]),
			.E(gen[8396]),

			.SO(gen[8489]),
			.S(gen[8490]),
			.SE(gen[8491]),

			.SELF(gen[8395]),
			.cell_state(gen[8395])
		); 

/******************* CELL 8396 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8396 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8300]),
			.N(gen[8301]),
			.NE(gen[8302]),

			.O(gen[8395]),
			.E(gen[8397]),

			.SO(gen[8490]),
			.S(gen[8491]),
			.SE(gen[8492]),

			.SELF(gen[8396]),
			.cell_state(gen[8396])
		); 

/******************* CELL 8397 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8397 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8301]),
			.N(gen[8302]),
			.NE(gen[8303]),

			.O(gen[8396]),
			.E(gen[8398]),

			.SO(gen[8491]),
			.S(gen[8492]),
			.SE(gen[8493]),

			.SELF(gen[8397]),
			.cell_state(gen[8397])
		); 

/******************* CELL 8398 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8398 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8302]),
			.N(gen[8303]),
			.NE(gen[8304]),

			.O(gen[8397]),
			.E(gen[8399]),

			.SO(gen[8492]),
			.S(gen[8493]),
			.SE(gen[8494]),

			.SELF(gen[8398]),
			.cell_state(gen[8398])
		); 

/******************* CELL 8399 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8399 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8303]),
			.N(gen[8304]),
			.NE(gen[8305]),

			.O(gen[8398]),
			.E(gen[8400]),

			.SO(gen[8493]),
			.S(gen[8494]),
			.SE(gen[8495]),

			.SELF(gen[8399]),
			.cell_state(gen[8399])
		); 

/******************* CELL 8400 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8400 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8304]),
			.N(gen[8305]),
			.NE(gen[8306]),

			.O(gen[8399]),
			.E(gen[8401]),

			.SO(gen[8494]),
			.S(gen[8495]),
			.SE(gen[8496]),

			.SELF(gen[8400]),
			.cell_state(gen[8400])
		); 

/******************* CELL 8401 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8401 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8305]),
			.N(gen[8306]),
			.NE(gen[8307]),

			.O(gen[8400]),
			.E(gen[8402]),

			.SO(gen[8495]),
			.S(gen[8496]),
			.SE(gen[8497]),

			.SELF(gen[8401]),
			.cell_state(gen[8401])
		); 

/******************* CELL 8402 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8402 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8306]),
			.N(gen[8307]),
			.NE(gen[8308]),

			.O(gen[8401]),
			.E(gen[8403]),

			.SO(gen[8496]),
			.S(gen[8497]),
			.SE(gen[8498]),

			.SELF(gen[8402]),
			.cell_state(gen[8402])
		); 

/******************* CELL 8403 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8403 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8307]),
			.N(gen[8308]),
			.NE(gen[8309]),

			.O(gen[8402]),
			.E(gen[8404]),

			.SO(gen[8497]),
			.S(gen[8498]),
			.SE(gen[8499]),

			.SELF(gen[8403]),
			.cell_state(gen[8403])
		); 

/******************* CELL 8404 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8404 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8308]),
			.N(gen[8309]),
			.NE(gen[8310]),

			.O(gen[8403]),
			.E(gen[8405]),

			.SO(gen[8498]),
			.S(gen[8499]),
			.SE(gen[8500]),

			.SELF(gen[8404]),
			.cell_state(gen[8404])
		); 

/******************* CELL 8405 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8405 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8309]),
			.N(gen[8310]),
			.NE(gen[8311]),

			.O(gen[8404]),
			.E(gen[8406]),

			.SO(gen[8499]),
			.S(gen[8500]),
			.SE(gen[8501]),

			.SELF(gen[8405]),
			.cell_state(gen[8405])
		); 

/******************* CELL 8406 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8406 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8310]),
			.N(gen[8311]),
			.NE(gen[8312]),

			.O(gen[8405]),
			.E(gen[8407]),

			.SO(gen[8500]),
			.S(gen[8501]),
			.SE(gen[8502]),

			.SELF(gen[8406]),
			.cell_state(gen[8406])
		); 

/******************* CELL 8407 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8407 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8311]),
			.N(gen[8312]),
			.NE(gen[8313]),

			.O(gen[8406]),
			.E(gen[8408]),

			.SO(gen[8501]),
			.S(gen[8502]),
			.SE(gen[8503]),

			.SELF(gen[8407]),
			.cell_state(gen[8407])
		); 

/******************* CELL 8408 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8408 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8312]),
			.N(gen[8313]),
			.NE(gen[8314]),

			.O(gen[8407]),
			.E(gen[8409]),

			.SO(gen[8502]),
			.S(gen[8503]),
			.SE(gen[8504]),

			.SELF(gen[8408]),
			.cell_state(gen[8408])
		); 

/******************* CELL 8409 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8409 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8313]),
			.N(gen[8314]),
			.NE(gen[8315]),

			.O(gen[8408]),
			.E(gen[8410]),

			.SO(gen[8503]),
			.S(gen[8504]),
			.SE(gen[8505]),

			.SELF(gen[8409]),
			.cell_state(gen[8409])
		); 

/******************* CELL 8410 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8410 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8314]),
			.N(gen[8315]),
			.NE(gen[8316]),

			.O(gen[8409]),
			.E(gen[8411]),

			.SO(gen[8504]),
			.S(gen[8505]),
			.SE(gen[8506]),

			.SELF(gen[8410]),
			.cell_state(gen[8410])
		); 

/******************* CELL 8411 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8411 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8315]),
			.N(gen[8316]),
			.NE(gen[8317]),

			.O(gen[8410]),
			.E(gen[8412]),

			.SO(gen[8505]),
			.S(gen[8506]),
			.SE(gen[8507]),

			.SELF(gen[8411]),
			.cell_state(gen[8411])
		); 

/******************* CELL 8412 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8412 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8316]),
			.N(gen[8317]),
			.NE(gen[8318]),

			.O(gen[8411]),
			.E(gen[8413]),

			.SO(gen[8506]),
			.S(gen[8507]),
			.SE(gen[8508]),

			.SELF(gen[8412]),
			.cell_state(gen[8412])
		); 

/******************* CELL 8413 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8413 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8317]),
			.N(gen[8318]),
			.NE(gen[8319]),

			.O(gen[8412]),
			.E(gen[8414]),

			.SO(gen[8507]),
			.S(gen[8508]),
			.SE(gen[8509]),

			.SELF(gen[8413]),
			.cell_state(gen[8413])
		); 

/******************* CELL 8414 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8414 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8318]),
			.N(gen[8319]),
			.NE(gen[8320]),

			.O(gen[8413]),
			.E(gen[8415]),

			.SO(gen[8508]),
			.S(gen[8509]),
			.SE(gen[8510]),

			.SELF(gen[8414]),
			.cell_state(gen[8414])
		); 

/******************* CELL 8415 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8415 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8319]),
			.N(gen[8320]),
			.NE(gen[8321]),

			.O(gen[8414]),
			.E(gen[8416]),

			.SO(gen[8509]),
			.S(gen[8510]),
			.SE(gen[8511]),

			.SELF(gen[8415]),
			.cell_state(gen[8415])
		); 

/******************* CELL 8416 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8416 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8320]),
			.N(gen[8321]),
			.NE(gen[8322]),

			.O(gen[8415]),
			.E(gen[8417]),

			.SO(gen[8510]),
			.S(gen[8511]),
			.SE(gen[8512]),

			.SELF(gen[8416]),
			.cell_state(gen[8416])
		); 

/******************* CELL 8417 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8417 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8321]),
			.N(gen[8322]),
			.NE(gen[8323]),

			.O(gen[8416]),
			.E(gen[8418]),

			.SO(gen[8511]),
			.S(gen[8512]),
			.SE(gen[8513]),

			.SELF(gen[8417]),
			.cell_state(gen[8417])
		); 

/******************* CELL 8418 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8418 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8322]),
			.N(gen[8323]),
			.NE(gen[8324]),

			.O(gen[8417]),
			.E(gen[8419]),

			.SO(gen[8512]),
			.S(gen[8513]),
			.SE(gen[8514]),

			.SELF(gen[8418]),
			.cell_state(gen[8418])
		); 

/******************* CELL 8419 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8419 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8323]),
			.N(gen[8324]),
			.NE(gen[8325]),

			.O(gen[8418]),
			.E(gen[8420]),

			.SO(gen[8513]),
			.S(gen[8514]),
			.SE(gen[8515]),

			.SELF(gen[8419]),
			.cell_state(gen[8419])
		); 

/******************* CELL 8420 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8420 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8324]),
			.N(gen[8325]),
			.NE(gen[8326]),

			.O(gen[8419]),
			.E(gen[8421]),

			.SO(gen[8514]),
			.S(gen[8515]),
			.SE(gen[8516]),

			.SELF(gen[8420]),
			.cell_state(gen[8420])
		); 

/******************* CELL 8421 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8421 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8325]),
			.N(gen[8326]),
			.NE(gen[8327]),

			.O(gen[8420]),
			.E(gen[8422]),

			.SO(gen[8515]),
			.S(gen[8516]),
			.SE(gen[8517]),

			.SELF(gen[8421]),
			.cell_state(gen[8421])
		); 

/******************* CELL 8422 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8422 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8326]),
			.N(gen[8327]),
			.NE(gen[8328]),

			.O(gen[8421]),
			.E(gen[8423]),

			.SO(gen[8516]),
			.S(gen[8517]),
			.SE(gen[8518]),

			.SELF(gen[8422]),
			.cell_state(gen[8422])
		); 

/******************* CELL 8423 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8423 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8327]),
			.N(gen[8328]),
			.NE(gen[8329]),

			.O(gen[8422]),
			.E(gen[8424]),

			.SO(gen[8517]),
			.S(gen[8518]),
			.SE(gen[8519]),

			.SELF(gen[8423]),
			.cell_state(gen[8423])
		); 

/******************* CELL 8424 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8424 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8328]),
			.N(gen[8329]),
			.NE(gen[8330]),

			.O(gen[8423]),
			.E(gen[8425]),

			.SO(gen[8518]),
			.S(gen[8519]),
			.SE(gen[8520]),

			.SELF(gen[8424]),
			.cell_state(gen[8424])
		); 

/******************* CELL 8425 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8425 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8329]),
			.N(gen[8330]),
			.NE(gen[8331]),

			.O(gen[8424]),
			.E(gen[8426]),

			.SO(gen[8519]),
			.S(gen[8520]),
			.SE(gen[8521]),

			.SELF(gen[8425]),
			.cell_state(gen[8425])
		); 

/******************* CELL 8426 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8426 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8330]),
			.N(gen[8331]),
			.NE(gen[8332]),

			.O(gen[8425]),
			.E(gen[8427]),

			.SO(gen[8520]),
			.S(gen[8521]),
			.SE(gen[8522]),

			.SELF(gen[8426]),
			.cell_state(gen[8426])
		); 

/******************* CELL 8427 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8427 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8331]),
			.N(gen[8332]),
			.NE(gen[8333]),

			.O(gen[8426]),
			.E(gen[8428]),

			.SO(gen[8521]),
			.S(gen[8522]),
			.SE(gen[8523]),

			.SELF(gen[8427]),
			.cell_state(gen[8427])
		); 

/******************* CELL 8428 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8428 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8332]),
			.N(gen[8333]),
			.NE(gen[8334]),

			.O(gen[8427]),
			.E(gen[8429]),

			.SO(gen[8522]),
			.S(gen[8523]),
			.SE(gen[8524]),

			.SELF(gen[8428]),
			.cell_state(gen[8428])
		); 

/******************* CELL 8429 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8429 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8333]),
			.N(gen[8334]),
			.NE(gen[8335]),

			.O(gen[8428]),
			.E(gen[8430]),

			.SO(gen[8523]),
			.S(gen[8524]),
			.SE(gen[8525]),

			.SELF(gen[8429]),
			.cell_state(gen[8429])
		); 

/******************* CELL 8430 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8430 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8334]),
			.N(gen[8335]),
			.NE(gen[8336]),

			.O(gen[8429]),
			.E(gen[8431]),

			.SO(gen[8524]),
			.S(gen[8525]),
			.SE(gen[8526]),

			.SELF(gen[8430]),
			.cell_state(gen[8430])
		); 

/******************* CELL 8431 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8431 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8335]),
			.N(gen[8336]),
			.NE(gen[8337]),

			.O(gen[8430]),
			.E(gen[8432]),

			.SO(gen[8525]),
			.S(gen[8526]),
			.SE(gen[8527]),

			.SELF(gen[8431]),
			.cell_state(gen[8431])
		); 

/******************* CELL 8432 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8432 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8336]),
			.N(gen[8337]),
			.NE(gen[8338]),

			.O(gen[8431]),
			.E(gen[8433]),

			.SO(gen[8526]),
			.S(gen[8527]),
			.SE(gen[8528]),

			.SELF(gen[8432]),
			.cell_state(gen[8432])
		); 

/******************* CELL 8433 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8433 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8337]),
			.N(gen[8338]),
			.NE(gen[8339]),

			.O(gen[8432]),
			.E(gen[8434]),

			.SO(gen[8527]),
			.S(gen[8528]),
			.SE(gen[8529]),

			.SELF(gen[8433]),
			.cell_state(gen[8433])
		); 

/******************* CELL 8434 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8434 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8338]),
			.N(gen[8339]),
			.NE(gen[8340]),

			.O(gen[8433]),
			.E(gen[8435]),

			.SO(gen[8528]),
			.S(gen[8529]),
			.SE(gen[8530]),

			.SELF(gen[8434]),
			.cell_state(gen[8434])
		); 

/******************* CELL 8435 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8435 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8339]),
			.N(gen[8340]),
			.NE(gen[8341]),

			.O(gen[8434]),
			.E(gen[8436]),

			.SO(gen[8529]),
			.S(gen[8530]),
			.SE(gen[8531]),

			.SELF(gen[8435]),
			.cell_state(gen[8435])
		); 

/******************* CELL 8436 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8436 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8340]),
			.N(gen[8341]),
			.NE(gen[8342]),

			.O(gen[8435]),
			.E(gen[8437]),

			.SO(gen[8530]),
			.S(gen[8531]),
			.SE(gen[8532]),

			.SELF(gen[8436]),
			.cell_state(gen[8436])
		); 

/******************* CELL 8437 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8437 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8341]),
			.N(gen[8342]),
			.NE(gen[8343]),

			.O(gen[8436]),
			.E(gen[8438]),

			.SO(gen[8531]),
			.S(gen[8532]),
			.SE(gen[8533]),

			.SELF(gen[8437]),
			.cell_state(gen[8437])
		); 

/******************* CELL 8438 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8438 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8342]),
			.N(gen[8343]),
			.NE(gen[8344]),

			.O(gen[8437]),
			.E(gen[8439]),

			.SO(gen[8532]),
			.S(gen[8533]),
			.SE(gen[8534]),

			.SELF(gen[8438]),
			.cell_state(gen[8438])
		); 

/******************* CELL 8439 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8439 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8343]),
			.N(gen[8344]),
			.NE(gen[8345]),

			.O(gen[8438]),
			.E(gen[8440]),

			.SO(gen[8533]),
			.S(gen[8534]),
			.SE(gen[8535]),

			.SELF(gen[8439]),
			.cell_state(gen[8439])
		); 

/******************* CELL 8440 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8440 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8344]),
			.N(gen[8345]),
			.NE(gen[8346]),

			.O(gen[8439]),
			.E(gen[8441]),

			.SO(gen[8534]),
			.S(gen[8535]),
			.SE(gen[8536]),

			.SELF(gen[8440]),
			.cell_state(gen[8440])
		); 

/******************* CELL 8441 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8441 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8345]),
			.N(gen[8346]),
			.NE(gen[8347]),

			.O(gen[8440]),
			.E(gen[8442]),

			.SO(gen[8535]),
			.S(gen[8536]),
			.SE(gen[8537]),

			.SELF(gen[8441]),
			.cell_state(gen[8441])
		); 

/******************* CELL 8442 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8442 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8346]),
			.N(gen[8347]),
			.NE(gen[8348]),

			.O(gen[8441]),
			.E(gen[8443]),

			.SO(gen[8536]),
			.S(gen[8537]),
			.SE(gen[8538]),

			.SELF(gen[8442]),
			.cell_state(gen[8442])
		); 

/******************* CELL 8443 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8443 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8347]),
			.N(gen[8348]),
			.NE(gen[8349]),

			.O(gen[8442]),
			.E(gen[8444]),

			.SO(gen[8537]),
			.S(gen[8538]),
			.SE(gen[8539]),

			.SELF(gen[8443]),
			.cell_state(gen[8443])
		); 

/******************* CELL 8444 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8444 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8348]),
			.N(gen[8349]),
			.NE(gen[8350]),

			.O(gen[8443]),
			.E(gen[8445]),

			.SO(gen[8538]),
			.S(gen[8539]),
			.SE(gen[8540]),

			.SELF(gen[8444]),
			.cell_state(gen[8444])
		); 

/******************* CELL 8445 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8445 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8349]),
			.N(gen[8350]),
			.NE(gen[8351]),

			.O(gen[8444]),
			.E(gen[8446]),

			.SO(gen[8539]),
			.S(gen[8540]),
			.SE(gen[8541]),

			.SELF(gen[8445]),
			.cell_state(gen[8445])
		); 

/******************* CELL 8446 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8446 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8350]),
			.N(gen[8351]),
			.NE(gen[8352]),

			.O(gen[8445]),
			.E(gen[8447]),

			.SO(gen[8540]),
			.S(gen[8541]),
			.SE(gen[8542]),

			.SELF(gen[8446]),
			.cell_state(gen[8446])
		); 

/******************* CELL 8447 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8447 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8351]),
			.N(gen[8352]),
			.NE(gen[8353]),

			.O(gen[8446]),
			.E(gen[8448]),

			.SO(gen[8541]),
			.S(gen[8542]),
			.SE(gen[8543]),

			.SELF(gen[8447]),
			.cell_state(gen[8447])
		); 

/******************* CELL 8448 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8448 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8352]),
			.N(gen[8353]),
			.NE(gen[8354]),

			.O(gen[8447]),
			.E(gen[8449]),

			.SO(gen[8542]),
			.S(gen[8543]),
			.SE(gen[8544]),

			.SELF(gen[8448]),
			.cell_state(gen[8448])
		); 

/******************* CELL 8449 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8449 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8353]),
			.N(gen[8354]),
			.NE(gen[8355]),

			.O(gen[8448]),
			.E(gen[8450]),

			.SO(gen[8543]),
			.S(gen[8544]),
			.SE(gen[8545]),

			.SELF(gen[8449]),
			.cell_state(gen[8449])
		); 

/******************* CELL 8450 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8450 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8354]),
			.N(gen[8355]),
			.NE(gen[8356]),

			.O(gen[8449]),
			.E(gen[8451]),

			.SO(gen[8544]),
			.S(gen[8545]),
			.SE(gen[8546]),

			.SELF(gen[8450]),
			.cell_state(gen[8450])
		); 

/******************* CELL 8451 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8451 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8355]),
			.N(gen[8356]),
			.NE(gen[8357]),

			.O(gen[8450]),
			.E(gen[8452]),

			.SO(gen[8545]),
			.S(gen[8546]),
			.SE(gen[8547]),

			.SELF(gen[8451]),
			.cell_state(gen[8451])
		); 

/******************* CELL 8452 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8452 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8356]),
			.N(gen[8357]),
			.NE(gen[8358]),

			.O(gen[8451]),
			.E(gen[8453]),

			.SO(gen[8546]),
			.S(gen[8547]),
			.SE(gen[8548]),

			.SELF(gen[8452]),
			.cell_state(gen[8452])
		); 

/******************* CELL 8453 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8453 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8357]),
			.N(gen[8358]),
			.NE(gen[8359]),

			.O(gen[8452]),
			.E(gen[8454]),

			.SO(gen[8547]),
			.S(gen[8548]),
			.SE(gen[8549]),

			.SELF(gen[8453]),
			.cell_state(gen[8453])
		); 

/******************* CELL 8454 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8454 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8358]),
			.N(gen[8359]),
			.NE(gen[8358]),

			.O(gen[8453]),
			.E(gen[8453]),

			.SO(gen[8548]),
			.S(gen[8549]),
			.SE(gen[8548]),

			.SELF(gen[8454]),
			.cell_state(gen[8454])
		); 

/******************* CELL 8455 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8455 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8361]),
			.N(gen[8360]),
			.NE(gen[8361]),

			.O(gen[8456]),
			.E(gen[8456]),

			.SO(gen[8551]),
			.S(gen[8550]),
			.SE(gen[8551]),

			.SELF(gen[8455]),
			.cell_state(gen[8455])
		); 

/******************* CELL 8456 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8456 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8360]),
			.N(gen[8361]),
			.NE(gen[8362]),

			.O(gen[8455]),
			.E(gen[8457]),

			.SO(gen[8550]),
			.S(gen[8551]),
			.SE(gen[8552]),

			.SELF(gen[8456]),
			.cell_state(gen[8456])
		); 

/******************* CELL 8457 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8457 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8361]),
			.N(gen[8362]),
			.NE(gen[8363]),

			.O(gen[8456]),
			.E(gen[8458]),

			.SO(gen[8551]),
			.S(gen[8552]),
			.SE(gen[8553]),

			.SELF(gen[8457]),
			.cell_state(gen[8457])
		); 

/******************* CELL 8458 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8458 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8362]),
			.N(gen[8363]),
			.NE(gen[8364]),

			.O(gen[8457]),
			.E(gen[8459]),

			.SO(gen[8552]),
			.S(gen[8553]),
			.SE(gen[8554]),

			.SELF(gen[8458]),
			.cell_state(gen[8458])
		); 

/******************* CELL 8459 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8459 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8363]),
			.N(gen[8364]),
			.NE(gen[8365]),

			.O(gen[8458]),
			.E(gen[8460]),

			.SO(gen[8553]),
			.S(gen[8554]),
			.SE(gen[8555]),

			.SELF(gen[8459]),
			.cell_state(gen[8459])
		); 

/******************* CELL 8460 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8460 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8364]),
			.N(gen[8365]),
			.NE(gen[8366]),

			.O(gen[8459]),
			.E(gen[8461]),

			.SO(gen[8554]),
			.S(gen[8555]),
			.SE(gen[8556]),

			.SELF(gen[8460]),
			.cell_state(gen[8460])
		); 

/******************* CELL 8461 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8461 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8365]),
			.N(gen[8366]),
			.NE(gen[8367]),

			.O(gen[8460]),
			.E(gen[8462]),

			.SO(gen[8555]),
			.S(gen[8556]),
			.SE(gen[8557]),

			.SELF(gen[8461]),
			.cell_state(gen[8461])
		); 

/******************* CELL 8462 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8462 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8366]),
			.N(gen[8367]),
			.NE(gen[8368]),

			.O(gen[8461]),
			.E(gen[8463]),

			.SO(gen[8556]),
			.S(gen[8557]),
			.SE(gen[8558]),

			.SELF(gen[8462]),
			.cell_state(gen[8462])
		); 

/******************* CELL 8463 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8463 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8367]),
			.N(gen[8368]),
			.NE(gen[8369]),

			.O(gen[8462]),
			.E(gen[8464]),

			.SO(gen[8557]),
			.S(gen[8558]),
			.SE(gen[8559]),

			.SELF(gen[8463]),
			.cell_state(gen[8463])
		); 

/******************* CELL 8464 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8464 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8368]),
			.N(gen[8369]),
			.NE(gen[8370]),

			.O(gen[8463]),
			.E(gen[8465]),

			.SO(gen[8558]),
			.S(gen[8559]),
			.SE(gen[8560]),

			.SELF(gen[8464]),
			.cell_state(gen[8464])
		); 

/******************* CELL 8465 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8465 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8369]),
			.N(gen[8370]),
			.NE(gen[8371]),

			.O(gen[8464]),
			.E(gen[8466]),

			.SO(gen[8559]),
			.S(gen[8560]),
			.SE(gen[8561]),

			.SELF(gen[8465]),
			.cell_state(gen[8465])
		); 

/******************* CELL 8466 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8466 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8370]),
			.N(gen[8371]),
			.NE(gen[8372]),

			.O(gen[8465]),
			.E(gen[8467]),

			.SO(gen[8560]),
			.S(gen[8561]),
			.SE(gen[8562]),

			.SELF(gen[8466]),
			.cell_state(gen[8466])
		); 

/******************* CELL 8467 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8467 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8371]),
			.N(gen[8372]),
			.NE(gen[8373]),

			.O(gen[8466]),
			.E(gen[8468]),

			.SO(gen[8561]),
			.S(gen[8562]),
			.SE(gen[8563]),

			.SELF(gen[8467]),
			.cell_state(gen[8467])
		); 

/******************* CELL 8468 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8468 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8372]),
			.N(gen[8373]),
			.NE(gen[8374]),

			.O(gen[8467]),
			.E(gen[8469]),

			.SO(gen[8562]),
			.S(gen[8563]),
			.SE(gen[8564]),

			.SELF(gen[8468]),
			.cell_state(gen[8468])
		); 

/******************* CELL 8469 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8469 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8373]),
			.N(gen[8374]),
			.NE(gen[8375]),

			.O(gen[8468]),
			.E(gen[8470]),

			.SO(gen[8563]),
			.S(gen[8564]),
			.SE(gen[8565]),

			.SELF(gen[8469]),
			.cell_state(gen[8469])
		); 

/******************* CELL 8470 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8470 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8374]),
			.N(gen[8375]),
			.NE(gen[8376]),

			.O(gen[8469]),
			.E(gen[8471]),

			.SO(gen[8564]),
			.S(gen[8565]),
			.SE(gen[8566]),

			.SELF(gen[8470]),
			.cell_state(gen[8470])
		); 

/******************* CELL 8471 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8471 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8375]),
			.N(gen[8376]),
			.NE(gen[8377]),

			.O(gen[8470]),
			.E(gen[8472]),

			.SO(gen[8565]),
			.S(gen[8566]),
			.SE(gen[8567]),

			.SELF(gen[8471]),
			.cell_state(gen[8471])
		); 

/******************* CELL 8472 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8472 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8376]),
			.N(gen[8377]),
			.NE(gen[8378]),

			.O(gen[8471]),
			.E(gen[8473]),

			.SO(gen[8566]),
			.S(gen[8567]),
			.SE(gen[8568]),

			.SELF(gen[8472]),
			.cell_state(gen[8472])
		); 

/******************* CELL 8473 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8473 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8377]),
			.N(gen[8378]),
			.NE(gen[8379]),

			.O(gen[8472]),
			.E(gen[8474]),

			.SO(gen[8567]),
			.S(gen[8568]),
			.SE(gen[8569]),

			.SELF(gen[8473]),
			.cell_state(gen[8473])
		); 

/******************* CELL 8474 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8474 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8378]),
			.N(gen[8379]),
			.NE(gen[8380]),

			.O(gen[8473]),
			.E(gen[8475]),

			.SO(gen[8568]),
			.S(gen[8569]),
			.SE(gen[8570]),

			.SELF(gen[8474]),
			.cell_state(gen[8474])
		); 

/******************* CELL 8475 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8475 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8379]),
			.N(gen[8380]),
			.NE(gen[8381]),

			.O(gen[8474]),
			.E(gen[8476]),

			.SO(gen[8569]),
			.S(gen[8570]),
			.SE(gen[8571]),

			.SELF(gen[8475]),
			.cell_state(gen[8475])
		); 

/******************* CELL 8476 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8476 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8380]),
			.N(gen[8381]),
			.NE(gen[8382]),

			.O(gen[8475]),
			.E(gen[8477]),

			.SO(gen[8570]),
			.S(gen[8571]),
			.SE(gen[8572]),

			.SELF(gen[8476]),
			.cell_state(gen[8476])
		); 

/******************* CELL 8477 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8477 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8381]),
			.N(gen[8382]),
			.NE(gen[8383]),

			.O(gen[8476]),
			.E(gen[8478]),

			.SO(gen[8571]),
			.S(gen[8572]),
			.SE(gen[8573]),

			.SELF(gen[8477]),
			.cell_state(gen[8477])
		); 

/******************* CELL 8478 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8478 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8382]),
			.N(gen[8383]),
			.NE(gen[8384]),

			.O(gen[8477]),
			.E(gen[8479]),

			.SO(gen[8572]),
			.S(gen[8573]),
			.SE(gen[8574]),

			.SELF(gen[8478]),
			.cell_state(gen[8478])
		); 

/******************* CELL 8479 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8479 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8383]),
			.N(gen[8384]),
			.NE(gen[8385]),

			.O(gen[8478]),
			.E(gen[8480]),

			.SO(gen[8573]),
			.S(gen[8574]),
			.SE(gen[8575]),

			.SELF(gen[8479]),
			.cell_state(gen[8479])
		); 

/******************* CELL 8480 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8480 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8384]),
			.N(gen[8385]),
			.NE(gen[8386]),

			.O(gen[8479]),
			.E(gen[8481]),

			.SO(gen[8574]),
			.S(gen[8575]),
			.SE(gen[8576]),

			.SELF(gen[8480]),
			.cell_state(gen[8480])
		); 

/******************* CELL 8481 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8481 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8385]),
			.N(gen[8386]),
			.NE(gen[8387]),

			.O(gen[8480]),
			.E(gen[8482]),

			.SO(gen[8575]),
			.S(gen[8576]),
			.SE(gen[8577]),

			.SELF(gen[8481]),
			.cell_state(gen[8481])
		); 

/******************* CELL 8482 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8482 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8386]),
			.N(gen[8387]),
			.NE(gen[8388]),

			.O(gen[8481]),
			.E(gen[8483]),

			.SO(gen[8576]),
			.S(gen[8577]),
			.SE(gen[8578]),

			.SELF(gen[8482]),
			.cell_state(gen[8482])
		); 

/******************* CELL 8483 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8483 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8387]),
			.N(gen[8388]),
			.NE(gen[8389]),

			.O(gen[8482]),
			.E(gen[8484]),

			.SO(gen[8577]),
			.S(gen[8578]),
			.SE(gen[8579]),

			.SELF(gen[8483]),
			.cell_state(gen[8483])
		); 

/******************* CELL 8484 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8484 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8388]),
			.N(gen[8389]),
			.NE(gen[8390]),

			.O(gen[8483]),
			.E(gen[8485]),

			.SO(gen[8578]),
			.S(gen[8579]),
			.SE(gen[8580]),

			.SELF(gen[8484]),
			.cell_state(gen[8484])
		); 

/******************* CELL 8485 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8485 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8389]),
			.N(gen[8390]),
			.NE(gen[8391]),

			.O(gen[8484]),
			.E(gen[8486]),

			.SO(gen[8579]),
			.S(gen[8580]),
			.SE(gen[8581]),

			.SELF(gen[8485]),
			.cell_state(gen[8485])
		); 

/******************* CELL 8486 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8486 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8390]),
			.N(gen[8391]),
			.NE(gen[8392]),

			.O(gen[8485]),
			.E(gen[8487]),

			.SO(gen[8580]),
			.S(gen[8581]),
			.SE(gen[8582]),

			.SELF(gen[8486]),
			.cell_state(gen[8486])
		); 

/******************* CELL 8487 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8487 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8391]),
			.N(gen[8392]),
			.NE(gen[8393]),

			.O(gen[8486]),
			.E(gen[8488]),

			.SO(gen[8581]),
			.S(gen[8582]),
			.SE(gen[8583]),

			.SELF(gen[8487]),
			.cell_state(gen[8487])
		); 

/******************* CELL 8488 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8488 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8392]),
			.N(gen[8393]),
			.NE(gen[8394]),

			.O(gen[8487]),
			.E(gen[8489]),

			.SO(gen[8582]),
			.S(gen[8583]),
			.SE(gen[8584]),

			.SELF(gen[8488]),
			.cell_state(gen[8488])
		); 

/******************* CELL 8489 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8489 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8393]),
			.N(gen[8394]),
			.NE(gen[8395]),

			.O(gen[8488]),
			.E(gen[8490]),

			.SO(gen[8583]),
			.S(gen[8584]),
			.SE(gen[8585]),

			.SELF(gen[8489]),
			.cell_state(gen[8489])
		); 

/******************* CELL 8490 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8490 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8394]),
			.N(gen[8395]),
			.NE(gen[8396]),

			.O(gen[8489]),
			.E(gen[8491]),

			.SO(gen[8584]),
			.S(gen[8585]),
			.SE(gen[8586]),

			.SELF(gen[8490]),
			.cell_state(gen[8490])
		); 

/******************* CELL 8491 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8491 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8395]),
			.N(gen[8396]),
			.NE(gen[8397]),

			.O(gen[8490]),
			.E(gen[8492]),

			.SO(gen[8585]),
			.S(gen[8586]),
			.SE(gen[8587]),

			.SELF(gen[8491]),
			.cell_state(gen[8491])
		); 

/******************* CELL 8492 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8492 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8396]),
			.N(gen[8397]),
			.NE(gen[8398]),

			.O(gen[8491]),
			.E(gen[8493]),

			.SO(gen[8586]),
			.S(gen[8587]),
			.SE(gen[8588]),

			.SELF(gen[8492]),
			.cell_state(gen[8492])
		); 

/******************* CELL 8493 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8493 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8397]),
			.N(gen[8398]),
			.NE(gen[8399]),

			.O(gen[8492]),
			.E(gen[8494]),

			.SO(gen[8587]),
			.S(gen[8588]),
			.SE(gen[8589]),

			.SELF(gen[8493]),
			.cell_state(gen[8493])
		); 

/******************* CELL 8494 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8494 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8398]),
			.N(gen[8399]),
			.NE(gen[8400]),

			.O(gen[8493]),
			.E(gen[8495]),

			.SO(gen[8588]),
			.S(gen[8589]),
			.SE(gen[8590]),

			.SELF(gen[8494]),
			.cell_state(gen[8494])
		); 

/******************* CELL 8495 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8495 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8399]),
			.N(gen[8400]),
			.NE(gen[8401]),

			.O(gen[8494]),
			.E(gen[8496]),

			.SO(gen[8589]),
			.S(gen[8590]),
			.SE(gen[8591]),

			.SELF(gen[8495]),
			.cell_state(gen[8495])
		); 

/******************* CELL 8496 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8496 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8400]),
			.N(gen[8401]),
			.NE(gen[8402]),

			.O(gen[8495]),
			.E(gen[8497]),

			.SO(gen[8590]),
			.S(gen[8591]),
			.SE(gen[8592]),

			.SELF(gen[8496]),
			.cell_state(gen[8496])
		); 

/******************* CELL 8497 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8497 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8401]),
			.N(gen[8402]),
			.NE(gen[8403]),

			.O(gen[8496]),
			.E(gen[8498]),

			.SO(gen[8591]),
			.S(gen[8592]),
			.SE(gen[8593]),

			.SELF(gen[8497]),
			.cell_state(gen[8497])
		); 

/******************* CELL 8498 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8498 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8402]),
			.N(gen[8403]),
			.NE(gen[8404]),

			.O(gen[8497]),
			.E(gen[8499]),

			.SO(gen[8592]),
			.S(gen[8593]),
			.SE(gen[8594]),

			.SELF(gen[8498]),
			.cell_state(gen[8498])
		); 

/******************* CELL 8499 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8499 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8403]),
			.N(gen[8404]),
			.NE(gen[8405]),

			.O(gen[8498]),
			.E(gen[8500]),

			.SO(gen[8593]),
			.S(gen[8594]),
			.SE(gen[8595]),

			.SELF(gen[8499]),
			.cell_state(gen[8499])
		); 

/******************* CELL 8500 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8500 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8404]),
			.N(gen[8405]),
			.NE(gen[8406]),

			.O(gen[8499]),
			.E(gen[8501]),

			.SO(gen[8594]),
			.S(gen[8595]),
			.SE(gen[8596]),

			.SELF(gen[8500]),
			.cell_state(gen[8500])
		); 

/******************* CELL 8501 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8501 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8405]),
			.N(gen[8406]),
			.NE(gen[8407]),

			.O(gen[8500]),
			.E(gen[8502]),

			.SO(gen[8595]),
			.S(gen[8596]),
			.SE(gen[8597]),

			.SELF(gen[8501]),
			.cell_state(gen[8501])
		); 

/******************* CELL 8502 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8502 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8406]),
			.N(gen[8407]),
			.NE(gen[8408]),

			.O(gen[8501]),
			.E(gen[8503]),

			.SO(gen[8596]),
			.S(gen[8597]),
			.SE(gen[8598]),

			.SELF(gen[8502]),
			.cell_state(gen[8502])
		); 

/******************* CELL 8503 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8503 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8407]),
			.N(gen[8408]),
			.NE(gen[8409]),

			.O(gen[8502]),
			.E(gen[8504]),

			.SO(gen[8597]),
			.S(gen[8598]),
			.SE(gen[8599]),

			.SELF(gen[8503]),
			.cell_state(gen[8503])
		); 

/******************* CELL 8504 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8504 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8408]),
			.N(gen[8409]),
			.NE(gen[8410]),

			.O(gen[8503]),
			.E(gen[8505]),

			.SO(gen[8598]),
			.S(gen[8599]),
			.SE(gen[8600]),

			.SELF(gen[8504]),
			.cell_state(gen[8504])
		); 

/******************* CELL 8505 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8505 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8409]),
			.N(gen[8410]),
			.NE(gen[8411]),

			.O(gen[8504]),
			.E(gen[8506]),

			.SO(gen[8599]),
			.S(gen[8600]),
			.SE(gen[8601]),

			.SELF(gen[8505]),
			.cell_state(gen[8505])
		); 

/******************* CELL 8506 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8506 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8410]),
			.N(gen[8411]),
			.NE(gen[8412]),

			.O(gen[8505]),
			.E(gen[8507]),

			.SO(gen[8600]),
			.S(gen[8601]),
			.SE(gen[8602]),

			.SELF(gen[8506]),
			.cell_state(gen[8506])
		); 

/******************* CELL 8507 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8507 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8411]),
			.N(gen[8412]),
			.NE(gen[8413]),

			.O(gen[8506]),
			.E(gen[8508]),

			.SO(gen[8601]),
			.S(gen[8602]),
			.SE(gen[8603]),

			.SELF(gen[8507]),
			.cell_state(gen[8507])
		); 

/******************* CELL 8508 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8508 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8412]),
			.N(gen[8413]),
			.NE(gen[8414]),

			.O(gen[8507]),
			.E(gen[8509]),

			.SO(gen[8602]),
			.S(gen[8603]),
			.SE(gen[8604]),

			.SELF(gen[8508]),
			.cell_state(gen[8508])
		); 

/******************* CELL 8509 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8509 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8413]),
			.N(gen[8414]),
			.NE(gen[8415]),

			.O(gen[8508]),
			.E(gen[8510]),

			.SO(gen[8603]),
			.S(gen[8604]),
			.SE(gen[8605]),

			.SELF(gen[8509]),
			.cell_state(gen[8509])
		); 

/******************* CELL 8510 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8510 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8414]),
			.N(gen[8415]),
			.NE(gen[8416]),

			.O(gen[8509]),
			.E(gen[8511]),

			.SO(gen[8604]),
			.S(gen[8605]),
			.SE(gen[8606]),

			.SELF(gen[8510]),
			.cell_state(gen[8510])
		); 

/******************* CELL 8511 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8511 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8415]),
			.N(gen[8416]),
			.NE(gen[8417]),

			.O(gen[8510]),
			.E(gen[8512]),

			.SO(gen[8605]),
			.S(gen[8606]),
			.SE(gen[8607]),

			.SELF(gen[8511]),
			.cell_state(gen[8511])
		); 

/******************* CELL 8512 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8512 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8416]),
			.N(gen[8417]),
			.NE(gen[8418]),

			.O(gen[8511]),
			.E(gen[8513]),

			.SO(gen[8606]),
			.S(gen[8607]),
			.SE(gen[8608]),

			.SELF(gen[8512]),
			.cell_state(gen[8512])
		); 

/******************* CELL 8513 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8513 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8417]),
			.N(gen[8418]),
			.NE(gen[8419]),

			.O(gen[8512]),
			.E(gen[8514]),

			.SO(gen[8607]),
			.S(gen[8608]),
			.SE(gen[8609]),

			.SELF(gen[8513]),
			.cell_state(gen[8513])
		); 

/******************* CELL 8514 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8514 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8418]),
			.N(gen[8419]),
			.NE(gen[8420]),

			.O(gen[8513]),
			.E(gen[8515]),

			.SO(gen[8608]),
			.S(gen[8609]),
			.SE(gen[8610]),

			.SELF(gen[8514]),
			.cell_state(gen[8514])
		); 

/******************* CELL 8515 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8515 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8419]),
			.N(gen[8420]),
			.NE(gen[8421]),

			.O(gen[8514]),
			.E(gen[8516]),

			.SO(gen[8609]),
			.S(gen[8610]),
			.SE(gen[8611]),

			.SELF(gen[8515]),
			.cell_state(gen[8515])
		); 

/******************* CELL 8516 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8516 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8420]),
			.N(gen[8421]),
			.NE(gen[8422]),

			.O(gen[8515]),
			.E(gen[8517]),

			.SO(gen[8610]),
			.S(gen[8611]),
			.SE(gen[8612]),

			.SELF(gen[8516]),
			.cell_state(gen[8516])
		); 

/******************* CELL 8517 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8517 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8421]),
			.N(gen[8422]),
			.NE(gen[8423]),

			.O(gen[8516]),
			.E(gen[8518]),

			.SO(gen[8611]),
			.S(gen[8612]),
			.SE(gen[8613]),

			.SELF(gen[8517]),
			.cell_state(gen[8517])
		); 

/******************* CELL 8518 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8518 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8422]),
			.N(gen[8423]),
			.NE(gen[8424]),

			.O(gen[8517]),
			.E(gen[8519]),

			.SO(gen[8612]),
			.S(gen[8613]),
			.SE(gen[8614]),

			.SELF(gen[8518]),
			.cell_state(gen[8518])
		); 

/******************* CELL 8519 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8519 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8423]),
			.N(gen[8424]),
			.NE(gen[8425]),

			.O(gen[8518]),
			.E(gen[8520]),

			.SO(gen[8613]),
			.S(gen[8614]),
			.SE(gen[8615]),

			.SELF(gen[8519]),
			.cell_state(gen[8519])
		); 

/******************* CELL 8520 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8520 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8424]),
			.N(gen[8425]),
			.NE(gen[8426]),

			.O(gen[8519]),
			.E(gen[8521]),

			.SO(gen[8614]),
			.S(gen[8615]),
			.SE(gen[8616]),

			.SELF(gen[8520]),
			.cell_state(gen[8520])
		); 

/******************* CELL 8521 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8521 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8425]),
			.N(gen[8426]),
			.NE(gen[8427]),

			.O(gen[8520]),
			.E(gen[8522]),

			.SO(gen[8615]),
			.S(gen[8616]),
			.SE(gen[8617]),

			.SELF(gen[8521]),
			.cell_state(gen[8521])
		); 

/******************* CELL 8522 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8522 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8426]),
			.N(gen[8427]),
			.NE(gen[8428]),

			.O(gen[8521]),
			.E(gen[8523]),

			.SO(gen[8616]),
			.S(gen[8617]),
			.SE(gen[8618]),

			.SELF(gen[8522]),
			.cell_state(gen[8522])
		); 

/******************* CELL 8523 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8523 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8427]),
			.N(gen[8428]),
			.NE(gen[8429]),

			.O(gen[8522]),
			.E(gen[8524]),

			.SO(gen[8617]),
			.S(gen[8618]),
			.SE(gen[8619]),

			.SELF(gen[8523]),
			.cell_state(gen[8523])
		); 

/******************* CELL 8524 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8524 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8428]),
			.N(gen[8429]),
			.NE(gen[8430]),

			.O(gen[8523]),
			.E(gen[8525]),

			.SO(gen[8618]),
			.S(gen[8619]),
			.SE(gen[8620]),

			.SELF(gen[8524]),
			.cell_state(gen[8524])
		); 

/******************* CELL 8525 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8525 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8429]),
			.N(gen[8430]),
			.NE(gen[8431]),

			.O(gen[8524]),
			.E(gen[8526]),

			.SO(gen[8619]),
			.S(gen[8620]),
			.SE(gen[8621]),

			.SELF(gen[8525]),
			.cell_state(gen[8525])
		); 

/******************* CELL 8526 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8526 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8430]),
			.N(gen[8431]),
			.NE(gen[8432]),

			.O(gen[8525]),
			.E(gen[8527]),

			.SO(gen[8620]),
			.S(gen[8621]),
			.SE(gen[8622]),

			.SELF(gen[8526]),
			.cell_state(gen[8526])
		); 

/******************* CELL 8527 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8527 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8431]),
			.N(gen[8432]),
			.NE(gen[8433]),

			.O(gen[8526]),
			.E(gen[8528]),

			.SO(gen[8621]),
			.S(gen[8622]),
			.SE(gen[8623]),

			.SELF(gen[8527]),
			.cell_state(gen[8527])
		); 

/******************* CELL 8528 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8528 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8432]),
			.N(gen[8433]),
			.NE(gen[8434]),

			.O(gen[8527]),
			.E(gen[8529]),

			.SO(gen[8622]),
			.S(gen[8623]),
			.SE(gen[8624]),

			.SELF(gen[8528]),
			.cell_state(gen[8528])
		); 

/******************* CELL 8529 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8529 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8433]),
			.N(gen[8434]),
			.NE(gen[8435]),

			.O(gen[8528]),
			.E(gen[8530]),

			.SO(gen[8623]),
			.S(gen[8624]),
			.SE(gen[8625]),

			.SELF(gen[8529]),
			.cell_state(gen[8529])
		); 

/******************* CELL 8530 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8530 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8434]),
			.N(gen[8435]),
			.NE(gen[8436]),

			.O(gen[8529]),
			.E(gen[8531]),

			.SO(gen[8624]),
			.S(gen[8625]),
			.SE(gen[8626]),

			.SELF(gen[8530]),
			.cell_state(gen[8530])
		); 

/******************* CELL 8531 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8531 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8435]),
			.N(gen[8436]),
			.NE(gen[8437]),

			.O(gen[8530]),
			.E(gen[8532]),

			.SO(gen[8625]),
			.S(gen[8626]),
			.SE(gen[8627]),

			.SELF(gen[8531]),
			.cell_state(gen[8531])
		); 

/******************* CELL 8532 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8532 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8436]),
			.N(gen[8437]),
			.NE(gen[8438]),

			.O(gen[8531]),
			.E(gen[8533]),

			.SO(gen[8626]),
			.S(gen[8627]),
			.SE(gen[8628]),

			.SELF(gen[8532]),
			.cell_state(gen[8532])
		); 

/******************* CELL 8533 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8533 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8437]),
			.N(gen[8438]),
			.NE(gen[8439]),

			.O(gen[8532]),
			.E(gen[8534]),

			.SO(gen[8627]),
			.S(gen[8628]),
			.SE(gen[8629]),

			.SELF(gen[8533]),
			.cell_state(gen[8533])
		); 

/******************* CELL 8534 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8534 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8438]),
			.N(gen[8439]),
			.NE(gen[8440]),

			.O(gen[8533]),
			.E(gen[8535]),

			.SO(gen[8628]),
			.S(gen[8629]),
			.SE(gen[8630]),

			.SELF(gen[8534]),
			.cell_state(gen[8534])
		); 

/******************* CELL 8535 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8535 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8439]),
			.N(gen[8440]),
			.NE(gen[8441]),

			.O(gen[8534]),
			.E(gen[8536]),

			.SO(gen[8629]),
			.S(gen[8630]),
			.SE(gen[8631]),

			.SELF(gen[8535]),
			.cell_state(gen[8535])
		); 

/******************* CELL 8536 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8536 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8440]),
			.N(gen[8441]),
			.NE(gen[8442]),

			.O(gen[8535]),
			.E(gen[8537]),

			.SO(gen[8630]),
			.S(gen[8631]),
			.SE(gen[8632]),

			.SELF(gen[8536]),
			.cell_state(gen[8536])
		); 

/******************* CELL 8537 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8537 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8441]),
			.N(gen[8442]),
			.NE(gen[8443]),

			.O(gen[8536]),
			.E(gen[8538]),

			.SO(gen[8631]),
			.S(gen[8632]),
			.SE(gen[8633]),

			.SELF(gen[8537]),
			.cell_state(gen[8537])
		); 

/******************* CELL 8538 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8538 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8442]),
			.N(gen[8443]),
			.NE(gen[8444]),

			.O(gen[8537]),
			.E(gen[8539]),

			.SO(gen[8632]),
			.S(gen[8633]),
			.SE(gen[8634]),

			.SELF(gen[8538]),
			.cell_state(gen[8538])
		); 

/******************* CELL 8539 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8539 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8443]),
			.N(gen[8444]),
			.NE(gen[8445]),

			.O(gen[8538]),
			.E(gen[8540]),

			.SO(gen[8633]),
			.S(gen[8634]),
			.SE(gen[8635]),

			.SELF(gen[8539]),
			.cell_state(gen[8539])
		); 

/******************* CELL 8540 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8540 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8444]),
			.N(gen[8445]),
			.NE(gen[8446]),

			.O(gen[8539]),
			.E(gen[8541]),

			.SO(gen[8634]),
			.S(gen[8635]),
			.SE(gen[8636]),

			.SELF(gen[8540]),
			.cell_state(gen[8540])
		); 

/******************* CELL 8541 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8541 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8445]),
			.N(gen[8446]),
			.NE(gen[8447]),

			.O(gen[8540]),
			.E(gen[8542]),

			.SO(gen[8635]),
			.S(gen[8636]),
			.SE(gen[8637]),

			.SELF(gen[8541]),
			.cell_state(gen[8541])
		); 

/******************* CELL 8542 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8542 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8446]),
			.N(gen[8447]),
			.NE(gen[8448]),

			.O(gen[8541]),
			.E(gen[8543]),

			.SO(gen[8636]),
			.S(gen[8637]),
			.SE(gen[8638]),

			.SELF(gen[8542]),
			.cell_state(gen[8542])
		); 

/******************* CELL 8543 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8543 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8447]),
			.N(gen[8448]),
			.NE(gen[8449]),

			.O(gen[8542]),
			.E(gen[8544]),

			.SO(gen[8637]),
			.S(gen[8638]),
			.SE(gen[8639]),

			.SELF(gen[8543]),
			.cell_state(gen[8543])
		); 

/******************* CELL 8544 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8544 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8448]),
			.N(gen[8449]),
			.NE(gen[8450]),

			.O(gen[8543]),
			.E(gen[8545]),

			.SO(gen[8638]),
			.S(gen[8639]),
			.SE(gen[8640]),

			.SELF(gen[8544]),
			.cell_state(gen[8544])
		); 

/******************* CELL 8545 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8545 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8449]),
			.N(gen[8450]),
			.NE(gen[8451]),

			.O(gen[8544]),
			.E(gen[8546]),

			.SO(gen[8639]),
			.S(gen[8640]),
			.SE(gen[8641]),

			.SELF(gen[8545]),
			.cell_state(gen[8545])
		); 

/******************* CELL 8546 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8546 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8450]),
			.N(gen[8451]),
			.NE(gen[8452]),

			.O(gen[8545]),
			.E(gen[8547]),

			.SO(gen[8640]),
			.S(gen[8641]),
			.SE(gen[8642]),

			.SELF(gen[8546]),
			.cell_state(gen[8546])
		); 

/******************* CELL 8547 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8547 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8451]),
			.N(gen[8452]),
			.NE(gen[8453]),

			.O(gen[8546]),
			.E(gen[8548]),

			.SO(gen[8641]),
			.S(gen[8642]),
			.SE(gen[8643]),

			.SELF(gen[8547]),
			.cell_state(gen[8547])
		); 

/******************* CELL 8548 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8548 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8452]),
			.N(gen[8453]),
			.NE(gen[8454]),

			.O(gen[8547]),
			.E(gen[8549]),

			.SO(gen[8642]),
			.S(gen[8643]),
			.SE(gen[8644]),

			.SELF(gen[8548]),
			.cell_state(gen[8548])
		); 

/******************* CELL 8549 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8549 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8453]),
			.N(gen[8454]),
			.NE(gen[8453]),

			.O(gen[8548]),
			.E(gen[8548]),

			.SO(gen[8643]),
			.S(gen[8644]),
			.SE(gen[8643]),

			.SELF(gen[8549]),
			.cell_state(gen[8549])
		); 

/******************* CELL 8550 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8550 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8456]),
			.N(gen[8455]),
			.NE(gen[8456]),

			.O(gen[8551]),
			.E(gen[8551]),

			.SO(gen[8646]),
			.S(gen[8645]),
			.SE(gen[8646]),

			.SELF(gen[8550]),
			.cell_state(gen[8550])
		); 

/******************* CELL 8551 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8551 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8455]),
			.N(gen[8456]),
			.NE(gen[8457]),

			.O(gen[8550]),
			.E(gen[8552]),

			.SO(gen[8645]),
			.S(gen[8646]),
			.SE(gen[8647]),

			.SELF(gen[8551]),
			.cell_state(gen[8551])
		); 

/******************* CELL 8552 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8552 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8456]),
			.N(gen[8457]),
			.NE(gen[8458]),

			.O(gen[8551]),
			.E(gen[8553]),

			.SO(gen[8646]),
			.S(gen[8647]),
			.SE(gen[8648]),

			.SELF(gen[8552]),
			.cell_state(gen[8552])
		); 

/******************* CELL 8553 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8553 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8457]),
			.N(gen[8458]),
			.NE(gen[8459]),

			.O(gen[8552]),
			.E(gen[8554]),

			.SO(gen[8647]),
			.S(gen[8648]),
			.SE(gen[8649]),

			.SELF(gen[8553]),
			.cell_state(gen[8553])
		); 

/******************* CELL 8554 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8554 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8458]),
			.N(gen[8459]),
			.NE(gen[8460]),

			.O(gen[8553]),
			.E(gen[8555]),

			.SO(gen[8648]),
			.S(gen[8649]),
			.SE(gen[8650]),

			.SELF(gen[8554]),
			.cell_state(gen[8554])
		); 

/******************* CELL 8555 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8555 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8459]),
			.N(gen[8460]),
			.NE(gen[8461]),

			.O(gen[8554]),
			.E(gen[8556]),

			.SO(gen[8649]),
			.S(gen[8650]),
			.SE(gen[8651]),

			.SELF(gen[8555]),
			.cell_state(gen[8555])
		); 

/******************* CELL 8556 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8556 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8460]),
			.N(gen[8461]),
			.NE(gen[8462]),

			.O(gen[8555]),
			.E(gen[8557]),

			.SO(gen[8650]),
			.S(gen[8651]),
			.SE(gen[8652]),

			.SELF(gen[8556]),
			.cell_state(gen[8556])
		); 

/******************* CELL 8557 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8557 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8461]),
			.N(gen[8462]),
			.NE(gen[8463]),

			.O(gen[8556]),
			.E(gen[8558]),

			.SO(gen[8651]),
			.S(gen[8652]),
			.SE(gen[8653]),

			.SELF(gen[8557]),
			.cell_state(gen[8557])
		); 

/******************* CELL 8558 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8558 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8462]),
			.N(gen[8463]),
			.NE(gen[8464]),

			.O(gen[8557]),
			.E(gen[8559]),

			.SO(gen[8652]),
			.S(gen[8653]),
			.SE(gen[8654]),

			.SELF(gen[8558]),
			.cell_state(gen[8558])
		); 

/******************* CELL 8559 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8559 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8463]),
			.N(gen[8464]),
			.NE(gen[8465]),

			.O(gen[8558]),
			.E(gen[8560]),

			.SO(gen[8653]),
			.S(gen[8654]),
			.SE(gen[8655]),

			.SELF(gen[8559]),
			.cell_state(gen[8559])
		); 

/******************* CELL 8560 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8560 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8464]),
			.N(gen[8465]),
			.NE(gen[8466]),

			.O(gen[8559]),
			.E(gen[8561]),

			.SO(gen[8654]),
			.S(gen[8655]),
			.SE(gen[8656]),

			.SELF(gen[8560]),
			.cell_state(gen[8560])
		); 

/******************* CELL 8561 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8561 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8465]),
			.N(gen[8466]),
			.NE(gen[8467]),

			.O(gen[8560]),
			.E(gen[8562]),

			.SO(gen[8655]),
			.S(gen[8656]),
			.SE(gen[8657]),

			.SELF(gen[8561]),
			.cell_state(gen[8561])
		); 

/******************* CELL 8562 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8562 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8466]),
			.N(gen[8467]),
			.NE(gen[8468]),

			.O(gen[8561]),
			.E(gen[8563]),

			.SO(gen[8656]),
			.S(gen[8657]),
			.SE(gen[8658]),

			.SELF(gen[8562]),
			.cell_state(gen[8562])
		); 

/******************* CELL 8563 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8563 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8467]),
			.N(gen[8468]),
			.NE(gen[8469]),

			.O(gen[8562]),
			.E(gen[8564]),

			.SO(gen[8657]),
			.S(gen[8658]),
			.SE(gen[8659]),

			.SELF(gen[8563]),
			.cell_state(gen[8563])
		); 

/******************* CELL 8564 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8564 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8468]),
			.N(gen[8469]),
			.NE(gen[8470]),

			.O(gen[8563]),
			.E(gen[8565]),

			.SO(gen[8658]),
			.S(gen[8659]),
			.SE(gen[8660]),

			.SELF(gen[8564]),
			.cell_state(gen[8564])
		); 

/******************* CELL 8565 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8565 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8469]),
			.N(gen[8470]),
			.NE(gen[8471]),

			.O(gen[8564]),
			.E(gen[8566]),

			.SO(gen[8659]),
			.S(gen[8660]),
			.SE(gen[8661]),

			.SELF(gen[8565]),
			.cell_state(gen[8565])
		); 

/******************* CELL 8566 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8566 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8470]),
			.N(gen[8471]),
			.NE(gen[8472]),

			.O(gen[8565]),
			.E(gen[8567]),

			.SO(gen[8660]),
			.S(gen[8661]),
			.SE(gen[8662]),

			.SELF(gen[8566]),
			.cell_state(gen[8566])
		); 

/******************* CELL 8567 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8567 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8471]),
			.N(gen[8472]),
			.NE(gen[8473]),

			.O(gen[8566]),
			.E(gen[8568]),

			.SO(gen[8661]),
			.S(gen[8662]),
			.SE(gen[8663]),

			.SELF(gen[8567]),
			.cell_state(gen[8567])
		); 

/******************* CELL 8568 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8568 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8472]),
			.N(gen[8473]),
			.NE(gen[8474]),

			.O(gen[8567]),
			.E(gen[8569]),

			.SO(gen[8662]),
			.S(gen[8663]),
			.SE(gen[8664]),

			.SELF(gen[8568]),
			.cell_state(gen[8568])
		); 

/******************* CELL 8569 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8569 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8473]),
			.N(gen[8474]),
			.NE(gen[8475]),

			.O(gen[8568]),
			.E(gen[8570]),

			.SO(gen[8663]),
			.S(gen[8664]),
			.SE(gen[8665]),

			.SELF(gen[8569]),
			.cell_state(gen[8569])
		); 

/******************* CELL 8570 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8570 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8474]),
			.N(gen[8475]),
			.NE(gen[8476]),

			.O(gen[8569]),
			.E(gen[8571]),

			.SO(gen[8664]),
			.S(gen[8665]),
			.SE(gen[8666]),

			.SELF(gen[8570]),
			.cell_state(gen[8570])
		); 

/******************* CELL 8571 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8571 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8475]),
			.N(gen[8476]),
			.NE(gen[8477]),

			.O(gen[8570]),
			.E(gen[8572]),

			.SO(gen[8665]),
			.S(gen[8666]),
			.SE(gen[8667]),

			.SELF(gen[8571]),
			.cell_state(gen[8571])
		); 

/******************* CELL 8572 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8572 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8476]),
			.N(gen[8477]),
			.NE(gen[8478]),

			.O(gen[8571]),
			.E(gen[8573]),

			.SO(gen[8666]),
			.S(gen[8667]),
			.SE(gen[8668]),

			.SELF(gen[8572]),
			.cell_state(gen[8572])
		); 

/******************* CELL 8573 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8573 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8477]),
			.N(gen[8478]),
			.NE(gen[8479]),

			.O(gen[8572]),
			.E(gen[8574]),

			.SO(gen[8667]),
			.S(gen[8668]),
			.SE(gen[8669]),

			.SELF(gen[8573]),
			.cell_state(gen[8573])
		); 

/******************* CELL 8574 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8574 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8478]),
			.N(gen[8479]),
			.NE(gen[8480]),

			.O(gen[8573]),
			.E(gen[8575]),

			.SO(gen[8668]),
			.S(gen[8669]),
			.SE(gen[8670]),

			.SELF(gen[8574]),
			.cell_state(gen[8574])
		); 

/******************* CELL 8575 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8575 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8479]),
			.N(gen[8480]),
			.NE(gen[8481]),

			.O(gen[8574]),
			.E(gen[8576]),

			.SO(gen[8669]),
			.S(gen[8670]),
			.SE(gen[8671]),

			.SELF(gen[8575]),
			.cell_state(gen[8575])
		); 

/******************* CELL 8576 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8576 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8480]),
			.N(gen[8481]),
			.NE(gen[8482]),

			.O(gen[8575]),
			.E(gen[8577]),

			.SO(gen[8670]),
			.S(gen[8671]),
			.SE(gen[8672]),

			.SELF(gen[8576]),
			.cell_state(gen[8576])
		); 

/******************* CELL 8577 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8577 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8481]),
			.N(gen[8482]),
			.NE(gen[8483]),

			.O(gen[8576]),
			.E(gen[8578]),

			.SO(gen[8671]),
			.S(gen[8672]),
			.SE(gen[8673]),

			.SELF(gen[8577]),
			.cell_state(gen[8577])
		); 

/******************* CELL 8578 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8578 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8482]),
			.N(gen[8483]),
			.NE(gen[8484]),

			.O(gen[8577]),
			.E(gen[8579]),

			.SO(gen[8672]),
			.S(gen[8673]),
			.SE(gen[8674]),

			.SELF(gen[8578]),
			.cell_state(gen[8578])
		); 

/******************* CELL 8579 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8579 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8483]),
			.N(gen[8484]),
			.NE(gen[8485]),

			.O(gen[8578]),
			.E(gen[8580]),

			.SO(gen[8673]),
			.S(gen[8674]),
			.SE(gen[8675]),

			.SELF(gen[8579]),
			.cell_state(gen[8579])
		); 

/******************* CELL 8580 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8580 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8484]),
			.N(gen[8485]),
			.NE(gen[8486]),

			.O(gen[8579]),
			.E(gen[8581]),

			.SO(gen[8674]),
			.S(gen[8675]),
			.SE(gen[8676]),

			.SELF(gen[8580]),
			.cell_state(gen[8580])
		); 

/******************* CELL 8581 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8581 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8485]),
			.N(gen[8486]),
			.NE(gen[8487]),

			.O(gen[8580]),
			.E(gen[8582]),

			.SO(gen[8675]),
			.S(gen[8676]),
			.SE(gen[8677]),

			.SELF(gen[8581]),
			.cell_state(gen[8581])
		); 

/******************* CELL 8582 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8582 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8486]),
			.N(gen[8487]),
			.NE(gen[8488]),

			.O(gen[8581]),
			.E(gen[8583]),

			.SO(gen[8676]),
			.S(gen[8677]),
			.SE(gen[8678]),

			.SELF(gen[8582]),
			.cell_state(gen[8582])
		); 

/******************* CELL 8583 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8583 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8487]),
			.N(gen[8488]),
			.NE(gen[8489]),

			.O(gen[8582]),
			.E(gen[8584]),

			.SO(gen[8677]),
			.S(gen[8678]),
			.SE(gen[8679]),

			.SELF(gen[8583]),
			.cell_state(gen[8583])
		); 

/******************* CELL 8584 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8584 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8488]),
			.N(gen[8489]),
			.NE(gen[8490]),

			.O(gen[8583]),
			.E(gen[8585]),

			.SO(gen[8678]),
			.S(gen[8679]),
			.SE(gen[8680]),

			.SELF(gen[8584]),
			.cell_state(gen[8584])
		); 

/******************* CELL 8585 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8585 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8489]),
			.N(gen[8490]),
			.NE(gen[8491]),

			.O(gen[8584]),
			.E(gen[8586]),

			.SO(gen[8679]),
			.S(gen[8680]),
			.SE(gen[8681]),

			.SELF(gen[8585]),
			.cell_state(gen[8585])
		); 

/******************* CELL 8586 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8586 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8490]),
			.N(gen[8491]),
			.NE(gen[8492]),

			.O(gen[8585]),
			.E(gen[8587]),

			.SO(gen[8680]),
			.S(gen[8681]),
			.SE(gen[8682]),

			.SELF(gen[8586]),
			.cell_state(gen[8586])
		); 

/******************* CELL 8587 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8587 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8491]),
			.N(gen[8492]),
			.NE(gen[8493]),

			.O(gen[8586]),
			.E(gen[8588]),

			.SO(gen[8681]),
			.S(gen[8682]),
			.SE(gen[8683]),

			.SELF(gen[8587]),
			.cell_state(gen[8587])
		); 

/******************* CELL 8588 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8588 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8492]),
			.N(gen[8493]),
			.NE(gen[8494]),

			.O(gen[8587]),
			.E(gen[8589]),

			.SO(gen[8682]),
			.S(gen[8683]),
			.SE(gen[8684]),

			.SELF(gen[8588]),
			.cell_state(gen[8588])
		); 

/******************* CELL 8589 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8589 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8493]),
			.N(gen[8494]),
			.NE(gen[8495]),

			.O(gen[8588]),
			.E(gen[8590]),

			.SO(gen[8683]),
			.S(gen[8684]),
			.SE(gen[8685]),

			.SELF(gen[8589]),
			.cell_state(gen[8589])
		); 

/******************* CELL 8590 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8590 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8494]),
			.N(gen[8495]),
			.NE(gen[8496]),

			.O(gen[8589]),
			.E(gen[8591]),

			.SO(gen[8684]),
			.S(gen[8685]),
			.SE(gen[8686]),

			.SELF(gen[8590]),
			.cell_state(gen[8590])
		); 

/******************* CELL 8591 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8591 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8495]),
			.N(gen[8496]),
			.NE(gen[8497]),

			.O(gen[8590]),
			.E(gen[8592]),

			.SO(gen[8685]),
			.S(gen[8686]),
			.SE(gen[8687]),

			.SELF(gen[8591]),
			.cell_state(gen[8591])
		); 

/******************* CELL 8592 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8592 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8496]),
			.N(gen[8497]),
			.NE(gen[8498]),

			.O(gen[8591]),
			.E(gen[8593]),

			.SO(gen[8686]),
			.S(gen[8687]),
			.SE(gen[8688]),

			.SELF(gen[8592]),
			.cell_state(gen[8592])
		); 

/******************* CELL 8593 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8593 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8497]),
			.N(gen[8498]),
			.NE(gen[8499]),

			.O(gen[8592]),
			.E(gen[8594]),

			.SO(gen[8687]),
			.S(gen[8688]),
			.SE(gen[8689]),

			.SELF(gen[8593]),
			.cell_state(gen[8593])
		); 

/******************* CELL 8594 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8594 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8498]),
			.N(gen[8499]),
			.NE(gen[8500]),

			.O(gen[8593]),
			.E(gen[8595]),

			.SO(gen[8688]),
			.S(gen[8689]),
			.SE(gen[8690]),

			.SELF(gen[8594]),
			.cell_state(gen[8594])
		); 

/******************* CELL 8595 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8595 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8499]),
			.N(gen[8500]),
			.NE(gen[8501]),

			.O(gen[8594]),
			.E(gen[8596]),

			.SO(gen[8689]),
			.S(gen[8690]),
			.SE(gen[8691]),

			.SELF(gen[8595]),
			.cell_state(gen[8595])
		); 

/******************* CELL 8596 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8596 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8500]),
			.N(gen[8501]),
			.NE(gen[8502]),

			.O(gen[8595]),
			.E(gen[8597]),

			.SO(gen[8690]),
			.S(gen[8691]),
			.SE(gen[8692]),

			.SELF(gen[8596]),
			.cell_state(gen[8596])
		); 

/******************* CELL 8597 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8597 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8501]),
			.N(gen[8502]),
			.NE(gen[8503]),

			.O(gen[8596]),
			.E(gen[8598]),

			.SO(gen[8691]),
			.S(gen[8692]),
			.SE(gen[8693]),

			.SELF(gen[8597]),
			.cell_state(gen[8597])
		); 

/******************* CELL 8598 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8598 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8502]),
			.N(gen[8503]),
			.NE(gen[8504]),

			.O(gen[8597]),
			.E(gen[8599]),

			.SO(gen[8692]),
			.S(gen[8693]),
			.SE(gen[8694]),

			.SELF(gen[8598]),
			.cell_state(gen[8598])
		); 

/******************* CELL 8599 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8599 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8503]),
			.N(gen[8504]),
			.NE(gen[8505]),

			.O(gen[8598]),
			.E(gen[8600]),

			.SO(gen[8693]),
			.S(gen[8694]),
			.SE(gen[8695]),

			.SELF(gen[8599]),
			.cell_state(gen[8599])
		); 

/******************* CELL 8600 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8600 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8504]),
			.N(gen[8505]),
			.NE(gen[8506]),

			.O(gen[8599]),
			.E(gen[8601]),

			.SO(gen[8694]),
			.S(gen[8695]),
			.SE(gen[8696]),

			.SELF(gen[8600]),
			.cell_state(gen[8600])
		); 

/******************* CELL 8601 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8601 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8505]),
			.N(gen[8506]),
			.NE(gen[8507]),

			.O(gen[8600]),
			.E(gen[8602]),

			.SO(gen[8695]),
			.S(gen[8696]),
			.SE(gen[8697]),

			.SELF(gen[8601]),
			.cell_state(gen[8601])
		); 

/******************* CELL 8602 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8602 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8506]),
			.N(gen[8507]),
			.NE(gen[8508]),

			.O(gen[8601]),
			.E(gen[8603]),

			.SO(gen[8696]),
			.S(gen[8697]),
			.SE(gen[8698]),

			.SELF(gen[8602]),
			.cell_state(gen[8602])
		); 

/******************* CELL 8603 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8603 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8507]),
			.N(gen[8508]),
			.NE(gen[8509]),

			.O(gen[8602]),
			.E(gen[8604]),

			.SO(gen[8697]),
			.S(gen[8698]),
			.SE(gen[8699]),

			.SELF(gen[8603]),
			.cell_state(gen[8603])
		); 

/******************* CELL 8604 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8604 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8508]),
			.N(gen[8509]),
			.NE(gen[8510]),

			.O(gen[8603]),
			.E(gen[8605]),

			.SO(gen[8698]),
			.S(gen[8699]),
			.SE(gen[8700]),

			.SELF(gen[8604]),
			.cell_state(gen[8604])
		); 

/******************* CELL 8605 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8605 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8509]),
			.N(gen[8510]),
			.NE(gen[8511]),

			.O(gen[8604]),
			.E(gen[8606]),

			.SO(gen[8699]),
			.S(gen[8700]),
			.SE(gen[8701]),

			.SELF(gen[8605]),
			.cell_state(gen[8605])
		); 

/******************* CELL 8606 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8606 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8510]),
			.N(gen[8511]),
			.NE(gen[8512]),

			.O(gen[8605]),
			.E(gen[8607]),

			.SO(gen[8700]),
			.S(gen[8701]),
			.SE(gen[8702]),

			.SELF(gen[8606]),
			.cell_state(gen[8606])
		); 

/******************* CELL 8607 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8607 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8511]),
			.N(gen[8512]),
			.NE(gen[8513]),

			.O(gen[8606]),
			.E(gen[8608]),

			.SO(gen[8701]),
			.S(gen[8702]),
			.SE(gen[8703]),

			.SELF(gen[8607]),
			.cell_state(gen[8607])
		); 

/******************* CELL 8608 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8608 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8512]),
			.N(gen[8513]),
			.NE(gen[8514]),

			.O(gen[8607]),
			.E(gen[8609]),

			.SO(gen[8702]),
			.S(gen[8703]),
			.SE(gen[8704]),

			.SELF(gen[8608]),
			.cell_state(gen[8608])
		); 

/******************* CELL 8609 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8609 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8513]),
			.N(gen[8514]),
			.NE(gen[8515]),

			.O(gen[8608]),
			.E(gen[8610]),

			.SO(gen[8703]),
			.S(gen[8704]),
			.SE(gen[8705]),

			.SELF(gen[8609]),
			.cell_state(gen[8609])
		); 

/******************* CELL 8610 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8610 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8514]),
			.N(gen[8515]),
			.NE(gen[8516]),

			.O(gen[8609]),
			.E(gen[8611]),

			.SO(gen[8704]),
			.S(gen[8705]),
			.SE(gen[8706]),

			.SELF(gen[8610]),
			.cell_state(gen[8610])
		); 

/******************* CELL 8611 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8611 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8515]),
			.N(gen[8516]),
			.NE(gen[8517]),

			.O(gen[8610]),
			.E(gen[8612]),

			.SO(gen[8705]),
			.S(gen[8706]),
			.SE(gen[8707]),

			.SELF(gen[8611]),
			.cell_state(gen[8611])
		); 

/******************* CELL 8612 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8612 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8516]),
			.N(gen[8517]),
			.NE(gen[8518]),

			.O(gen[8611]),
			.E(gen[8613]),

			.SO(gen[8706]),
			.S(gen[8707]),
			.SE(gen[8708]),

			.SELF(gen[8612]),
			.cell_state(gen[8612])
		); 

/******************* CELL 8613 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8613 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8517]),
			.N(gen[8518]),
			.NE(gen[8519]),

			.O(gen[8612]),
			.E(gen[8614]),

			.SO(gen[8707]),
			.S(gen[8708]),
			.SE(gen[8709]),

			.SELF(gen[8613]),
			.cell_state(gen[8613])
		); 

/******************* CELL 8614 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8614 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8518]),
			.N(gen[8519]),
			.NE(gen[8520]),

			.O(gen[8613]),
			.E(gen[8615]),

			.SO(gen[8708]),
			.S(gen[8709]),
			.SE(gen[8710]),

			.SELF(gen[8614]),
			.cell_state(gen[8614])
		); 

/******************* CELL 8615 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8615 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8519]),
			.N(gen[8520]),
			.NE(gen[8521]),

			.O(gen[8614]),
			.E(gen[8616]),

			.SO(gen[8709]),
			.S(gen[8710]),
			.SE(gen[8711]),

			.SELF(gen[8615]),
			.cell_state(gen[8615])
		); 

/******************* CELL 8616 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8616 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8520]),
			.N(gen[8521]),
			.NE(gen[8522]),

			.O(gen[8615]),
			.E(gen[8617]),

			.SO(gen[8710]),
			.S(gen[8711]),
			.SE(gen[8712]),

			.SELF(gen[8616]),
			.cell_state(gen[8616])
		); 

/******************* CELL 8617 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8617 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8521]),
			.N(gen[8522]),
			.NE(gen[8523]),

			.O(gen[8616]),
			.E(gen[8618]),

			.SO(gen[8711]),
			.S(gen[8712]),
			.SE(gen[8713]),

			.SELF(gen[8617]),
			.cell_state(gen[8617])
		); 

/******************* CELL 8618 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8618 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8522]),
			.N(gen[8523]),
			.NE(gen[8524]),

			.O(gen[8617]),
			.E(gen[8619]),

			.SO(gen[8712]),
			.S(gen[8713]),
			.SE(gen[8714]),

			.SELF(gen[8618]),
			.cell_state(gen[8618])
		); 

/******************* CELL 8619 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8619 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8523]),
			.N(gen[8524]),
			.NE(gen[8525]),

			.O(gen[8618]),
			.E(gen[8620]),

			.SO(gen[8713]),
			.S(gen[8714]),
			.SE(gen[8715]),

			.SELF(gen[8619]),
			.cell_state(gen[8619])
		); 

/******************* CELL 8620 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8620 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8524]),
			.N(gen[8525]),
			.NE(gen[8526]),

			.O(gen[8619]),
			.E(gen[8621]),

			.SO(gen[8714]),
			.S(gen[8715]),
			.SE(gen[8716]),

			.SELF(gen[8620]),
			.cell_state(gen[8620])
		); 

/******************* CELL 8621 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8621 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8525]),
			.N(gen[8526]),
			.NE(gen[8527]),

			.O(gen[8620]),
			.E(gen[8622]),

			.SO(gen[8715]),
			.S(gen[8716]),
			.SE(gen[8717]),

			.SELF(gen[8621]),
			.cell_state(gen[8621])
		); 

/******************* CELL 8622 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8622 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8526]),
			.N(gen[8527]),
			.NE(gen[8528]),

			.O(gen[8621]),
			.E(gen[8623]),

			.SO(gen[8716]),
			.S(gen[8717]),
			.SE(gen[8718]),

			.SELF(gen[8622]),
			.cell_state(gen[8622])
		); 

/******************* CELL 8623 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8623 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8527]),
			.N(gen[8528]),
			.NE(gen[8529]),

			.O(gen[8622]),
			.E(gen[8624]),

			.SO(gen[8717]),
			.S(gen[8718]),
			.SE(gen[8719]),

			.SELF(gen[8623]),
			.cell_state(gen[8623])
		); 

/******************* CELL 8624 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8624 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8528]),
			.N(gen[8529]),
			.NE(gen[8530]),

			.O(gen[8623]),
			.E(gen[8625]),

			.SO(gen[8718]),
			.S(gen[8719]),
			.SE(gen[8720]),

			.SELF(gen[8624]),
			.cell_state(gen[8624])
		); 

/******************* CELL 8625 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8625 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8529]),
			.N(gen[8530]),
			.NE(gen[8531]),

			.O(gen[8624]),
			.E(gen[8626]),

			.SO(gen[8719]),
			.S(gen[8720]),
			.SE(gen[8721]),

			.SELF(gen[8625]),
			.cell_state(gen[8625])
		); 

/******************* CELL 8626 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8626 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8530]),
			.N(gen[8531]),
			.NE(gen[8532]),

			.O(gen[8625]),
			.E(gen[8627]),

			.SO(gen[8720]),
			.S(gen[8721]),
			.SE(gen[8722]),

			.SELF(gen[8626]),
			.cell_state(gen[8626])
		); 

/******************* CELL 8627 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8627 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8531]),
			.N(gen[8532]),
			.NE(gen[8533]),

			.O(gen[8626]),
			.E(gen[8628]),

			.SO(gen[8721]),
			.S(gen[8722]),
			.SE(gen[8723]),

			.SELF(gen[8627]),
			.cell_state(gen[8627])
		); 

/******************* CELL 8628 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8628 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8532]),
			.N(gen[8533]),
			.NE(gen[8534]),

			.O(gen[8627]),
			.E(gen[8629]),

			.SO(gen[8722]),
			.S(gen[8723]),
			.SE(gen[8724]),

			.SELF(gen[8628]),
			.cell_state(gen[8628])
		); 

/******************* CELL 8629 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8629 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8533]),
			.N(gen[8534]),
			.NE(gen[8535]),

			.O(gen[8628]),
			.E(gen[8630]),

			.SO(gen[8723]),
			.S(gen[8724]),
			.SE(gen[8725]),

			.SELF(gen[8629]),
			.cell_state(gen[8629])
		); 

/******************* CELL 8630 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8630 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8534]),
			.N(gen[8535]),
			.NE(gen[8536]),

			.O(gen[8629]),
			.E(gen[8631]),

			.SO(gen[8724]),
			.S(gen[8725]),
			.SE(gen[8726]),

			.SELF(gen[8630]),
			.cell_state(gen[8630])
		); 

/******************* CELL 8631 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8631 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8535]),
			.N(gen[8536]),
			.NE(gen[8537]),

			.O(gen[8630]),
			.E(gen[8632]),

			.SO(gen[8725]),
			.S(gen[8726]),
			.SE(gen[8727]),

			.SELF(gen[8631]),
			.cell_state(gen[8631])
		); 

/******************* CELL 8632 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8632 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8536]),
			.N(gen[8537]),
			.NE(gen[8538]),

			.O(gen[8631]),
			.E(gen[8633]),

			.SO(gen[8726]),
			.S(gen[8727]),
			.SE(gen[8728]),

			.SELF(gen[8632]),
			.cell_state(gen[8632])
		); 

/******************* CELL 8633 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8633 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8537]),
			.N(gen[8538]),
			.NE(gen[8539]),

			.O(gen[8632]),
			.E(gen[8634]),

			.SO(gen[8727]),
			.S(gen[8728]),
			.SE(gen[8729]),

			.SELF(gen[8633]),
			.cell_state(gen[8633])
		); 

/******************* CELL 8634 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8634 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8538]),
			.N(gen[8539]),
			.NE(gen[8540]),

			.O(gen[8633]),
			.E(gen[8635]),

			.SO(gen[8728]),
			.S(gen[8729]),
			.SE(gen[8730]),

			.SELF(gen[8634]),
			.cell_state(gen[8634])
		); 

/******************* CELL 8635 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8635 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8539]),
			.N(gen[8540]),
			.NE(gen[8541]),

			.O(gen[8634]),
			.E(gen[8636]),

			.SO(gen[8729]),
			.S(gen[8730]),
			.SE(gen[8731]),

			.SELF(gen[8635]),
			.cell_state(gen[8635])
		); 

/******************* CELL 8636 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8636 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8540]),
			.N(gen[8541]),
			.NE(gen[8542]),

			.O(gen[8635]),
			.E(gen[8637]),

			.SO(gen[8730]),
			.S(gen[8731]),
			.SE(gen[8732]),

			.SELF(gen[8636]),
			.cell_state(gen[8636])
		); 

/******************* CELL 8637 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8637 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8541]),
			.N(gen[8542]),
			.NE(gen[8543]),

			.O(gen[8636]),
			.E(gen[8638]),

			.SO(gen[8731]),
			.S(gen[8732]),
			.SE(gen[8733]),

			.SELF(gen[8637]),
			.cell_state(gen[8637])
		); 

/******************* CELL 8638 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8638 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8542]),
			.N(gen[8543]),
			.NE(gen[8544]),

			.O(gen[8637]),
			.E(gen[8639]),

			.SO(gen[8732]),
			.S(gen[8733]),
			.SE(gen[8734]),

			.SELF(gen[8638]),
			.cell_state(gen[8638])
		); 

/******************* CELL 8639 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8639 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8543]),
			.N(gen[8544]),
			.NE(gen[8545]),

			.O(gen[8638]),
			.E(gen[8640]),

			.SO(gen[8733]),
			.S(gen[8734]),
			.SE(gen[8735]),

			.SELF(gen[8639]),
			.cell_state(gen[8639])
		); 

/******************* CELL 8640 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8640 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8544]),
			.N(gen[8545]),
			.NE(gen[8546]),

			.O(gen[8639]),
			.E(gen[8641]),

			.SO(gen[8734]),
			.S(gen[8735]),
			.SE(gen[8736]),

			.SELF(gen[8640]),
			.cell_state(gen[8640])
		); 

/******************* CELL 8641 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8641 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8545]),
			.N(gen[8546]),
			.NE(gen[8547]),

			.O(gen[8640]),
			.E(gen[8642]),

			.SO(gen[8735]),
			.S(gen[8736]),
			.SE(gen[8737]),

			.SELF(gen[8641]),
			.cell_state(gen[8641])
		); 

/******************* CELL 8642 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8642 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8546]),
			.N(gen[8547]),
			.NE(gen[8548]),

			.O(gen[8641]),
			.E(gen[8643]),

			.SO(gen[8736]),
			.S(gen[8737]),
			.SE(gen[8738]),

			.SELF(gen[8642]),
			.cell_state(gen[8642])
		); 

/******************* CELL 8643 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8643 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8547]),
			.N(gen[8548]),
			.NE(gen[8549]),

			.O(gen[8642]),
			.E(gen[8644]),

			.SO(gen[8737]),
			.S(gen[8738]),
			.SE(gen[8739]),

			.SELF(gen[8643]),
			.cell_state(gen[8643])
		); 

/******************* CELL 8644 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8644 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8548]),
			.N(gen[8549]),
			.NE(gen[8548]),

			.O(gen[8643]),
			.E(gen[8643]),

			.SO(gen[8738]),
			.S(gen[8739]),
			.SE(gen[8738]),

			.SELF(gen[8644]),
			.cell_state(gen[8644])
		); 

/******************* CELL 8645 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8645 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8551]),
			.N(gen[8550]),
			.NE(gen[8551]),

			.O(gen[8646]),
			.E(gen[8646]),

			.SO(gen[8741]),
			.S(gen[8740]),
			.SE(gen[8741]),

			.SELF(gen[8645]),
			.cell_state(gen[8645])
		); 

/******************* CELL 8646 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8646 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8550]),
			.N(gen[8551]),
			.NE(gen[8552]),

			.O(gen[8645]),
			.E(gen[8647]),

			.SO(gen[8740]),
			.S(gen[8741]),
			.SE(gen[8742]),

			.SELF(gen[8646]),
			.cell_state(gen[8646])
		); 

/******************* CELL 8647 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8647 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8551]),
			.N(gen[8552]),
			.NE(gen[8553]),

			.O(gen[8646]),
			.E(gen[8648]),

			.SO(gen[8741]),
			.S(gen[8742]),
			.SE(gen[8743]),

			.SELF(gen[8647]),
			.cell_state(gen[8647])
		); 

/******************* CELL 8648 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8648 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8552]),
			.N(gen[8553]),
			.NE(gen[8554]),

			.O(gen[8647]),
			.E(gen[8649]),

			.SO(gen[8742]),
			.S(gen[8743]),
			.SE(gen[8744]),

			.SELF(gen[8648]),
			.cell_state(gen[8648])
		); 

/******************* CELL 8649 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8649 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8553]),
			.N(gen[8554]),
			.NE(gen[8555]),

			.O(gen[8648]),
			.E(gen[8650]),

			.SO(gen[8743]),
			.S(gen[8744]),
			.SE(gen[8745]),

			.SELF(gen[8649]),
			.cell_state(gen[8649])
		); 

/******************* CELL 8650 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8650 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8554]),
			.N(gen[8555]),
			.NE(gen[8556]),

			.O(gen[8649]),
			.E(gen[8651]),

			.SO(gen[8744]),
			.S(gen[8745]),
			.SE(gen[8746]),

			.SELF(gen[8650]),
			.cell_state(gen[8650])
		); 

/******************* CELL 8651 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8651 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8555]),
			.N(gen[8556]),
			.NE(gen[8557]),

			.O(gen[8650]),
			.E(gen[8652]),

			.SO(gen[8745]),
			.S(gen[8746]),
			.SE(gen[8747]),

			.SELF(gen[8651]),
			.cell_state(gen[8651])
		); 

/******************* CELL 8652 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8652 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8556]),
			.N(gen[8557]),
			.NE(gen[8558]),

			.O(gen[8651]),
			.E(gen[8653]),

			.SO(gen[8746]),
			.S(gen[8747]),
			.SE(gen[8748]),

			.SELF(gen[8652]),
			.cell_state(gen[8652])
		); 

/******************* CELL 8653 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8653 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8557]),
			.N(gen[8558]),
			.NE(gen[8559]),

			.O(gen[8652]),
			.E(gen[8654]),

			.SO(gen[8747]),
			.S(gen[8748]),
			.SE(gen[8749]),

			.SELF(gen[8653]),
			.cell_state(gen[8653])
		); 

/******************* CELL 8654 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8654 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8558]),
			.N(gen[8559]),
			.NE(gen[8560]),

			.O(gen[8653]),
			.E(gen[8655]),

			.SO(gen[8748]),
			.S(gen[8749]),
			.SE(gen[8750]),

			.SELF(gen[8654]),
			.cell_state(gen[8654])
		); 

/******************* CELL 8655 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8655 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8559]),
			.N(gen[8560]),
			.NE(gen[8561]),

			.O(gen[8654]),
			.E(gen[8656]),

			.SO(gen[8749]),
			.S(gen[8750]),
			.SE(gen[8751]),

			.SELF(gen[8655]),
			.cell_state(gen[8655])
		); 

/******************* CELL 8656 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8656 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8560]),
			.N(gen[8561]),
			.NE(gen[8562]),

			.O(gen[8655]),
			.E(gen[8657]),

			.SO(gen[8750]),
			.S(gen[8751]),
			.SE(gen[8752]),

			.SELF(gen[8656]),
			.cell_state(gen[8656])
		); 

/******************* CELL 8657 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8657 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8561]),
			.N(gen[8562]),
			.NE(gen[8563]),

			.O(gen[8656]),
			.E(gen[8658]),

			.SO(gen[8751]),
			.S(gen[8752]),
			.SE(gen[8753]),

			.SELF(gen[8657]),
			.cell_state(gen[8657])
		); 

/******************* CELL 8658 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8658 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8562]),
			.N(gen[8563]),
			.NE(gen[8564]),

			.O(gen[8657]),
			.E(gen[8659]),

			.SO(gen[8752]),
			.S(gen[8753]),
			.SE(gen[8754]),

			.SELF(gen[8658]),
			.cell_state(gen[8658])
		); 

/******************* CELL 8659 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8659 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8563]),
			.N(gen[8564]),
			.NE(gen[8565]),

			.O(gen[8658]),
			.E(gen[8660]),

			.SO(gen[8753]),
			.S(gen[8754]),
			.SE(gen[8755]),

			.SELF(gen[8659]),
			.cell_state(gen[8659])
		); 

/******************* CELL 8660 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8660 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8564]),
			.N(gen[8565]),
			.NE(gen[8566]),

			.O(gen[8659]),
			.E(gen[8661]),

			.SO(gen[8754]),
			.S(gen[8755]),
			.SE(gen[8756]),

			.SELF(gen[8660]),
			.cell_state(gen[8660])
		); 

/******************* CELL 8661 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8661 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8565]),
			.N(gen[8566]),
			.NE(gen[8567]),

			.O(gen[8660]),
			.E(gen[8662]),

			.SO(gen[8755]),
			.S(gen[8756]),
			.SE(gen[8757]),

			.SELF(gen[8661]),
			.cell_state(gen[8661])
		); 

/******************* CELL 8662 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8662 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8566]),
			.N(gen[8567]),
			.NE(gen[8568]),

			.O(gen[8661]),
			.E(gen[8663]),

			.SO(gen[8756]),
			.S(gen[8757]),
			.SE(gen[8758]),

			.SELF(gen[8662]),
			.cell_state(gen[8662])
		); 

/******************* CELL 8663 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8663 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8567]),
			.N(gen[8568]),
			.NE(gen[8569]),

			.O(gen[8662]),
			.E(gen[8664]),

			.SO(gen[8757]),
			.S(gen[8758]),
			.SE(gen[8759]),

			.SELF(gen[8663]),
			.cell_state(gen[8663])
		); 

/******************* CELL 8664 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8664 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8568]),
			.N(gen[8569]),
			.NE(gen[8570]),

			.O(gen[8663]),
			.E(gen[8665]),

			.SO(gen[8758]),
			.S(gen[8759]),
			.SE(gen[8760]),

			.SELF(gen[8664]),
			.cell_state(gen[8664])
		); 

/******************* CELL 8665 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8665 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8569]),
			.N(gen[8570]),
			.NE(gen[8571]),

			.O(gen[8664]),
			.E(gen[8666]),

			.SO(gen[8759]),
			.S(gen[8760]),
			.SE(gen[8761]),

			.SELF(gen[8665]),
			.cell_state(gen[8665])
		); 

/******************* CELL 8666 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8666 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8570]),
			.N(gen[8571]),
			.NE(gen[8572]),

			.O(gen[8665]),
			.E(gen[8667]),

			.SO(gen[8760]),
			.S(gen[8761]),
			.SE(gen[8762]),

			.SELF(gen[8666]),
			.cell_state(gen[8666])
		); 

/******************* CELL 8667 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8667 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8571]),
			.N(gen[8572]),
			.NE(gen[8573]),

			.O(gen[8666]),
			.E(gen[8668]),

			.SO(gen[8761]),
			.S(gen[8762]),
			.SE(gen[8763]),

			.SELF(gen[8667]),
			.cell_state(gen[8667])
		); 

/******************* CELL 8668 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8668 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8572]),
			.N(gen[8573]),
			.NE(gen[8574]),

			.O(gen[8667]),
			.E(gen[8669]),

			.SO(gen[8762]),
			.S(gen[8763]),
			.SE(gen[8764]),

			.SELF(gen[8668]),
			.cell_state(gen[8668])
		); 

/******************* CELL 8669 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8669 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8573]),
			.N(gen[8574]),
			.NE(gen[8575]),

			.O(gen[8668]),
			.E(gen[8670]),

			.SO(gen[8763]),
			.S(gen[8764]),
			.SE(gen[8765]),

			.SELF(gen[8669]),
			.cell_state(gen[8669])
		); 

/******************* CELL 8670 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8670 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8574]),
			.N(gen[8575]),
			.NE(gen[8576]),

			.O(gen[8669]),
			.E(gen[8671]),

			.SO(gen[8764]),
			.S(gen[8765]),
			.SE(gen[8766]),

			.SELF(gen[8670]),
			.cell_state(gen[8670])
		); 

/******************* CELL 8671 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8671 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8575]),
			.N(gen[8576]),
			.NE(gen[8577]),

			.O(gen[8670]),
			.E(gen[8672]),

			.SO(gen[8765]),
			.S(gen[8766]),
			.SE(gen[8767]),

			.SELF(gen[8671]),
			.cell_state(gen[8671])
		); 

/******************* CELL 8672 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8672 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8576]),
			.N(gen[8577]),
			.NE(gen[8578]),

			.O(gen[8671]),
			.E(gen[8673]),

			.SO(gen[8766]),
			.S(gen[8767]),
			.SE(gen[8768]),

			.SELF(gen[8672]),
			.cell_state(gen[8672])
		); 

/******************* CELL 8673 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8673 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8577]),
			.N(gen[8578]),
			.NE(gen[8579]),

			.O(gen[8672]),
			.E(gen[8674]),

			.SO(gen[8767]),
			.S(gen[8768]),
			.SE(gen[8769]),

			.SELF(gen[8673]),
			.cell_state(gen[8673])
		); 

/******************* CELL 8674 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8674 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8578]),
			.N(gen[8579]),
			.NE(gen[8580]),

			.O(gen[8673]),
			.E(gen[8675]),

			.SO(gen[8768]),
			.S(gen[8769]),
			.SE(gen[8770]),

			.SELF(gen[8674]),
			.cell_state(gen[8674])
		); 

/******************* CELL 8675 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8675 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8579]),
			.N(gen[8580]),
			.NE(gen[8581]),

			.O(gen[8674]),
			.E(gen[8676]),

			.SO(gen[8769]),
			.S(gen[8770]),
			.SE(gen[8771]),

			.SELF(gen[8675]),
			.cell_state(gen[8675])
		); 

/******************* CELL 8676 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8676 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8580]),
			.N(gen[8581]),
			.NE(gen[8582]),

			.O(gen[8675]),
			.E(gen[8677]),

			.SO(gen[8770]),
			.S(gen[8771]),
			.SE(gen[8772]),

			.SELF(gen[8676]),
			.cell_state(gen[8676])
		); 

/******************* CELL 8677 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8677 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8581]),
			.N(gen[8582]),
			.NE(gen[8583]),

			.O(gen[8676]),
			.E(gen[8678]),

			.SO(gen[8771]),
			.S(gen[8772]),
			.SE(gen[8773]),

			.SELF(gen[8677]),
			.cell_state(gen[8677])
		); 

/******************* CELL 8678 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8678 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8582]),
			.N(gen[8583]),
			.NE(gen[8584]),

			.O(gen[8677]),
			.E(gen[8679]),

			.SO(gen[8772]),
			.S(gen[8773]),
			.SE(gen[8774]),

			.SELF(gen[8678]),
			.cell_state(gen[8678])
		); 

/******************* CELL 8679 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8679 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8583]),
			.N(gen[8584]),
			.NE(gen[8585]),

			.O(gen[8678]),
			.E(gen[8680]),

			.SO(gen[8773]),
			.S(gen[8774]),
			.SE(gen[8775]),

			.SELF(gen[8679]),
			.cell_state(gen[8679])
		); 

/******************* CELL 8680 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8680 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8584]),
			.N(gen[8585]),
			.NE(gen[8586]),

			.O(gen[8679]),
			.E(gen[8681]),

			.SO(gen[8774]),
			.S(gen[8775]),
			.SE(gen[8776]),

			.SELF(gen[8680]),
			.cell_state(gen[8680])
		); 

/******************* CELL 8681 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8681 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8585]),
			.N(gen[8586]),
			.NE(gen[8587]),

			.O(gen[8680]),
			.E(gen[8682]),

			.SO(gen[8775]),
			.S(gen[8776]),
			.SE(gen[8777]),

			.SELF(gen[8681]),
			.cell_state(gen[8681])
		); 

/******************* CELL 8682 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8682 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8586]),
			.N(gen[8587]),
			.NE(gen[8588]),

			.O(gen[8681]),
			.E(gen[8683]),

			.SO(gen[8776]),
			.S(gen[8777]),
			.SE(gen[8778]),

			.SELF(gen[8682]),
			.cell_state(gen[8682])
		); 

/******************* CELL 8683 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8683 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8587]),
			.N(gen[8588]),
			.NE(gen[8589]),

			.O(gen[8682]),
			.E(gen[8684]),

			.SO(gen[8777]),
			.S(gen[8778]),
			.SE(gen[8779]),

			.SELF(gen[8683]),
			.cell_state(gen[8683])
		); 

/******************* CELL 8684 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8684 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8588]),
			.N(gen[8589]),
			.NE(gen[8590]),

			.O(gen[8683]),
			.E(gen[8685]),

			.SO(gen[8778]),
			.S(gen[8779]),
			.SE(gen[8780]),

			.SELF(gen[8684]),
			.cell_state(gen[8684])
		); 

/******************* CELL 8685 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8685 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8589]),
			.N(gen[8590]),
			.NE(gen[8591]),

			.O(gen[8684]),
			.E(gen[8686]),

			.SO(gen[8779]),
			.S(gen[8780]),
			.SE(gen[8781]),

			.SELF(gen[8685]),
			.cell_state(gen[8685])
		); 

/******************* CELL 8686 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8686 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8590]),
			.N(gen[8591]),
			.NE(gen[8592]),

			.O(gen[8685]),
			.E(gen[8687]),

			.SO(gen[8780]),
			.S(gen[8781]),
			.SE(gen[8782]),

			.SELF(gen[8686]),
			.cell_state(gen[8686])
		); 

/******************* CELL 8687 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8687 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8591]),
			.N(gen[8592]),
			.NE(gen[8593]),

			.O(gen[8686]),
			.E(gen[8688]),

			.SO(gen[8781]),
			.S(gen[8782]),
			.SE(gen[8783]),

			.SELF(gen[8687]),
			.cell_state(gen[8687])
		); 

/******************* CELL 8688 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8688 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8592]),
			.N(gen[8593]),
			.NE(gen[8594]),

			.O(gen[8687]),
			.E(gen[8689]),

			.SO(gen[8782]),
			.S(gen[8783]),
			.SE(gen[8784]),

			.SELF(gen[8688]),
			.cell_state(gen[8688])
		); 

/******************* CELL 8689 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8689 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8593]),
			.N(gen[8594]),
			.NE(gen[8595]),

			.O(gen[8688]),
			.E(gen[8690]),

			.SO(gen[8783]),
			.S(gen[8784]),
			.SE(gen[8785]),

			.SELF(gen[8689]),
			.cell_state(gen[8689])
		); 

/******************* CELL 8690 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8690 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8594]),
			.N(gen[8595]),
			.NE(gen[8596]),

			.O(gen[8689]),
			.E(gen[8691]),

			.SO(gen[8784]),
			.S(gen[8785]),
			.SE(gen[8786]),

			.SELF(gen[8690]),
			.cell_state(gen[8690])
		); 

/******************* CELL 8691 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8691 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8595]),
			.N(gen[8596]),
			.NE(gen[8597]),

			.O(gen[8690]),
			.E(gen[8692]),

			.SO(gen[8785]),
			.S(gen[8786]),
			.SE(gen[8787]),

			.SELF(gen[8691]),
			.cell_state(gen[8691])
		); 

/******************* CELL 8692 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8692 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8596]),
			.N(gen[8597]),
			.NE(gen[8598]),

			.O(gen[8691]),
			.E(gen[8693]),

			.SO(gen[8786]),
			.S(gen[8787]),
			.SE(gen[8788]),

			.SELF(gen[8692]),
			.cell_state(gen[8692])
		); 

/******************* CELL 8693 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8693 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8597]),
			.N(gen[8598]),
			.NE(gen[8599]),

			.O(gen[8692]),
			.E(gen[8694]),

			.SO(gen[8787]),
			.S(gen[8788]),
			.SE(gen[8789]),

			.SELF(gen[8693]),
			.cell_state(gen[8693])
		); 

/******************* CELL 8694 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8694 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8598]),
			.N(gen[8599]),
			.NE(gen[8600]),

			.O(gen[8693]),
			.E(gen[8695]),

			.SO(gen[8788]),
			.S(gen[8789]),
			.SE(gen[8790]),

			.SELF(gen[8694]),
			.cell_state(gen[8694])
		); 

/******************* CELL 8695 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8695 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8599]),
			.N(gen[8600]),
			.NE(gen[8601]),

			.O(gen[8694]),
			.E(gen[8696]),

			.SO(gen[8789]),
			.S(gen[8790]),
			.SE(gen[8791]),

			.SELF(gen[8695]),
			.cell_state(gen[8695])
		); 

/******************* CELL 8696 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8696 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8600]),
			.N(gen[8601]),
			.NE(gen[8602]),

			.O(gen[8695]),
			.E(gen[8697]),

			.SO(gen[8790]),
			.S(gen[8791]),
			.SE(gen[8792]),

			.SELF(gen[8696]),
			.cell_state(gen[8696])
		); 

/******************* CELL 8697 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8697 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8601]),
			.N(gen[8602]),
			.NE(gen[8603]),

			.O(gen[8696]),
			.E(gen[8698]),

			.SO(gen[8791]),
			.S(gen[8792]),
			.SE(gen[8793]),

			.SELF(gen[8697]),
			.cell_state(gen[8697])
		); 

/******************* CELL 8698 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8698 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8602]),
			.N(gen[8603]),
			.NE(gen[8604]),

			.O(gen[8697]),
			.E(gen[8699]),

			.SO(gen[8792]),
			.S(gen[8793]),
			.SE(gen[8794]),

			.SELF(gen[8698]),
			.cell_state(gen[8698])
		); 

/******************* CELL 8699 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8699 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8603]),
			.N(gen[8604]),
			.NE(gen[8605]),

			.O(gen[8698]),
			.E(gen[8700]),

			.SO(gen[8793]),
			.S(gen[8794]),
			.SE(gen[8795]),

			.SELF(gen[8699]),
			.cell_state(gen[8699])
		); 

/******************* CELL 8700 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8700 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8604]),
			.N(gen[8605]),
			.NE(gen[8606]),

			.O(gen[8699]),
			.E(gen[8701]),

			.SO(gen[8794]),
			.S(gen[8795]),
			.SE(gen[8796]),

			.SELF(gen[8700]),
			.cell_state(gen[8700])
		); 

/******************* CELL 8701 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8701 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8605]),
			.N(gen[8606]),
			.NE(gen[8607]),

			.O(gen[8700]),
			.E(gen[8702]),

			.SO(gen[8795]),
			.S(gen[8796]),
			.SE(gen[8797]),

			.SELF(gen[8701]),
			.cell_state(gen[8701])
		); 

/******************* CELL 8702 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8702 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8606]),
			.N(gen[8607]),
			.NE(gen[8608]),

			.O(gen[8701]),
			.E(gen[8703]),

			.SO(gen[8796]),
			.S(gen[8797]),
			.SE(gen[8798]),

			.SELF(gen[8702]),
			.cell_state(gen[8702])
		); 

/******************* CELL 8703 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8703 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8607]),
			.N(gen[8608]),
			.NE(gen[8609]),

			.O(gen[8702]),
			.E(gen[8704]),

			.SO(gen[8797]),
			.S(gen[8798]),
			.SE(gen[8799]),

			.SELF(gen[8703]),
			.cell_state(gen[8703])
		); 

/******************* CELL 8704 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8704 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8608]),
			.N(gen[8609]),
			.NE(gen[8610]),

			.O(gen[8703]),
			.E(gen[8705]),

			.SO(gen[8798]),
			.S(gen[8799]),
			.SE(gen[8800]),

			.SELF(gen[8704]),
			.cell_state(gen[8704])
		); 

/******************* CELL 8705 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8705 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8609]),
			.N(gen[8610]),
			.NE(gen[8611]),

			.O(gen[8704]),
			.E(gen[8706]),

			.SO(gen[8799]),
			.S(gen[8800]),
			.SE(gen[8801]),

			.SELF(gen[8705]),
			.cell_state(gen[8705])
		); 

/******************* CELL 8706 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8706 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8610]),
			.N(gen[8611]),
			.NE(gen[8612]),

			.O(gen[8705]),
			.E(gen[8707]),

			.SO(gen[8800]),
			.S(gen[8801]),
			.SE(gen[8802]),

			.SELF(gen[8706]),
			.cell_state(gen[8706])
		); 

/******************* CELL 8707 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8707 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8611]),
			.N(gen[8612]),
			.NE(gen[8613]),

			.O(gen[8706]),
			.E(gen[8708]),

			.SO(gen[8801]),
			.S(gen[8802]),
			.SE(gen[8803]),

			.SELF(gen[8707]),
			.cell_state(gen[8707])
		); 

/******************* CELL 8708 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8708 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8612]),
			.N(gen[8613]),
			.NE(gen[8614]),

			.O(gen[8707]),
			.E(gen[8709]),

			.SO(gen[8802]),
			.S(gen[8803]),
			.SE(gen[8804]),

			.SELF(gen[8708]),
			.cell_state(gen[8708])
		); 

/******************* CELL 8709 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8709 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8613]),
			.N(gen[8614]),
			.NE(gen[8615]),

			.O(gen[8708]),
			.E(gen[8710]),

			.SO(gen[8803]),
			.S(gen[8804]),
			.SE(gen[8805]),

			.SELF(gen[8709]),
			.cell_state(gen[8709])
		); 

/******************* CELL 8710 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8710 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8614]),
			.N(gen[8615]),
			.NE(gen[8616]),

			.O(gen[8709]),
			.E(gen[8711]),

			.SO(gen[8804]),
			.S(gen[8805]),
			.SE(gen[8806]),

			.SELF(gen[8710]),
			.cell_state(gen[8710])
		); 

/******************* CELL 8711 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8711 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8615]),
			.N(gen[8616]),
			.NE(gen[8617]),

			.O(gen[8710]),
			.E(gen[8712]),

			.SO(gen[8805]),
			.S(gen[8806]),
			.SE(gen[8807]),

			.SELF(gen[8711]),
			.cell_state(gen[8711])
		); 

/******************* CELL 8712 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8712 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8616]),
			.N(gen[8617]),
			.NE(gen[8618]),

			.O(gen[8711]),
			.E(gen[8713]),

			.SO(gen[8806]),
			.S(gen[8807]),
			.SE(gen[8808]),

			.SELF(gen[8712]),
			.cell_state(gen[8712])
		); 

/******************* CELL 8713 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8713 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8617]),
			.N(gen[8618]),
			.NE(gen[8619]),

			.O(gen[8712]),
			.E(gen[8714]),

			.SO(gen[8807]),
			.S(gen[8808]),
			.SE(gen[8809]),

			.SELF(gen[8713]),
			.cell_state(gen[8713])
		); 

/******************* CELL 8714 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8714 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8618]),
			.N(gen[8619]),
			.NE(gen[8620]),

			.O(gen[8713]),
			.E(gen[8715]),

			.SO(gen[8808]),
			.S(gen[8809]),
			.SE(gen[8810]),

			.SELF(gen[8714]),
			.cell_state(gen[8714])
		); 

/******************* CELL 8715 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8715 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8619]),
			.N(gen[8620]),
			.NE(gen[8621]),

			.O(gen[8714]),
			.E(gen[8716]),

			.SO(gen[8809]),
			.S(gen[8810]),
			.SE(gen[8811]),

			.SELF(gen[8715]),
			.cell_state(gen[8715])
		); 

/******************* CELL 8716 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8716 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8620]),
			.N(gen[8621]),
			.NE(gen[8622]),

			.O(gen[8715]),
			.E(gen[8717]),

			.SO(gen[8810]),
			.S(gen[8811]),
			.SE(gen[8812]),

			.SELF(gen[8716]),
			.cell_state(gen[8716])
		); 

/******************* CELL 8717 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8717 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8621]),
			.N(gen[8622]),
			.NE(gen[8623]),

			.O(gen[8716]),
			.E(gen[8718]),

			.SO(gen[8811]),
			.S(gen[8812]),
			.SE(gen[8813]),

			.SELF(gen[8717]),
			.cell_state(gen[8717])
		); 

/******************* CELL 8718 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8718 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8622]),
			.N(gen[8623]),
			.NE(gen[8624]),

			.O(gen[8717]),
			.E(gen[8719]),

			.SO(gen[8812]),
			.S(gen[8813]),
			.SE(gen[8814]),

			.SELF(gen[8718]),
			.cell_state(gen[8718])
		); 

/******************* CELL 8719 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8719 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8623]),
			.N(gen[8624]),
			.NE(gen[8625]),

			.O(gen[8718]),
			.E(gen[8720]),

			.SO(gen[8813]),
			.S(gen[8814]),
			.SE(gen[8815]),

			.SELF(gen[8719]),
			.cell_state(gen[8719])
		); 

/******************* CELL 8720 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8720 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8624]),
			.N(gen[8625]),
			.NE(gen[8626]),

			.O(gen[8719]),
			.E(gen[8721]),

			.SO(gen[8814]),
			.S(gen[8815]),
			.SE(gen[8816]),

			.SELF(gen[8720]),
			.cell_state(gen[8720])
		); 

/******************* CELL 8721 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8721 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8625]),
			.N(gen[8626]),
			.NE(gen[8627]),

			.O(gen[8720]),
			.E(gen[8722]),

			.SO(gen[8815]),
			.S(gen[8816]),
			.SE(gen[8817]),

			.SELF(gen[8721]),
			.cell_state(gen[8721])
		); 

/******************* CELL 8722 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8722 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8626]),
			.N(gen[8627]),
			.NE(gen[8628]),

			.O(gen[8721]),
			.E(gen[8723]),

			.SO(gen[8816]),
			.S(gen[8817]),
			.SE(gen[8818]),

			.SELF(gen[8722]),
			.cell_state(gen[8722])
		); 

/******************* CELL 8723 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8723 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8627]),
			.N(gen[8628]),
			.NE(gen[8629]),

			.O(gen[8722]),
			.E(gen[8724]),

			.SO(gen[8817]),
			.S(gen[8818]),
			.SE(gen[8819]),

			.SELF(gen[8723]),
			.cell_state(gen[8723])
		); 

/******************* CELL 8724 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8724 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8628]),
			.N(gen[8629]),
			.NE(gen[8630]),

			.O(gen[8723]),
			.E(gen[8725]),

			.SO(gen[8818]),
			.S(gen[8819]),
			.SE(gen[8820]),

			.SELF(gen[8724]),
			.cell_state(gen[8724])
		); 

/******************* CELL 8725 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8725 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8629]),
			.N(gen[8630]),
			.NE(gen[8631]),

			.O(gen[8724]),
			.E(gen[8726]),

			.SO(gen[8819]),
			.S(gen[8820]),
			.SE(gen[8821]),

			.SELF(gen[8725]),
			.cell_state(gen[8725])
		); 

/******************* CELL 8726 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8726 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8630]),
			.N(gen[8631]),
			.NE(gen[8632]),

			.O(gen[8725]),
			.E(gen[8727]),

			.SO(gen[8820]),
			.S(gen[8821]),
			.SE(gen[8822]),

			.SELF(gen[8726]),
			.cell_state(gen[8726])
		); 

/******************* CELL 8727 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8727 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8631]),
			.N(gen[8632]),
			.NE(gen[8633]),

			.O(gen[8726]),
			.E(gen[8728]),

			.SO(gen[8821]),
			.S(gen[8822]),
			.SE(gen[8823]),

			.SELF(gen[8727]),
			.cell_state(gen[8727])
		); 

/******************* CELL 8728 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8728 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8632]),
			.N(gen[8633]),
			.NE(gen[8634]),

			.O(gen[8727]),
			.E(gen[8729]),

			.SO(gen[8822]),
			.S(gen[8823]),
			.SE(gen[8824]),

			.SELF(gen[8728]),
			.cell_state(gen[8728])
		); 

/******************* CELL 8729 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8729 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8633]),
			.N(gen[8634]),
			.NE(gen[8635]),

			.O(gen[8728]),
			.E(gen[8730]),

			.SO(gen[8823]),
			.S(gen[8824]),
			.SE(gen[8825]),

			.SELF(gen[8729]),
			.cell_state(gen[8729])
		); 

/******************* CELL 8730 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8730 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8634]),
			.N(gen[8635]),
			.NE(gen[8636]),

			.O(gen[8729]),
			.E(gen[8731]),

			.SO(gen[8824]),
			.S(gen[8825]),
			.SE(gen[8826]),

			.SELF(gen[8730]),
			.cell_state(gen[8730])
		); 

/******************* CELL 8731 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8731 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8635]),
			.N(gen[8636]),
			.NE(gen[8637]),

			.O(gen[8730]),
			.E(gen[8732]),

			.SO(gen[8825]),
			.S(gen[8826]),
			.SE(gen[8827]),

			.SELF(gen[8731]),
			.cell_state(gen[8731])
		); 

/******************* CELL 8732 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8732 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8636]),
			.N(gen[8637]),
			.NE(gen[8638]),

			.O(gen[8731]),
			.E(gen[8733]),

			.SO(gen[8826]),
			.S(gen[8827]),
			.SE(gen[8828]),

			.SELF(gen[8732]),
			.cell_state(gen[8732])
		); 

/******************* CELL 8733 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8733 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8637]),
			.N(gen[8638]),
			.NE(gen[8639]),

			.O(gen[8732]),
			.E(gen[8734]),

			.SO(gen[8827]),
			.S(gen[8828]),
			.SE(gen[8829]),

			.SELF(gen[8733]),
			.cell_state(gen[8733])
		); 

/******************* CELL 8734 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8734 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8638]),
			.N(gen[8639]),
			.NE(gen[8640]),

			.O(gen[8733]),
			.E(gen[8735]),

			.SO(gen[8828]),
			.S(gen[8829]),
			.SE(gen[8830]),

			.SELF(gen[8734]),
			.cell_state(gen[8734])
		); 

/******************* CELL 8735 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8735 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8639]),
			.N(gen[8640]),
			.NE(gen[8641]),

			.O(gen[8734]),
			.E(gen[8736]),

			.SO(gen[8829]),
			.S(gen[8830]),
			.SE(gen[8831]),

			.SELF(gen[8735]),
			.cell_state(gen[8735])
		); 

/******************* CELL 8736 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8736 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8640]),
			.N(gen[8641]),
			.NE(gen[8642]),

			.O(gen[8735]),
			.E(gen[8737]),

			.SO(gen[8830]),
			.S(gen[8831]),
			.SE(gen[8832]),

			.SELF(gen[8736]),
			.cell_state(gen[8736])
		); 

/******************* CELL 8737 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8737 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8641]),
			.N(gen[8642]),
			.NE(gen[8643]),

			.O(gen[8736]),
			.E(gen[8738]),

			.SO(gen[8831]),
			.S(gen[8832]),
			.SE(gen[8833]),

			.SELF(gen[8737]),
			.cell_state(gen[8737])
		); 

/******************* CELL 8738 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8738 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8642]),
			.N(gen[8643]),
			.NE(gen[8644]),

			.O(gen[8737]),
			.E(gen[8739]),

			.SO(gen[8832]),
			.S(gen[8833]),
			.SE(gen[8834]),

			.SELF(gen[8738]),
			.cell_state(gen[8738])
		); 

/******************* CELL 8739 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8739 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8643]),
			.N(gen[8644]),
			.NE(gen[8643]),

			.O(gen[8738]),
			.E(gen[8738]),

			.SO(gen[8833]),
			.S(gen[8834]),
			.SE(gen[8833]),

			.SELF(gen[8739]),
			.cell_state(gen[8739])
		); 

/******************* CELL 8740 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8740 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8646]),
			.N(gen[8645]),
			.NE(gen[8646]),

			.O(gen[8741]),
			.E(gen[8741]),

			.SO(gen[8836]),
			.S(gen[8835]),
			.SE(gen[8836]),

			.SELF(gen[8740]),
			.cell_state(gen[8740])
		); 

/******************* CELL 8741 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8741 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8645]),
			.N(gen[8646]),
			.NE(gen[8647]),

			.O(gen[8740]),
			.E(gen[8742]),

			.SO(gen[8835]),
			.S(gen[8836]),
			.SE(gen[8837]),

			.SELF(gen[8741]),
			.cell_state(gen[8741])
		); 

/******************* CELL 8742 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8742 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8646]),
			.N(gen[8647]),
			.NE(gen[8648]),

			.O(gen[8741]),
			.E(gen[8743]),

			.SO(gen[8836]),
			.S(gen[8837]),
			.SE(gen[8838]),

			.SELF(gen[8742]),
			.cell_state(gen[8742])
		); 

/******************* CELL 8743 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8743 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8647]),
			.N(gen[8648]),
			.NE(gen[8649]),

			.O(gen[8742]),
			.E(gen[8744]),

			.SO(gen[8837]),
			.S(gen[8838]),
			.SE(gen[8839]),

			.SELF(gen[8743]),
			.cell_state(gen[8743])
		); 

/******************* CELL 8744 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8744 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8648]),
			.N(gen[8649]),
			.NE(gen[8650]),

			.O(gen[8743]),
			.E(gen[8745]),

			.SO(gen[8838]),
			.S(gen[8839]),
			.SE(gen[8840]),

			.SELF(gen[8744]),
			.cell_state(gen[8744])
		); 

/******************* CELL 8745 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8745 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8649]),
			.N(gen[8650]),
			.NE(gen[8651]),

			.O(gen[8744]),
			.E(gen[8746]),

			.SO(gen[8839]),
			.S(gen[8840]),
			.SE(gen[8841]),

			.SELF(gen[8745]),
			.cell_state(gen[8745])
		); 

/******************* CELL 8746 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8746 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8650]),
			.N(gen[8651]),
			.NE(gen[8652]),

			.O(gen[8745]),
			.E(gen[8747]),

			.SO(gen[8840]),
			.S(gen[8841]),
			.SE(gen[8842]),

			.SELF(gen[8746]),
			.cell_state(gen[8746])
		); 

/******************* CELL 8747 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8747 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8651]),
			.N(gen[8652]),
			.NE(gen[8653]),

			.O(gen[8746]),
			.E(gen[8748]),

			.SO(gen[8841]),
			.S(gen[8842]),
			.SE(gen[8843]),

			.SELF(gen[8747]),
			.cell_state(gen[8747])
		); 

/******************* CELL 8748 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8748 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8652]),
			.N(gen[8653]),
			.NE(gen[8654]),

			.O(gen[8747]),
			.E(gen[8749]),

			.SO(gen[8842]),
			.S(gen[8843]),
			.SE(gen[8844]),

			.SELF(gen[8748]),
			.cell_state(gen[8748])
		); 

/******************* CELL 8749 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8749 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8653]),
			.N(gen[8654]),
			.NE(gen[8655]),

			.O(gen[8748]),
			.E(gen[8750]),

			.SO(gen[8843]),
			.S(gen[8844]),
			.SE(gen[8845]),

			.SELF(gen[8749]),
			.cell_state(gen[8749])
		); 

/******************* CELL 8750 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8750 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8654]),
			.N(gen[8655]),
			.NE(gen[8656]),

			.O(gen[8749]),
			.E(gen[8751]),

			.SO(gen[8844]),
			.S(gen[8845]),
			.SE(gen[8846]),

			.SELF(gen[8750]),
			.cell_state(gen[8750])
		); 

/******************* CELL 8751 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8751 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8655]),
			.N(gen[8656]),
			.NE(gen[8657]),

			.O(gen[8750]),
			.E(gen[8752]),

			.SO(gen[8845]),
			.S(gen[8846]),
			.SE(gen[8847]),

			.SELF(gen[8751]),
			.cell_state(gen[8751])
		); 

/******************* CELL 8752 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8752 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8656]),
			.N(gen[8657]),
			.NE(gen[8658]),

			.O(gen[8751]),
			.E(gen[8753]),

			.SO(gen[8846]),
			.S(gen[8847]),
			.SE(gen[8848]),

			.SELF(gen[8752]),
			.cell_state(gen[8752])
		); 

/******************* CELL 8753 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8753 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8657]),
			.N(gen[8658]),
			.NE(gen[8659]),

			.O(gen[8752]),
			.E(gen[8754]),

			.SO(gen[8847]),
			.S(gen[8848]),
			.SE(gen[8849]),

			.SELF(gen[8753]),
			.cell_state(gen[8753])
		); 

/******************* CELL 8754 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8754 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8658]),
			.N(gen[8659]),
			.NE(gen[8660]),

			.O(gen[8753]),
			.E(gen[8755]),

			.SO(gen[8848]),
			.S(gen[8849]),
			.SE(gen[8850]),

			.SELF(gen[8754]),
			.cell_state(gen[8754])
		); 

/******************* CELL 8755 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8755 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8659]),
			.N(gen[8660]),
			.NE(gen[8661]),

			.O(gen[8754]),
			.E(gen[8756]),

			.SO(gen[8849]),
			.S(gen[8850]),
			.SE(gen[8851]),

			.SELF(gen[8755]),
			.cell_state(gen[8755])
		); 

/******************* CELL 8756 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8756 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8660]),
			.N(gen[8661]),
			.NE(gen[8662]),

			.O(gen[8755]),
			.E(gen[8757]),

			.SO(gen[8850]),
			.S(gen[8851]),
			.SE(gen[8852]),

			.SELF(gen[8756]),
			.cell_state(gen[8756])
		); 

/******************* CELL 8757 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8757 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8661]),
			.N(gen[8662]),
			.NE(gen[8663]),

			.O(gen[8756]),
			.E(gen[8758]),

			.SO(gen[8851]),
			.S(gen[8852]),
			.SE(gen[8853]),

			.SELF(gen[8757]),
			.cell_state(gen[8757])
		); 

/******************* CELL 8758 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8758 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8662]),
			.N(gen[8663]),
			.NE(gen[8664]),

			.O(gen[8757]),
			.E(gen[8759]),

			.SO(gen[8852]),
			.S(gen[8853]),
			.SE(gen[8854]),

			.SELF(gen[8758]),
			.cell_state(gen[8758])
		); 

/******************* CELL 8759 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8759 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8663]),
			.N(gen[8664]),
			.NE(gen[8665]),

			.O(gen[8758]),
			.E(gen[8760]),

			.SO(gen[8853]),
			.S(gen[8854]),
			.SE(gen[8855]),

			.SELF(gen[8759]),
			.cell_state(gen[8759])
		); 

/******************* CELL 8760 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8760 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8664]),
			.N(gen[8665]),
			.NE(gen[8666]),

			.O(gen[8759]),
			.E(gen[8761]),

			.SO(gen[8854]),
			.S(gen[8855]),
			.SE(gen[8856]),

			.SELF(gen[8760]),
			.cell_state(gen[8760])
		); 

/******************* CELL 8761 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8761 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8665]),
			.N(gen[8666]),
			.NE(gen[8667]),

			.O(gen[8760]),
			.E(gen[8762]),

			.SO(gen[8855]),
			.S(gen[8856]),
			.SE(gen[8857]),

			.SELF(gen[8761]),
			.cell_state(gen[8761])
		); 

/******************* CELL 8762 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8762 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8666]),
			.N(gen[8667]),
			.NE(gen[8668]),

			.O(gen[8761]),
			.E(gen[8763]),

			.SO(gen[8856]),
			.S(gen[8857]),
			.SE(gen[8858]),

			.SELF(gen[8762]),
			.cell_state(gen[8762])
		); 

/******************* CELL 8763 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8763 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8667]),
			.N(gen[8668]),
			.NE(gen[8669]),

			.O(gen[8762]),
			.E(gen[8764]),

			.SO(gen[8857]),
			.S(gen[8858]),
			.SE(gen[8859]),

			.SELF(gen[8763]),
			.cell_state(gen[8763])
		); 

/******************* CELL 8764 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8764 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8668]),
			.N(gen[8669]),
			.NE(gen[8670]),

			.O(gen[8763]),
			.E(gen[8765]),

			.SO(gen[8858]),
			.S(gen[8859]),
			.SE(gen[8860]),

			.SELF(gen[8764]),
			.cell_state(gen[8764])
		); 

/******************* CELL 8765 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8765 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8669]),
			.N(gen[8670]),
			.NE(gen[8671]),

			.O(gen[8764]),
			.E(gen[8766]),

			.SO(gen[8859]),
			.S(gen[8860]),
			.SE(gen[8861]),

			.SELF(gen[8765]),
			.cell_state(gen[8765])
		); 

/******************* CELL 8766 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8766 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8670]),
			.N(gen[8671]),
			.NE(gen[8672]),

			.O(gen[8765]),
			.E(gen[8767]),

			.SO(gen[8860]),
			.S(gen[8861]),
			.SE(gen[8862]),

			.SELF(gen[8766]),
			.cell_state(gen[8766])
		); 

/******************* CELL 8767 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8767 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8671]),
			.N(gen[8672]),
			.NE(gen[8673]),

			.O(gen[8766]),
			.E(gen[8768]),

			.SO(gen[8861]),
			.S(gen[8862]),
			.SE(gen[8863]),

			.SELF(gen[8767]),
			.cell_state(gen[8767])
		); 

/******************* CELL 8768 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8768 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8672]),
			.N(gen[8673]),
			.NE(gen[8674]),

			.O(gen[8767]),
			.E(gen[8769]),

			.SO(gen[8862]),
			.S(gen[8863]),
			.SE(gen[8864]),

			.SELF(gen[8768]),
			.cell_state(gen[8768])
		); 

/******************* CELL 8769 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8769 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8673]),
			.N(gen[8674]),
			.NE(gen[8675]),

			.O(gen[8768]),
			.E(gen[8770]),

			.SO(gen[8863]),
			.S(gen[8864]),
			.SE(gen[8865]),

			.SELF(gen[8769]),
			.cell_state(gen[8769])
		); 

/******************* CELL 8770 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8770 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8674]),
			.N(gen[8675]),
			.NE(gen[8676]),

			.O(gen[8769]),
			.E(gen[8771]),

			.SO(gen[8864]),
			.S(gen[8865]),
			.SE(gen[8866]),

			.SELF(gen[8770]),
			.cell_state(gen[8770])
		); 

/******************* CELL 8771 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8771 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8675]),
			.N(gen[8676]),
			.NE(gen[8677]),

			.O(gen[8770]),
			.E(gen[8772]),

			.SO(gen[8865]),
			.S(gen[8866]),
			.SE(gen[8867]),

			.SELF(gen[8771]),
			.cell_state(gen[8771])
		); 

/******************* CELL 8772 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8772 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8676]),
			.N(gen[8677]),
			.NE(gen[8678]),

			.O(gen[8771]),
			.E(gen[8773]),

			.SO(gen[8866]),
			.S(gen[8867]),
			.SE(gen[8868]),

			.SELF(gen[8772]),
			.cell_state(gen[8772])
		); 

/******************* CELL 8773 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8773 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8677]),
			.N(gen[8678]),
			.NE(gen[8679]),

			.O(gen[8772]),
			.E(gen[8774]),

			.SO(gen[8867]),
			.S(gen[8868]),
			.SE(gen[8869]),

			.SELF(gen[8773]),
			.cell_state(gen[8773])
		); 

/******************* CELL 8774 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8774 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8678]),
			.N(gen[8679]),
			.NE(gen[8680]),

			.O(gen[8773]),
			.E(gen[8775]),

			.SO(gen[8868]),
			.S(gen[8869]),
			.SE(gen[8870]),

			.SELF(gen[8774]),
			.cell_state(gen[8774])
		); 

/******************* CELL 8775 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8775 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8679]),
			.N(gen[8680]),
			.NE(gen[8681]),

			.O(gen[8774]),
			.E(gen[8776]),

			.SO(gen[8869]),
			.S(gen[8870]),
			.SE(gen[8871]),

			.SELF(gen[8775]),
			.cell_state(gen[8775])
		); 

/******************* CELL 8776 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8776 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8680]),
			.N(gen[8681]),
			.NE(gen[8682]),

			.O(gen[8775]),
			.E(gen[8777]),

			.SO(gen[8870]),
			.S(gen[8871]),
			.SE(gen[8872]),

			.SELF(gen[8776]),
			.cell_state(gen[8776])
		); 

/******************* CELL 8777 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8777 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8681]),
			.N(gen[8682]),
			.NE(gen[8683]),

			.O(gen[8776]),
			.E(gen[8778]),

			.SO(gen[8871]),
			.S(gen[8872]),
			.SE(gen[8873]),

			.SELF(gen[8777]),
			.cell_state(gen[8777])
		); 

/******************* CELL 8778 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8778 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8682]),
			.N(gen[8683]),
			.NE(gen[8684]),

			.O(gen[8777]),
			.E(gen[8779]),

			.SO(gen[8872]),
			.S(gen[8873]),
			.SE(gen[8874]),

			.SELF(gen[8778]),
			.cell_state(gen[8778])
		); 

/******************* CELL 8779 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8779 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8683]),
			.N(gen[8684]),
			.NE(gen[8685]),

			.O(gen[8778]),
			.E(gen[8780]),

			.SO(gen[8873]),
			.S(gen[8874]),
			.SE(gen[8875]),

			.SELF(gen[8779]),
			.cell_state(gen[8779])
		); 

/******************* CELL 8780 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8780 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8684]),
			.N(gen[8685]),
			.NE(gen[8686]),

			.O(gen[8779]),
			.E(gen[8781]),

			.SO(gen[8874]),
			.S(gen[8875]),
			.SE(gen[8876]),

			.SELF(gen[8780]),
			.cell_state(gen[8780])
		); 

/******************* CELL 8781 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8781 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8685]),
			.N(gen[8686]),
			.NE(gen[8687]),

			.O(gen[8780]),
			.E(gen[8782]),

			.SO(gen[8875]),
			.S(gen[8876]),
			.SE(gen[8877]),

			.SELF(gen[8781]),
			.cell_state(gen[8781])
		); 

/******************* CELL 8782 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8782 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8686]),
			.N(gen[8687]),
			.NE(gen[8688]),

			.O(gen[8781]),
			.E(gen[8783]),

			.SO(gen[8876]),
			.S(gen[8877]),
			.SE(gen[8878]),

			.SELF(gen[8782]),
			.cell_state(gen[8782])
		); 

/******************* CELL 8783 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8783 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8687]),
			.N(gen[8688]),
			.NE(gen[8689]),

			.O(gen[8782]),
			.E(gen[8784]),

			.SO(gen[8877]),
			.S(gen[8878]),
			.SE(gen[8879]),

			.SELF(gen[8783]),
			.cell_state(gen[8783])
		); 

/******************* CELL 8784 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8784 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8688]),
			.N(gen[8689]),
			.NE(gen[8690]),

			.O(gen[8783]),
			.E(gen[8785]),

			.SO(gen[8878]),
			.S(gen[8879]),
			.SE(gen[8880]),

			.SELF(gen[8784]),
			.cell_state(gen[8784])
		); 

/******************* CELL 8785 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8785 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8689]),
			.N(gen[8690]),
			.NE(gen[8691]),

			.O(gen[8784]),
			.E(gen[8786]),

			.SO(gen[8879]),
			.S(gen[8880]),
			.SE(gen[8881]),

			.SELF(gen[8785]),
			.cell_state(gen[8785])
		); 

/******************* CELL 8786 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8786 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8690]),
			.N(gen[8691]),
			.NE(gen[8692]),

			.O(gen[8785]),
			.E(gen[8787]),

			.SO(gen[8880]),
			.S(gen[8881]),
			.SE(gen[8882]),

			.SELF(gen[8786]),
			.cell_state(gen[8786])
		); 

/******************* CELL 8787 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8787 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8691]),
			.N(gen[8692]),
			.NE(gen[8693]),

			.O(gen[8786]),
			.E(gen[8788]),

			.SO(gen[8881]),
			.S(gen[8882]),
			.SE(gen[8883]),

			.SELF(gen[8787]),
			.cell_state(gen[8787])
		); 

/******************* CELL 8788 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8788 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8692]),
			.N(gen[8693]),
			.NE(gen[8694]),

			.O(gen[8787]),
			.E(gen[8789]),

			.SO(gen[8882]),
			.S(gen[8883]),
			.SE(gen[8884]),

			.SELF(gen[8788]),
			.cell_state(gen[8788])
		); 

/******************* CELL 8789 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8789 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8693]),
			.N(gen[8694]),
			.NE(gen[8695]),

			.O(gen[8788]),
			.E(gen[8790]),

			.SO(gen[8883]),
			.S(gen[8884]),
			.SE(gen[8885]),

			.SELF(gen[8789]),
			.cell_state(gen[8789])
		); 

/******************* CELL 8790 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8790 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8694]),
			.N(gen[8695]),
			.NE(gen[8696]),

			.O(gen[8789]),
			.E(gen[8791]),

			.SO(gen[8884]),
			.S(gen[8885]),
			.SE(gen[8886]),

			.SELF(gen[8790]),
			.cell_state(gen[8790])
		); 

/******************* CELL 8791 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8791 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8695]),
			.N(gen[8696]),
			.NE(gen[8697]),

			.O(gen[8790]),
			.E(gen[8792]),

			.SO(gen[8885]),
			.S(gen[8886]),
			.SE(gen[8887]),

			.SELF(gen[8791]),
			.cell_state(gen[8791])
		); 

/******************* CELL 8792 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8792 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8696]),
			.N(gen[8697]),
			.NE(gen[8698]),

			.O(gen[8791]),
			.E(gen[8793]),

			.SO(gen[8886]),
			.S(gen[8887]),
			.SE(gen[8888]),

			.SELF(gen[8792]),
			.cell_state(gen[8792])
		); 

/******************* CELL 8793 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8793 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8697]),
			.N(gen[8698]),
			.NE(gen[8699]),

			.O(gen[8792]),
			.E(gen[8794]),

			.SO(gen[8887]),
			.S(gen[8888]),
			.SE(gen[8889]),

			.SELF(gen[8793]),
			.cell_state(gen[8793])
		); 

/******************* CELL 8794 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8794 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8698]),
			.N(gen[8699]),
			.NE(gen[8700]),

			.O(gen[8793]),
			.E(gen[8795]),

			.SO(gen[8888]),
			.S(gen[8889]),
			.SE(gen[8890]),

			.SELF(gen[8794]),
			.cell_state(gen[8794])
		); 

/******************* CELL 8795 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8795 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8699]),
			.N(gen[8700]),
			.NE(gen[8701]),

			.O(gen[8794]),
			.E(gen[8796]),

			.SO(gen[8889]),
			.S(gen[8890]),
			.SE(gen[8891]),

			.SELF(gen[8795]),
			.cell_state(gen[8795])
		); 

/******************* CELL 8796 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8796 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8700]),
			.N(gen[8701]),
			.NE(gen[8702]),

			.O(gen[8795]),
			.E(gen[8797]),

			.SO(gen[8890]),
			.S(gen[8891]),
			.SE(gen[8892]),

			.SELF(gen[8796]),
			.cell_state(gen[8796])
		); 

/******************* CELL 8797 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8797 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8701]),
			.N(gen[8702]),
			.NE(gen[8703]),

			.O(gen[8796]),
			.E(gen[8798]),

			.SO(gen[8891]),
			.S(gen[8892]),
			.SE(gen[8893]),

			.SELF(gen[8797]),
			.cell_state(gen[8797])
		); 

/******************* CELL 8798 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8798 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8702]),
			.N(gen[8703]),
			.NE(gen[8704]),

			.O(gen[8797]),
			.E(gen[8799]),

			.SO(gen[8892]),
			.S(gen[8893]),
			.SE(gen[8894]),

			.SELF(gen[8798]),
			.cell_state(gen[8798])
		); 

/******************* CELL 8799 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8799 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8703]),
			.N(gen[8704]),
			.NE(gen[8705]),

			.O(gen[8798]),
			.E(gen[8800]),

			.SO(gen[8893]),
			.S(gen[8894]),
			.SE(gen[8895]),

			.SELF(gen[8799]),
			.cell_state(gen[8799])
		); 

/******************* CELL 8800 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8800 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8704]),
			.N(gen[8705]),
			.NE(gen[8706]),

			.O(gen[8799]),
			.E(gen[8801]),

			.SO(gen[8894]),
			.S(gen[8895]),
			.SE(gen[8896]),

			.SELF(gen[8800]),
			.cell_state(gen[8800])
		); 

/******************* CELL 8801 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8801 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8705]),
			.N(gen[8706]),
			.NE(gen[8707]),

			.O(gen[8800]),
			.E(gen[8802]),

			.SO(gen[8895]),
			.S(gen[8896]),
			.SE(gen[8897]),

			.SELF(gen[8801]),
			.cell_state(gen[8801])
		); 

/******************* CELL 8802 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8802 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8706]),
			.N(gen[8707]),
			.NE(gen[8708]),

			.O(gen[8801]),
			.E(gen[8803]),

			.SO(gen[8896]),
			.S(gen[8897]),
			.SE(gen[8898]),

			.SELF(gen[8802]),
			.cell_state(gen[8802])
		); 

/******************* CELL 8803 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8803 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8707]),
			.N(gen[8708]),
			.NE(gen[8709]),

			.O(gen[8802]),
			.E(gen[8804]),

			.SO(gen[8897]),
			.S(gen[8898]),
			.SE(gen[8899]),

			.SELF(gen[8803]),
			.cell_state(gen[8803])
		); 

/******************* CELL 8804 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8804 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8708]),
			.N(gen[8709]),
			.NE(gen[8710]),

			.O(gen[8803]),
			.E(gen[8805]),

			.SO(gen[8898]),
			.S(gen[8899]),
			.SE(gen[8900]),

			.SELF(gen[8804]),
			.cell_state(gen[8804])
		); 

/******************* CELL 8805 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8805 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8709]),
			.N(gen[8710]),
			.NE(gen[8711]),

			.O(gen[8804]),
			.E(gen[8806]),

			.SO(gen[8899]),
			.S(gen[8900]),
			.SE(gen[8901]),

			.SELF(gen[8805]),
			.cell_state(gen[8805])
		); 

/******************* CELL 8806 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8806 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8710]),
			.N(gen[8711]),
			.NE(gen[8712]),

			.O(gen[8805]),
			.E(gen[8807]),

			.SO(gen[8900]),
			.S(gen[8901]),
			.SE(gen[8902]),

			.SELF(gen[8806]),
			.cell_state(gen[8806])
		); 

/******************* CELL 8807 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8807 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8711]),
			.N(gen[8712]),
			.NE(gen[8713]),

			.O(gen[8806]),
			.E(gen[8808]),

			.SO(gen[8901]),
			.S(gen[8902]),
			.SE(gen[8903]),

			.SELF(gen[8807]),
			.cell_state(gen[8807])
		); 

/******************* CELL 8808 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8808 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8712]),
			.N(gen[8713]),
			.NE(gen[8714]),

			.O(gen[8807]),
			.E(gen[8809]),

			.SO(gen[8902]),
			.S(gen[8903]),
			.SE(gen[8904]),

			.SELF(gen[8808]),
			.cell_state(gen[8808])
		); 

/******************* CELL 8809 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8809 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8713]),
			.N(gen[8714]),
			.NE(gen[8715]),

			.O(gen[8808]),
			.E(gen[8810]),

			.SO(gen[8903]),
			.S(gen[8904]),
			.SE(gen[8905]),

			.SELF(gen[8809]),
			.cell_state(gen[8809])
		); 

/******************* CELL 8810 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8810 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8714]),
			.N(gen[8715]),
			.NE(gen[8716]),

			.O(gen[8809]),
			.E(gen[8811]),

			.SO(gen[8904]),
			.S(gen[8905]),
			.SE(gen[8906]),

			.SELF(gen[8810]),
			.cell_state(gen[8810])
		); 

/******************* CELL 8811 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8811 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8715]),
			.N(gen[8716]),
			.NE(gen[8717]),

			.O(gen[8810]),
			.E(gen[8812]),

			.SO(gen[8905]),
			.S(gen[8906]),
			.SE(gen[8907]),

			.SELF(gen[8811]),
			.cell_state(gen[8811])
		); 

/******************* CELL 8812 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8812 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8716]),
			.N(gen[8717]),
			.NE(gen[8718]),

			.O(gen[8811]),
			.E(gen[8813]),

			.SO(gen[8906]),
			.S(gen[8907]),
			.SE(gen[8908]),

			.SELF(gen[8812]),
			.cell_state(gen[8812])
		); 

/******************* CELL 8813 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8813 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8717]),
			.N(gen[8718]),
			.NE(gen[8719]),

			.O(gen[8812]),
			.E(gen[8814]),

			.SO(gen[8907]),
			.S(gen[8908]),
			.SE(gen[8909]),

			.SELF(gen[8813]),
			.cell_state(gen[8813])
		); 

/******************* CELL 8814 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8814 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8718]),
			.N(gen[8719]),
			.NE(gen[8720]),

			.O(gen[8813]),
			.E(gen[8815]),

			.SO(gen[8908]),
			.S(gen[8909]),
			.SE(gen[8910]),

			.SELF(gen[8814]),
			.cell_state(gen[8814])
		); 

/******************* CELL 8815 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8815 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8719]),
			.N(gen[8720]),
			.NE(gen[8721]),

			.O(gen[8814]),
			.E(gen[8816]),

			.SO(gen[8909]),
			.S(gen[8910]),
			.SE(gen[8911]),

			.SELF(gen[8815]),
			.cell_state(gen[8815])
		); 

/******************* CELL 8816 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8816 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8720]),
			.N(gen[8721]),
			.NE(gen[8722]),

			.O(gen[8815]),
			.E(gen[8817]),

			.SO(gen[8910]),
			.S(gen[8911]),
			.SE(gen[8912]),

			.SELF(gen[8816]),
			.cell_state(gen[8816])
		); 

/******************* CELL 8817 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8817 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8721]),
			.N(gen[8722]),
			.NE(gen[8723]),

			.O(gen[8816]),
			.E(gen[8818]),

			.SO(gen[8911]),
			.S(gen[8912]),
			.SE(gen[8913]),

			.SELF(gen[8817]),
			.cell_state(gen[8817])
		); 

/******************* CELL 8818 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8818 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8722]),
			.N(gen[8723]),
			.NE(gen[8724]),

			.O(gen[8817]),
			.E(gen[8819]),

			.SO(gen[8912]),
			.S(gen[8913]),
			.SE(gen[8914]),

			.SELF(gen[8818]),
			.cell_state(gen[8818])
		); 

/******************* CELL 8819 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8819 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8723]),
			.N(gen[8724]),
			.NE(gen[8725]),

			.O(gen[8818]),
			.E(gen[8820]),

			.SO(gen[8913]),
			.S(gen[8914]),
			.SE(gen[8915]),

			.SELF(gen[8819]),
			.cell_state(gen[8819])
		); 

/******************* CELL 8820 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8820 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8724]),
			.N(gen[8725]),
			.NE(gen[8726]),

			.O(gen[8819]),
			.E(gen[8821]),

			.SO(gen[8914]),
			.S(gen[8915]),
			.SE(gen[8916]),

			.SELF(gen[8820]),
			.cell_state(gen[8820])
		); 

/******************* CELL 8821 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8821 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8725]),
			.N(gen[8726]),
			.NE(gen[8727]),

			.O(gen[8820]),
			.E(gen[8822]),

			.SO(gen[8915]),
			.S(gen[8916]),
			.SE(gen[8917]),

			.SELF(gen[8821]),
			.cell_state(gen[8821])
		); 

/******************* CELL 8822 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8822 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8726]),
			.N(gen[8727]),
			.NE(gen[8728]),

			.O(gen[8821]),
			.E(gen[8823]),

			.SO(gen[8916]),
			.S(gen[8917]),
			.SE(gen[8918]),

			.SELF(gen[8822]),
			.cell_state(gen[8822])
		); 

/******************* CELL 8823 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8823 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8727]),
			.N(gen[8728]),
			.NE(gen[8729]),

			.O(gen[8822]),
			.E(gen[8824]),

			.SO(gen[8917]),
			.S(gen[8918]),
			.SE(gen[8919]),

			.SELF(gen[8823]),
			.cell_state(gen[8823])
		); 

/******************* CELL 8824 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8824 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8728]),
			.N(gen[8729]),
			.NE(gen[8730]),

			.O(gen[8823]),
			.E(gen[8825]),

			.SO(gen[8918]),
			.S(gen[8919]),
			.SE(gen[8920]),

			.SELF(gen[8824]),
			.cell_state(gen[8824])
		); 

/******************* CELL 8825 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8825 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8729]),
			.N(gen[8730]),
			.NE(gen[8731]),

			.O(gen[8824]),
			.E(gen[8826]),

			.SO(gen[8919]),
			.S(gen[8920]),
			.SE(gen[8921]),

			.SELF(gen[8825]),
			.cell_state(gen[8825])
		); 

/******************* CELL 8826 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8826 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8730]),
			.N(gen[8731]),
			.NE(gen[8732]),

			.O(gen[8825]),
			.E(gen[8827]),

			.SO(gen[8920]),
			.S(gen[8921]),
			.SE(gen[8922]),

			.SELF(gen[8826]),
			.cell_state(gen[8826])
		); 

/******************* CELL 8827 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8827 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8731]),
			.N(gen[8732]),
			.NE(gen[8733]),

			.O(gen[8826]),
			.E(gen[8828]),

			.SO(gen[8921]),
			.S(gen[8922]),
			.SE(gen[8923]),

			.SELF(gen[8827]),
			.cell_state(gen[8827])
		); 

/******************* CELL 8828 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8828 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8732]),
			.N(gen[8733]),
			.NE(gen[8734]),

			.O(gen[8827]),
			.E(gen[8829]),

			.SO(gen[8922]),
			.S(gen[8923]),
			.SE(gen[8924]),

			.SELF(gen[8828]),
			.cell_state(gen[8828])
		); 

/******************* CELL 8829 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8829 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8733]),
			.N(gen[8734]),
			.NE(gen[8735]),

			.O(gen[8828]),
			.E(gen[8830]),

			.SO(gen[8923]),
			.S(gen[8924]),
			.SE(gen[8925]),

			.SELF(gen[8829]),
			.cell_state(gen[8829])
		); 

/******************* CELL 8830 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8830 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8734]),
			.N(gen[8735]),
			.NE(gen[8736]),

			.O(gen[8829]),
			.E(gen[8831]),

			.SO(gen[8924]),
			.S(gen[8925]),
			.SE(gen[8926]),

			.SELF(gen[8830]),
			.cell_state(gen[8830])
		); 

/******************* CELL 8831 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8831 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8735]),
			.N(gen[8736]),
			.NE(gen[8737]),

			.O(gen[8830]),
			.E(gen[8832]),

			.SO(gen[8925]),
			.S(gen[8926]),
			.SE(gen[8927]),

			.SELF(gen[8831]),
			.cell_state(gen[8831])
		); 

/******************* CELL 8832 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8832 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8736]),
			.N(gen[8737]),
			.NE(gen[8738]),

			.O(gen[8831]),
			.E(gen[8833]),

			.SO(gen[8926]),
			.S(gen[8927]),
			.SE(gen[8928]),

			.SELF(gen[8832]),
			.cell_state(gen[8832])
		); 

/******************* CELL 8833 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8833 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8737]),
			.N(gen[8738]),
			.NE(gen[8739]),

			.O(gen[8832]),
			.E(gen[8834]),

			.SO(gen[8927]),
			.S(gen[8928]),
			.SE(gen[8929]),

			.SELF(gen[8833]),
			.cell_state(gen[8833])
		); 

/******************* CELL 8834 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8834 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8738]),
			.N(gen[8739]),
			.NE(gen[8738]),

			.O(gen[8833]),
			.E(gen[8833]),

			.SO(gen[8928]),
			.S(gen[8929]),
			.SE(gen[8928]),

			.SELF(gen[8834]),
			.cell_state(gen[8834])
		); 

/******************* CELL 8835 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8835 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8741]),
			.N(gen[8740]),
			.NE(gen[8741]),

			.O(gen[8836]),
			.E(gen[8836]),

			.SO(gen[8931]),
			.S(gen[8930]),
			.SE(gen[8931]),

			.SELF(gen[8835]),
			.cell_state(gen[8835])
		); 

/******************* CELL 8836 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8836 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8740]),
			.N(gen[8741]),
			.NE(gen[8742]),

			.O(gen[8835]),
			.E(gen[8837]),

			.SO(gen[8930]),
			.S(gen[8931]),
			.SE(gen[8932]),

			.SELF(gen[8836]),
			.cell_state(gen[8836])
		); 

/******************* CELL 8837 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8837 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8741]),
			.N(gen[8742]),
			.NE(gen[8743]),

			.O(gen[8836]),
			.E(gen[8838]),

			.SO(gen[8931]),
			.S(gen[8932]),
			.SE(gen[8933]),

			.SELF(gen[8837]),
			.cell_state(gen[8837])
		); 

/******************* CELL 8838 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8838 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8742]),
			.N(gen[8743]),
			.NE(gen[8744]),

			.O(gen[8837]),
			.E(gen[8839]),

			.SO(gen[8932]),
			.S(gen[8933]),
			.SE(gen[8934]),

			.SELF(gen[8838]),
			.cell_state(gen[8838])
		); 

/******************* CELL 8839 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8839 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8743]),
			.N(gen[8744]),
			.NE(gen[8745]),

			.O(gen[8838]),
			.E(gen[8840]),

			.SO(gen[8933]),
			.S(gen[8934]),
			.SE(gen[8935]),

			.SELF(gen[8839]),
			.cell_state(gen[8839])
		); 

/******************* CELL 8840 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8840 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8744]),
			.N(gen[8745]),
			.NE(gen[8746]),

			.O(gen[8839]),
			.E(gen[8841]),

			.SO(gen[8934]),
			.S(gen[8935]),
			.SE(gen[8936]),

			.SELF(gen[8840]),
			.cell_state(gen[8840])
		); 

/******************* CELL 8841 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8841 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8745]),
			.N(gen[8746]),
			.NE(gen[8747]),

			.O(gen[8840]),
			.E(gen[8842]),

			.SO(gen[8935]),
			.S(gen[8936]),
			.SE(gen[8937]),

			.SELF(gen[8841]),
			.cell_state(gen[8841])
		); 

/******************* CELL 8842 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8842 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8746]),
			.N(gen[8747]),
			.NE(gen[8748]),

			.O(gen[8841]),
			.E(gen[8843]),

			.SO(gen[8936]),
			.S(gen[8937]),
			.SE(gen[8938]),

			.SELF(gen[8842]),
			.cell_state(gen[8842])
		); 

/******************* CELL 8843 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8843 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8747]),
			.N(gen[8748]),
			.NE(gen[8749]),

			.O(gen[8842]),
			.E(gen[8844]),

			.SO(gen[8937]),
			.S(gen[8938]),
			.SE(gen[8939]),

			.SELF(gen[8843]),
			.cell_state(gen[8843])
		); 

/******************* CELL 8844 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8844 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8748]),
			.N(gen[8749]),
			.NE(gen[8750]),

			.O(gen[8843]),
			.E(gen[8845]),

			.SO(gen[8938]),
			.S(gen[8939]),
			.SE(gen[8940]),

			.SELF(gen[8844]),
			.cell_state(gen[8844])
		); 

/******************* CELL 8845 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8845 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8749]),
			.N(gen[8750]),
			.NE(gen[8751]),

			.O(gen[8844]),
			.E(gen[8846]),

			.SO(gen[8939]),
			.S(gen[8940]),
			.SE(gen[8941]),

			.SELF(gen[8845]),
			.cell_state(gen[8845])
		); 

/******************* CELL 8846 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8846 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8750]),
			.N(gen[8751]),
			.NE(gen[8752]),

			.O(gen[8845]),
			.E(gen[8847]),

			.SO(gen[8940]),
			.S(gen[8941]),
			.SE(gen[8942]),

			.SELF(gen[8846]),
			.cell_state(gen[8846])
		); 

/******************* CELL 8847 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8847 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8751]),
			.N(gen[8752]),
			.NE(gen[8753]),

			.O(gen[8846]),
			.E(gen[8848]),

			.SO(gen[8941]),
			.S(gen[8942]),
			.SE(gen[8943]),

			.SELF(gen[8847]),
			.cell_state(gen[8847])
		); 

/******************* CELL 8848 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8848 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8752]),
			.N(gen[8753]),
			.NE(gen[8754]),

			.O(gen[8847]),
			.E(gen[8849]),

			.SO(gen[8942]),
			.S(gen[8943]),
			.SE(gen[8944]),

			.SELF(gen[8848]),
			.cell_state(gen[8848])
		); 

/******************* CELL 8849 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8849 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8753]),
			.N(gen[8754]),
			.NE(gen[8755]),

			.O(gen[8848]),
			.E(gen[8850]),

			.SO(gen[8943]),
			.S(gen[8944]),
			.SE(gen[8945]),

			.SELF(gen[8849]),
			.cell_state(gen[8849])
		); 

/******************* CELL 8850 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8850 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8754]),
			.N(gen[8755]),
			.NE(gen[8756]),

			.O(gen[8849]),
			.E(gen[8851]),

			.SO(gen[8944]),
			.S(gen[8945]),
			.SE(gen[8946]),

			.SELF(gen[8850]),
			.cell_state(gen[8850])
		); 

/******************* CELL 8851 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8851 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8755]),
			.N(gen[8756]),
			.NE(gen[8757]),

			.O(gen[8850]),
			.E(gen[8852]),

			.SO(gen[8945]),
			.S(gen[8946]),
			.SE(gen[8947]),

			.SELF(gen[8851]),
			.cell_state(gen[8851])
		); 

/******************* CELL 8852 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8852 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8756]),
			.N(gen[8757]),
			.NE(gen[8758]),

			.O(gen[8851]),
			.E(gen[8853]),

			.SO(gen[8946]),
			.S(gen[8947]),
			.SE(gen[8948]),

			.SELF(gen[8852]),
			.cell_state(gen[8852])
		); 

/******************* CELL 8853 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8853 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8757]),
			.N(gen[8758]),
			.NE(gen[8759]),

			.O(gen[8852]),
			.E(gen[8854]),

			.SO(gen[8947]),
			.S(gen[8948]),
			.SE(gen[8949]),

			.SELF(gen[8853]),
			.cell_state(gen[8853])
		); 

/******************* CELL 8854 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8854 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8758]),
			.N(gen[8759]),
			.NE(gen[8760]),

			.O(gen[8853]),
			.E(gen[8855]),

			.SO(gen[8948]),
			.S(gen[8949]),
			.SE(gen[8950]),

			.SELF(gen[8854]),
			.cell_state(gen[8854])
		); 

/******************* CELL 8855 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8855 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8759]),
			.N(gen[8760]),
			.NE(gen[8761]),

			.O(gen[8854]),
			.E(gen[8856]),

			.SO(gen[8949]),
			.S(gen[8950]),
			.SE(gen[8951]),

			.SELF(gen[8855]),
			.cell_state(gen[8855])
		); 

/******************* CELL 8856 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8856 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8760]),
			.N(gen[8761]),
			.NE(gen[8762]),

			.O(gen[8855]),
			.E(gen[8857]),

			.SO(gen[8950]),
			.S(gen[8951]),
			.SE(gen[8952]),

			.SELF(gen[8856]),
			.cell_state(gen[8856])
		); 

/******************* CELL 8857 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8857 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8761]),
			.N(gen[8762]),
			.NE(gen[8763]),

			.O(gen[8856]),
			.E(gen[8858]),

			.SO(gen[8951]),
			.S(gen[8952]),
			.SE(gen[8953]),

			.SELF(gen[8857]),
			.cell_state(gen[8857])
		); 

/******************* CELL 8858 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8858 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8762]),
			.N(gen[8763]),
			.NE(gen[8764]),

			.O(gen[8857]),
			.E(gen[8859]),

			.SO(gen[8952]),
			.S(gen[8953]),
			.SE(gen[8954]),

			.SELF(gen[8858]),
			.cell_state(gen[8858])
		); 

/******************* CELL 8859 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8859 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8763]),
			.N(gen[8764]),
			.NE(gen[8765]),

			.O(gen[8858]),
			.E(gen[8860]),

			.SO(gen[8953]),
			.S(gen[8954]),
			.SE(gen[8955]),

			.SELF(gen[8859]),
			.cell_state(gen[8859])
		); 

/******************* CELL 8860 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8860 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8764]),
			.N(gen[8765]),
			.NE(gen[8766]),

			.O(gen[8859]),
			.E(gen[8861]),

			.SO(gen[8954]),
			.S(gen[8955]),
			.SE(gen[8956]),

			.SELF(gen[8860]),
			.cell_state(gen[8860])
		); 

/******************* CELL 8861 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8861 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8765]),
			.N(gen[8766]),
			.NE(gen[8767]),

			.O(gen[8860]),
			.E(gen[8862]),

			.SO(gen[8955]),
			.S(gen[8956]),
			.SE(gen[8957]),

			.SELF(gen[8861]),
			.cell_state(gen[8861])
		); 

/******************* CELL 8862 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8862 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8766]),
			.N(gen[8767]),
			.NE(gen[8768]),

			.O(gen[8861]),
			.E(gen[8863]),

			.SO(gen[8956]),
			.S(gen[8957]),
			.SE(gen[8958]),

			.SELF(gen[8862]),
			.cell_state(gen[8862])
		); 

/******************* CELL 8863 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8863 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8767]),
			.N(gen[8768]),
			.NE(gen[8769]),

			.O(gen[8862]),
			.E(gen[8864]),

			.SO(gen[8957]),
			.S(gen[8958]),
			.SE(gen[8959]),

			.SELF(gen[8863]),
			.cell_state(gen[8863])
		); 

/******************* CELL 8864 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8864 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8768]),
			.N(gen[8769]),
			.NE(gen[8770]),

			.O(gen[8863]),
			.E(gen[8865]),

			.SO(gen[8958]),
			.S(gen[8959]),
			.SE(gen[8960]),

			.SELF(gen[8864]),
			.cell_state(gen[8864])
		); 

/******************* CELL 8865 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8865 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8769]),
			.N(gen[8770]),
			.NE(gen[8771]),

			.O(gen[8864]),
			.E(gen[8866]),

			.SO(gen[8959]),
			.S(gen[8960]),
			.SE(gen[8961]),

			.SELF(gen[8865]),
			.cell_state(gen[8865])
		); 

/******************* CELL 8866 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8866 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8770]),
			.N(gen[8771]),
			.NE(gen[8772]),

			.O(gen[8865]),
			.E(gen[8867]),

			.SO(gen[8960]),
			.S(gen[8961]),
			.SE(gen[8962]),

			.SELF(gen[8866]),
			.cell_state(gen[8866])
		); 

/******************* CELL 8867 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8867 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8771]),
			.N(gen[8772]),
			.NE(gen[8773]),

			.O(gen[8866]),
			.E(gen[8868]),

			.SO(gen[8961]),
			.S(gen[8962]),
			.SE(gen[8963]),

			.SELF(gen[8867]),
			.cell_state(gen[8867])
		); 

/******************* CELL 8868 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8868 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8772]),
			.N(gen[8773]),
			.NE(gen[8774]),

			.O(gen[8867]),
			.E(gen[8869]),

			.SO(gen[8962]),
			.S(gen[8963]),
			.SE(gen[8964]),

			.SELF(gen[8868]),
			.cell_state(gen[8868])
		); 

/******************* CELL 8869 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8869 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8773]),
			.N(gen[8774]),
			.NE(gen[8775]),

			.O(gen[8868]),
			.E(gen[8870]),

			.SO(gen[8963]),
			.S(gen[8964]),
			.SE(gen[8965]),

			.SELF(gen[8869]),
			.cell_state(gen[8869])
		); 

/******************* CELL 8870 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8870 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8774]),
			.N(gen[8775]),
			.NE(gen[8776]),

			.O(gen[8869]),
			.E(gen[8871]),

			.SO(gen[8964]),
			.S(gen[8965]),
			.SE(gen[8966]),

			.SELF(gen[8870]),
			.cell_state(gen[8870])
		); 

/******************* CELL 8871 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8871 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8775]),
			.N(gen[8776]),
			.NE(gen[8777]),

			.O(gen[8870]),
			.E(gen[8872]),

			.SO(gen[8965]),
			.S(gen[8966]),
			.SE(gen[8967]),

			.SELF(gen[8871]),
			.cell_state(gen[8871])
		); 

/******************* CELL 8872 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8872 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8776]),
			.N(gen[8777]),
			.NE(gen[8778]),

			.O(gen[8871]),
			.E(gen[8873]),

			.SO(gen[8966]),
			.S(gen[8967]),
			.SE(gen[8968]),

			.SELF(gen[8872]),
			.cell_state(gen[8872])
		); 

/******************* CELL 8873 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8873 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8777]),
			.N(gen[8778]),
			.NE(gen[8779]),

			.O(gen[8872]),
			.E(gen[8874]),

			.SO(gen[8967]),
			.S(gen[8968]),
			.SE(gen[8969]),

			.SELF(gen[8873]),
			.cell_state(gen[8873])
		); 

/******************* CELL 8874 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8874 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8778]),
			.N(gen[8779]),
			.NE(gen[8780]),

			.O(gen[8873]),
			.E(gen[8875]),

			.SO(gen[8968]),
			.S(gen[8969]),
			.SE(gen[8970]),

			.SELF(gen[8874]),
			.cell_state(gen[8874])
		); 

/******************* CELL 8875 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8875 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8779]),
			.N(gen[8780]),
			.NE(gen[8781]),

			.O(gen[8874]),
			.E(gen[8876]),

			.SO(gen[8969]),
			.S(gen[8970]),
			.SE(gen[8971]),

			.SELF(gen[8875]),
			.cell_state(gen[8875])
		); 

/******************* CELL 8876 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8876 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8780]),
			.N(gen[8781]),
			.NE(gen[8782]),

			.O(gen[8875]),
			.E(gen[8877]),

			.SO(gen[8970]),
			.S(gen[8971]),
			.SE(gen[8972]),

			.SELF(gen[8876]),
			.cell_state(gen[8876])
		); 

/******************* CELL 8877 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8877 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8781]),
			.N(gen[8782]),
			.NE(gen[8783]),

			.O(gen[8876]),
			.E(gen[8878]),

			.SO(gen[8971]),
			.S(gen[8972]),
			.SE(gen[8973]),

			.SELF(gen[8877]),
			.cell_state(gen[8877])
		); 

/******************* CELL 8878 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8878 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8782]),
			.N(gen[8783]),
			.NE(gen[8784]),

			.O(gen[8877]),
			.E(gen[8879]),

			.SO(gen[8972]),
			.S(gen[8973]),
			.SE(gen[8974]),

			.SELF(gen[8878]),
			.cell_state(gen[8878])
		); 

/******************* CELL 8879 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8879 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8783]),
			.N(gen[8784]),
			.NE(gen[8785]),

			.O(gen[8878]),
			.E(gen[8880]),

			.SO(gen[8973]),
			.S(gen[8974]),
			.SE(gen[8975]),

			.SELF(gen[8879]),
			.cell_state(gen[8879])
		); 

/******************* CELL 8880 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8880 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8784]),
			.N(gen[8785]),
			.NE(gen[8786]),

			.O(gen[8879]),
			.E(gen[8881]),

			.SO(gen[8974]),
			.S(gen[8975]),
			.SE(gen[8976]),

			.SELF(gen[8880]),
			.cell_state(gen[8880])
		); 

/******************* CELL 8881 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8881 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8785]),
			.N(gen[8786]),
			.NE(gen[8787]),

			.O(gen[8880]),
			.E(gen[8882]),

			.SO(gen[8975]),
			.S(gen[8976]),
			.SE(gen[8977]),

			.SELF(gen[8881]),
			.cell_state(gen[8881])
		); 

/******************* CELL 8882 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8882 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8786]),
			.N(gen[8787]),
			.NE(gen[8788]),

			.O(gen[8881]),
			.E(gen[8883]),

			.SO(gen[8976]),
			.S(gen[8977]),
			.SE(gen[8978]),

			.SELF(gen[8882]),
			.cell_state(gen[8882])
		); 

/******************* CELL 8883 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8883 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8787]),
			.N(gen[8788]),
			.NE(gen[8789]),

			.O(gen[8882]),
			.E(gen[8884]),

			.SO(gen[8977]),
			.S(gen[8978]),
			.SE(gen[8979]),

			.SELF(gen[8883]),
			.cell_state(gen[8883])
		); 

/******************* CELL 8884 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8884 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8788]),
			.N(gen[8789]),
			.NE(gen[8790]),

			.O(gen[8883]),
			.E(gen[8885]),

			.SO(gen[8978]),
			.S(gen[8979]),
			.SE(gen[8980]),

			.SELF(gen[8884]),
			.cell_state(gen[8884])
		); 

/******************* CELL 8885 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8885 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8789]),
			.N(gen[8790]),
			.NE(gen[8791]),

			.O(gen[8884]),
			.E(gen[8886]),

			.SO(gen[8979]),
			.S(gen[8980]),
			.SE(gen[8981]),

			.SELF(gen[8885]),
			.cell_state(gen[8885])
		); 

/******************* CELL 8886 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8886 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8790]),
			.N(gen[8791]),
			.NE(gen[8792]),

			.O(gen[8885]),
			.E(gen[8887]),

			.SO(gen[8980]),
			.S(gen[8981]),
			.SE(gen[8982]),

			.SELF(gen[8886]),
			.cell_state(gen[8886])
		); 

/******************* CELL 8887 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8887 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8791]),
			.N(gen[8792]),
			.NE(gen[8793]),

			.O(gen[8886]),
			.E(gen[8888]),

			.SO(gen[8981]),
			.S(gen[8982]),
			.SE(gen[8983]),

			.SELF(gen[8887]),
			.cell_state(gen[8887])
		); 

/******************* CELL 8888 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8888 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8792]),
			.N(gen[8793]),
			.NE(gen[8794]),

			.O(gen[8887]),
			.E(gen[8889]),

			.SO(gen[8982]),
			.S(gen[8983]),
			.SE(gen[8984]),

			.SELF(gen[8888]),
			.cell_state(gen[8888])
		); 

/******************* CELL 8889 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8889 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8793]),
			.N(gen[8794]),
			.NE(gen[8795]),

			.O(gen[8888]),
			.E(gen[8890]),

			.SO(gen[8983]),
			.S(gen[8984]),
			.SE(gen[8985]),

			.SELF(gen[8889]),
			.cell_state(gen[8889])
		); 

/******************* CELL 8890 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8890 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8794]),
			.N(gen[8795]),
			.NE(gen[8796]),

			.O(gen[8889]),
			.E(gen[8891]),

			.SO(gen[8984]),
			.S(gen[8985]),
			.SE(gen[8986]),

			.SELF(gen[8890]),
			.cell_state(gen[8890])
		); 

/******************* CELL 8891 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8891 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8795]),
			.N(gen[8796]),
			.NE(gen[8797]),

			.O(gen[8890]),
			.E(gen[8892]),

			.SO(gen[8985]),
			.S(gen[8986]),
			.SE(gen[8987]),

			.SELF(gen[8891]),
			.cell_state(gen[8891])
		); 

/******************* CELL 8892 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8892 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8796]),
			.N(gen[8797]),
			.NE(gen[8798]),

			.O(gen[8891]),
			.E(gen[8893]),

			.SO(gen[8986]),
			.S(gen[8987]),
			.SE(gen[8988]),

			.SELF(gen[8892]),
			.cell_state(gen[8892])
		); 

/******************* CELL 8893 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8893 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8797]),
			.N(gen[8798]),
			.NE(gen[8799]),

			.O(gen[8892]),
			.E(gen[8894]),

			.SO(gen[8987]),
			.S(gen[8988]),
			.SE(gen[8989]),

			.SELF(gen[8893]),
			.cell_state(gen[8893])
		); 

/******************* CELL 8894 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8894 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8798]),
			.N(gen[8799]),
			.NE(gen[8800]),

			.O(gen[8893]),
			.E(gen[8895]),

			.SO(gen[8988]),
			.S(gen[8989]),
			.SE(gen[8990]),

			.SELF(gen[8894]),
			.cell_state(gen[8894])
		); 

/******************* CELL 8895 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8895 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8799]),
			.N(gen[8800]),
			.NE(gen[8801]),

			.O(gen[8894]),
			.E(gen[8896]),

			.SO(gen[8989]),
			.S(gen[8990]),
			.SE(gen[8991]),

			.SELF(gen[8895]),
			.cell_state(gen[8895])
		); 

/******************* CELL 8896 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8896 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8800]),
			.N(gen[8801]),
			.NE(gen[8802]),

			.O(gen[8895]),
			.E(gen[8897]),

			.SO(gen[8990]),
			.S(gen[8991]),
			.SE(gen[8992]),

			.SELF(gen[8896]),
			.cell_state(gen[8896])
		); 

/******************* CELL 8897 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8897 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8801]),
			.N(gen[8802]),
			.NE(gen[8803]),

			.O(gen[8896]),
			.E(gen[8898]),

			.SO(gen[8991]),
			.S(gen[8992]),
			.SE(gen[8993]),

			.SELF(gen[8897]),
			.cell_state(gen[8897])
		); 

/******************* CELL 8898 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8898 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8802]),
			.N(gen[8803]),
			.NE(gen[8804]),

			.O(gen[8897]),
			.E(gen[8899]),

			.SO(gen[8992]),
			.S(gen[8993]),
			.SE(gen[8994]),

			.SELF(gen[8898]),
			.cell_state(gen[8898])
		); 

/******************* CELL 8899 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8899 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8803]),
			.N(gen[8804]),
			.NE(gen[8805]),

			.O(gen[8898]),
			.E(gen[8900]),

			.SO(gen[8993]),
			.S(gen[8994]),
			.SE(gen[8995]),

			.SELF(gen[8899]),
			.cell_state(gen[8899])
		); 

/******************* CELL 8900 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8900 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8804]),
			.N(gen[8805]),
			.NE(gen[8806]),

			.O(gen[8899]),
			.E(gen[8901]),

			.SO(gen[8994]),
			.S(gen[8995]),
			.SE(gen[8996]),

			.SELF(gen[8900]),
			.cell_state(gen[8900])
		); 

/******************* CELL 8901 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8901 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8805]),
			.N(gen[8806]),
			.NE(gen[8807]),

			.O(gen[8900]),
			.E(gen[8902]),

			.SO(gen[8995]),
			.S(gen[8996]),
			.SE(gen[8997]),

			.SELF(gen[8901]),
			.cell_state(gen[8901])
		); 

/******************* CELL 8902 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8902 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8806]),
			.N(gen[8807]),
			.NE(gen[8808]),

			.O(gen[8901]),
			.E(gen[8903]),

			.SO(gen[8996]),
			.S(gen[8997]),
			.SE(gen[8998]),

			.SELF(gen[8902]),
			.cell_state(gen[8902])
		); 

/******************* CELL 8903 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8903 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8807]),
			.N(gen[8808]),
			.NE(gen[8809]),

			.O(gen[8902]),
			.E(gen[8904]),

			.SO(gen[8997]),
			.S(gen[8998]),
			.SE(gen[8999]),

			.SELF(gen[8903]),
			.cell_state(gen[8903])
		); 

/******************* CELL 8904 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8904 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8808]),
			.N(gen[8809]),
			.NE(gen[8810]),

			.O(gen[8903]),
			.E(gen[8905]),

			.SO(gen[8998]),
			.S(gen[8999]),
			.SE(gen[9000]),

			.SELF(gen[8904]),
			.cell_state(gen[8904])
		); 

/******************* CELL 8905 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8905 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8809]),
			.N(gen[8810]),
			.NE(gen[8811]),

			.O(gen[8904]),
			.E(gen[8906]),

			.SO(gen[8999]),
			.S(gen[9000]),
			.SE(gen[9001]),

			.SELF(gen[8905]),
			.cell_state(gen[8905])
		); 

/******************* CELL 8906 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8906 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8810]),
			.N(gen[8811]),
			.NE(gen[8812]),

			.O(gen[8905]),
			.E(gen[8907]),

			.SO(gen[9000]),
			.S(gen[9001]),
			.SE(gen[9002]),

			.SELF(gen[8906]),
			.cell_state(gen[8906])
		); 

/******************* CELL 8907 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8907 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8811]),
			.N(gen[8812]),
			.NE(gen[8813]),

			.O(gen[8906]),
			.E(gen[8908]),

			.SO(gen[9001]),
			.S(gen[9002]),
			.SE(gen[9003]),

			.SELF(gen[8907]),
			.cell_state(gen[8907])
		); 

/******************* CELL 8908 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8908 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8812]),
			.N(gen[8813]),
			.NE(gen[8814]),

			.O(gen[8907]),
			.E(gen[8909]),

			.SO(gen[9002]),
			.S(gen[9003]),
			.SE(gen[9004]),

			.SELF(gen[8908]),
			.cell_state(gen[8908])
		); 

/******************* CELL 8909 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8909 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8813]),
			.N(gen[8814]),
			.NE(gen[8815]),

			.O(gen[8908]),
			.E(gen[8910]),

			.SO(gen[9003]),
			.S(gen[9004]),
			.SE(gen[9005]),

			.SELF(gen[8909]),
			.cell_state(gen[8909])
		); 

/******************* CELL 8910 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8910 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8814]),
			.N(gen[8815]),
			.NE(gen[8816]),

			.O(gen[8909]),
			.E(gen[8911]),

			.SO(gen[9004]),
			.S(gen[9005]),
			.SE(gen[9006]),

			.SELF(gen[8910]),
			.cell_state(gen[8910])
		); 

/******************* CELL 8911 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8911 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8815]),
			.N(gen[8816]),
			.NE(gen[8817]),

			.O(gen[8910]),
			.E(gen[8912]),

			.SO(gen[9005]),
			.S(gen[9006]),
			.SE(gen[9007]),

			.SELF(gen[8911]),
			.cell_state(gen[8911])
		); 

/******************* CELL 8912 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8912 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8816]),
			.N(gen[8817]),
			.NE(gen[8818]),

			.O(gen[8911]),
			.E(gen[8913]),

			.SO(gen[9006]),
			.S(gen[9007]),
			.SE(gen[9008]),

			.SELF(gen[8912]),
			.cell_state(gen[8912])
		); 

/******************* CELL 8913 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8913 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8817]),
			.N(gen[8818]),
			.NE(gen[8819]),

			.O(gen[8912]),
			.E(gen[8914]),

			.SO(gen[9007]),
			.S(gen[9008]),
			.SE(gen[9009]),

			.SELF(gen[8913]),
			.cell_state(gen[8913])
		); 

/******************* CELL 8914 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8914 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8818]),
			.N(gen[8819]),
			.NE(gen[8820]),

			.O(gen[8913]),
			.E(gen[8915]),

			.SO(gen[9008]),
			.S(gen[9009]),
			.SE(gen[9010]),

			.SELF(gen[8914]),
			.cell_state(gen[8914])
		); 

/******************* CELL 8915 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8915 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8819]),
			.N(gen[8820]),
			.NE(gen[8821]),

			.O(gen[8914]),
			.E(gen[8916]),

			.SO(gen[9009]),
			.S(gen[9010]),
			.SE(gen[9011]),

			.SELF(gen[8915]),
			.cell_state(gen[8915])
		); 

/******************* CELL 8916 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8916 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8820]),
			.N(gen[8821]),
			.NE(gen[8822]),

			.O(gen[8915]),
			.E(gen[8917]),

			.SO(gen[9010]),
			.S(gen[9011]),
			.SE(gen[9012]),

			.SELF(gen[8916]),
			.cell_state(gen[8916])
		); 

/******************* CELL 8917 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8917 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8821]),
			.N(gen[8822]),
			.NE(gen[8823]),

			.O(gen[8916]),
			.E(gen[8918]),

			.SO(gen[9011]),
			.S(gen[9012]),
			.SE(gen[9013]),

			.SELF(gen[8917]),
			.cell_state(gen[8917])
		); 

/******************* CELL 8918 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8918 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8822]),
			.N(gen[8823]),
			.NE(gen[8824]),

			.O(gen[8917]),
			.E(gen[8919]),

			.SO(gen[9012]),
			.S(gen[9013]),
			.SE(gen[9014]),

			.SELF(gen[8918]),
			.cell_state(gen[8918])
		); 

/******************* CELL 8919 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8919 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8823]),
			.N(gen[8824]),
			.NE(gen[8825]),

			.O(gen[8918]),
			.E(gen[8920]),

			.SO(gen[9013]),
			.S(gen[9014]),
			.SE(gen[9015]),

			.SELF(gen[8919]),
			.cell_state(gen[8919])
		); 

/******************* CELL 8920 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8920 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8824]),
			.N(gen[8825]),
			.NE(gen[8826]),

			.O(gen[8919]),
			.E(gen[8921]),

			.SO(gen[9014]),
			.S(gen[9015]),
			.SE(gen[9016]),

			.SELF(gen[8920]),
			.cell_state(gen[8920])
		); 

/******************* CELL 8921 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8921 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8825]),
			.N(gen[8826]),
			.NE(gen[8827]),

			.O(gen[8920]),
			.E(gen[8922]),

			.SO(gen[9015]),
			.S(gen[9016]),
			.SE(gen[9017]),

			.SELF(gen[8921]),
			.cell_state(gen[8921])
		); 

/******************* CELL 8922 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8922 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8826]),
			.N(gen[8827]),
			.NE(gen[8828]),

			.O(gen[8921]),
			.E(gen[8923]),

			.SO(gen[9016]),
			.S(gen[9017]),
			.SE(gen[9018]),

			.SELF(gen[8922]),
			.cell_state(gen[8922])
		); 

/******************* CELL 8923 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8923 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8827]),
			.N(gen[8828]),
			.NE(gen[8829]),

			.O(gen[8922]),
			.E(gen[8924]),

			.SO(gen[9017]),
			.S(gen[9018]),
			.SE(gen[9019]),

			.SELF(gen[8923]),
			.cell_state(gen[8923])
		); 

/******************* CELL 8924 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8924 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8828]),
			.N(gen[8829]),
			.NE(gen[8830]),

			.O(gen[8923]),
			.E(gen[8925]),

			.SO(gen[9018]),
			.S(gen[9019]),
			.SE(gen[9020]),

			.SELF(gen[8924]),
			.cell_state(gen[8924])
		); 

/******************* CELL 8925 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8925 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8829]),
			.N(gen[8830]),
			.NE(gen[8831]),

			.O(gen[8924]),
			.E(gen[8926]),

			.SO(gen[9019]),
			.S(gen[9020]),
			.SE(gen[9021]),

			.SELF(gen[8925]),
			.cell_state(gen[8925])
		); 

/******************* CELL 8926 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8926 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8830]),
			.N(gen[8831]),
			.NE(gen[8832]),

			.O(gen[8925]),
			.E(gen[8927]),

			.SO(gen[9020]),
			.S(gen[9021]),
			.SE(gen[9022]),

			.SELF(gen[8926]),
			.cell_state(gen[8926])
		); 

/******************* CELL 8927 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8927 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8831]),
			.N(gen[8832]),
			.NE(gen[8833]),

			.O(gen[8926]),
			.E(gen[8928]),

			.SO(gen[9021]),
			.S(gen[9022]),
			.SE(gen[9023]),

			.SELF(gen[8927]),
			.cell_state(gen[8927])
		); 

/******************* CELL 8928 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8928 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8832]),
			.N(gen[8833]),
			.NE(gen[8834]),

			.O(gen[8927]),
			.E(gen[8929]),

			.SO(gen[9022]),
			.S(gen[9023]),
			.SE(gen[9024]),

			.SELF(gen[8928]),
			.cell_state(gen[8928])
		); 

/******************* CELL 8929 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell8929 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8833]),
			.N(gen[8834]),
			.NE(gen[8833]),

			.O(gen[8928]),
			.E(gen[8928]),

			.SO(gen[9023]),
			.S(gen[9024]),
			.SE(gen[9023]),

			.SELF(gen[8929]),
			.cell_state(gen[8929])
		); 

/******************* CELL 8930 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8930 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8836]),
			.N(gen[8835]),
			.NE(gen[8836]),

			.O(gen[8931]),
			.E(gen[8931]),

			.SO(gen[8836]),
			.S(gen[8835]),
			.SE(gen[8836]),

			.SELF(gen[8930]),
			.cell_state(gen[8930])
		); 

/******************* CELL 8931 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8931 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8835]),
			.N(gen[8836]),
			.NE(gen[8837]),

			.O(gen[8930]),
			.E(gen[8932]),

			.SO(gen[8835]),
			.S(gen[8836]),
			.SE(gen[8837]),

			.SELF(gen[8931]),
			.cell_state(gen[8931])
		); 

/******************* CELL 8932 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8932 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8836]),
			.N(gen[8837]),
			.NE(gen[8838]),

			.O(gen[8931]),
			.E(gen[8933]),

			.SO(gen[8836]),
			.S(gen[8837]),
			.SE(gen[8838]),

			.SELF(gen[8932]),
			.cell_state(gen[8932])
		); 

/******************* CELL 8933 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8933 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8837]),
			.N(gen[8838]),
			.NE(gen[8839]),

			.O(gen[8932]),
			.E(gen[8934]),

			.SO(gen[8837]),
			.S(gen[8838]),
			.SE(gen[8839]),

			.SELF(gen[8933]),
			.cell_state(gen[8933])
		); 

/******************* CELL 8934 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8934 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8838]),
			.N(gen[8839]),
			.NE(gen[8840]),

			.O(gen[8933]),
			.E(gen[8935]),

			.SO(gen[8838]),
			.S(gen[8839]),
			.SE(gen[8840]),

			.SELF(gen[8934]),
			.cell_state(gen[8934])
		); 

/******************* CELL 8935 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8935 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8839]),
			.N(gen[8840]),
			.NE(gen[8841]),

			.O(gen[8934]),
			.E(gen[8936]),

			.SO(gen[8839]),
			.S(gen[8840]),
			.SE(gen[8841]),

			.SELF(gen[8935]),
			.cell_state(gen[8935])
		); 

/******************* CELL 8936 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8936 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8840]),
			.N(gen[8841]),
			.NE(gen[8842]),

			.O(gen[8935]),
			.E(gen[8937]),

			.SO(gen[8840]),
			.S(gen[8841]),
			.SE(gen[8842]),

			.SELF(gen[8936]),
			.cell_state(gen[8936])
		); 

/******************* CELL 8937 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8937 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8841]),
			.N(gen[8842]),
			.NE(gen[8843]),

			.O(gen[8936]),
			.E(gen[8938]),

			.SO(gen[8841]),
			.S(gen[8842]),
			.SE(gen[8843]),

			.SELF(gen[8937]),
			.cell_state(gen[8937])
		); 

/******************* CELL 8938 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8938 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8842]),
			.N(gen[8843]),
			.NE(gen[8844]),

			.O(gen[8937]),
			.E(gen[8939]),

			.SO(gen[8842]),
			.S(gen[8843]),
			.SE(gen[8844]),

			.SELF(gen[8938]),
			.cell_state(gen[8938])
		); 

/******************* CELL 8939 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8939 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8843]),
			.N(gen[8844]),
			.NE(gen[8845]),

			.O(gen[8938]),
			.E(gen[8940]),

			.SO(gen[8843]),
			.S(gen[8844]),
			.SE(gen[8845]),

			.SELF(gen[8939]),
			.cell_state(gen[8939])
		); 

/******************* CELL 8940 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8940 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8844]),
			.N(gen[8845]),
			.NE(gen[8846]),

			.O(gen[8939]),
			.E(gen[8941]),

			.SO(gen[8844]),
			.S(gen[8845]),
			.SE(gen[8846]),

			.SELF(gen[8940]),
			.cell_state(gen[8940])
		); 

/******************* CELL 8941 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8941 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8845]),
			.N(gen[8846]),
			.NE(gen[8847]),

			.O(gen[8940]),
			.E(gen[8942]),

			.SO(gen[8845]),
			.S(gen[8846]),
			.SE(gen[8847]),

			.SELF(gen[8941]),
			.cell_state(gen[8941])
		); 

/******************* CELL 8942 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8942 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8846]),
			.N(gen[8847]),
			.NE(gen[8848]),

			.O(gen[8941]),
			.E(gen[8943]),

			.SO(gen[8846]),
			.S(gen[8847]),
			.SE(gen[8848]),

			.SELF(gen[8942]),
			.cell_state(gen[8942])
		); 

/******************* CELL 8943 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8943 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8847]),
			.N(gen[8848]),
			.NE(gen[8849]),

			.O(gen[8942]),
			.E(gen[8944]),

			.SO(gen[8847]),
			.S(gen[8848]),
			.SE(gen[8849]),

			.SELF(gen[8943]),
			.cell_state(gen[8943])
		); 

/******************* CELL 8944 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8944 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8848]),
			.N(gen[8849]),
			.NE(gen[8850]),

			.O(gen[8943]),
			.E(gen[8945]),

			.SO(gen[8848]),
			.S(gen[8849]),
			.SE(gen[8850]),

			.SELF(gen[8944]),
			.cell_state(gen[8944])
		); 

/******************* CELL 8945 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8945 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8849]),
			.N(gen[8850]),
			.NE(gen[8851]),

			.O(gen[8944]),
			.E(gen[8946]),

			.SO(gen[8849]),
			.S(gen[8850]),
			.SE(gen[8851]),

			.SELF(gen[8945]),
			.cell_state(gen[8945])
		); 

/******************* CELL 8946 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8946 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8850]),
			.N(gen[8851]),
			.NE(gen[8852]),

			.O(gen[8945]),
			.E(gen[8947]),

			.SO(gen[8850]),
			.S(gen[8851]),
			.SE(gen[8852]),

			.SELF(gen[8946]),
			.cell_state(gen[8946])
		); 

/******************* CELL 8947 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8947 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8851]),
			.N(gen[8852]),
			.NE(gen[8853]),

			.O(gen[8946]),
			.E(gen[8948]),

			.SO(gen[8851]),
			.S(gen[8852]),
			.SE(gen[8853]),

			.SELF(gen[8947]),
			.cell_state(gen[8947])
		); 

/******************* CELL 8948 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8948 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8852]),
			.N(gen[8853]),
			.NE(gen[8854]),

			.O(gen[8947]),
			.E(gen[8949]),

			.SO(gen[8852]),
			.S(gen[8853]),
			.SE(gen[8854]),

			.SELF(gen[8948]),
			.cell_state(gen[8948])
		); 

/******************* CELL 8949 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8949 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8853]),
			.N(gen[8854]),
			.NE(gen[8855]),

			.O(gen[8948]),
			.E(gen[8950]),

			.SO(gen[8853]),
			.S(gen[8854]),
			.SE(gen[8855]),

			.SELF(gen[8949]),
			.cell_state(gen[8949])
		); 

/******************* CELL 8950 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8950 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8854]),
			.N(gen[8855]),
			.NE(gen[8856]),

			.O(gen[8949]),
			.E(gen[8951]),

			.SO(gen[8854]),
			.S(gen[8855]),
			.SE(gen[8856]),

			.SELF(gen[8950]),
			.cell_state(gen[8950])
		); 

/******************* CELL 8951 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8951 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8855]),
			.N(gen[8856]),
			.NE(gen[8857]),

			.O(gen[8950]),
			.E(gen[8952]),

			.SO(gen[8855]),
			.S(gen[8856]),
			.SE(gen[8857]),

			.SELF(gen[8951]),
			.cell_state(gen[8951])
		); 

/******************* CELL 8952 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8952 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8856]),
			.N(gen[8857]),
			.NE(gen[8858]),

			.O(gen[8951]),
			.E(gen[8953]),

			.SO(gen[8856]),
			.S(gen[8857]),
			.SE(gen[8858]),

			.SELF(gen[8952]),
			.cell_state(gen[8952])
		); 

/******************* CELL 8953 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8953 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8857]),
			.N(gen[8858]),
			.NE(gen[8859]),

			.O(gen[8952]),
			.E(gen[8954]),

			.SO(gen[8857]),
			.S(gen[8858]),
			.SE(gen[8859]),

			.SELF(gen[8953]),
			.cell_state(gen[8953])
		); 

/******************* CELL 8954 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8954 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8858]),
			.N(gen[8859]),
			.NE(gen[8860]),

			.O(gen[8953]),
			.E(gen[8955]),

			.SO(gen[8858]),
			.S(gen[8859]),
			.SE(gen[8860]),

			.SELF(gen[8954]),
			.cell_state(gen[8954])
		); 

/******************* CELL 8955 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8955 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8859]),
			.N(gen[8860]),
			.NE(gen[8861]),

			.O(gen[8954]),
			.E(gen[8956]),

			.SO(gen[8859]),
			.S(gen[8860]),
			.SE(gen[8861]),

			.SELF(gen[8955]),
			.cell_state(gen[8955])
		); 

/******************* CELL 8956 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8956 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8860]),
			.N(gen[8861]),
			.NE(gen[8862]),

			.O(gen[8955]),
			.E(gen[8957]),

			.SO(gen[8860]),
			.S(gen[8861]),
			.SE(gen[8862]),

			.SELF(gen[8956]),
			.cell_state(gen[8956])
		); 

/******************* CELL 8957 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8957 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8861]),
			.N(gen[8862]),
			.NE(gen[8863]),

			.O(gen[8956]),
			.E(gen[8958]),

			.SO(gen[8861]),
			.S(gen[8862]),
			.SE(gen[8863]),

			.SELF(gen[8957]),
			.cell_state(gen[8957])
		); 

/******************* CELL 8958 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8958 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8862]),
			.N(gen[8863]),
			.NE(gen[8864]),

			.O(gen[8957]),
			.E(gen[8959]),

			.SO(gen[8862]),
			.S(gen[8863]),
			.SE(gen[8864]),

			.SELF(gen[8958]),
			.cell_state(gen[8958])
		); 

/******************* CELL 8959 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8959 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8863]),
			.N(gen[8864]),
			.NE(gen[8865]),

			.O(gen[8958]),
			.E(gen[8960]),

			.SO(gen[8863]),
			.S(gen[8864]),
			.SE(gen[8865]),

			.SELF(gen[8959]),
			.cell_state(gen[8959])
		); 

/******************* CELL 8960 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8960 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8864]),
			.N(gen[8865]),
			.NE(gen[8866]),

			.O(gen[8959]),
			.E(gen[8961]),

			.SO(gen[8864]),
			.S(gen[8865]),
			.SE(gen[8866]),

			.SELF(gen[8960]),
			.cell_state(gen[8960])
		); 

/******************* CELL 8961 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8961 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8865]),
			.N(gen[8866]),
			.NE(gen[8867]),

			.O(gen[8960]),
			.E(gen[8962]),

			.SO(gen[8865]),
			.S(gen[8866]),
			.SE(gen[8867]),

			.SELF(gen[8961]),
			.cell_state(gen[8961])
		); 

/******************* CELL 8962 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8962 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8866]),
			.N(gen[8867]),
			.NE(gen[8868]),

			.O(gen[8961]),
			.E(gen[8963]),

			.SO(gen[8866]),
			.S(gen[8867]),
			.SE(gen[8868]),

			.SELF(gen[8962]),
			.cell_state(gen[8962])
		); 

/******************* CELL 8963 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8963 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8867]),
			.N(gen[8868]),
			.NE(gen[8869]),

			.O(gen[8962]),
			.E(gen[8964]),

			.SO(gen[8867]),
			.S(gen[8868]),
			.SE(gen[8869]),

			.SELF(gen[8963]),
			.cell_state(gen[8963])
		); 

/******************* CELL 8964 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8964 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8868]),
			.N(gen[8869]),
			.NE(gen[8870]),

			.O(gen[8963]),
			.E(gen[8965]),

			.SO(gen[8868]),
			.S(gen[8869]),
			.SE(gen[8870]),

			.SELF(gen[8964]),
			.cell_state(gen[8964])
		); 

/******************* CELL 8965 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8965 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8869]),
			.N(gen[8870]),
			.NE(gen[8871]),

			.O(gen[8964]),
			.E(gen[8966]),

			.SO(gen[8869]),
			.S(gen[8870]),
			.SE(gen[8871]),

			.SELF(gen[8965]),
			.cell_state(gen[8965])
		); 

/******************* CELL 8966 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8966 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8870]),
			.N(gen[8871]),
			.NE(gen[8872]),

			.O(gen[8965]),
			.E(gen[8967]),

			.SO(gen[8870]),
			.S(gen[8871]),
			.SE(gen[8872]),

			.SELF(gen[8966]),
			.cell_state(gen[8966])
		); 

/******************* CELL 8967 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8967 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8871]),
			.N(gen[8872]),
			.NE(gen[8873]),

			.O(gen[8966]),
			.E(gen[8968]),

			.SO(gen[8871]),
			.S(gen[8872]),
			.SE(gen[8873]),

			.SELF(gen[8967]),
			.cell_state(gen[8967])
		); 

/******************* CELL 8968 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8968 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8872]),
			.N(gen[8873]),
			.NE(gen[8874]),

			.O(gen[8967]),
			.E(gen[8969]),

			.SO(gen[8872]),
			.S(gen[8873]),
			.SE(gen[8874]),

			.SELF(gen[8968]),
			.cell_state(gen[8968])
		); 

/******************* CELL 8969 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8969 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8873]),
			.N(gen[8874]),
			.NE(gen[8875]),

			.O(gen[8968]),
			.E(gen[8970]),

			.SO(gen[8873]),
			.S(gen[8874]),
			.SE(gen[8875]),

			.SELF(gen[8969]),
			.cell_state(gen[8969])
		); 

/******************* CELL 8970 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8970 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8874]),
			.N(gen[8875]),
			.NE(gen[8876]),

			.O(gen[8969]),
			.E(gen[8971]),

			.SO(gen[8874]),
			.S(gen[8875]),
			.SE(gen[8876]),

			.SELF(gen[8970]),
			.cell_state(gen[8970])
		); 

/******************* CELL 8971 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8971 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8875]),
			.N(gen[8876]),
			.NE(gen[8877]),

			.O(gen[8970]),
			.E(gen[8972]),

			.SO(gen[8875]),
			.S(gen[8876]),
			.SE(gen[8877]),

			.SELF(gen[8971]),
			.cell_state(gen[8971])
		); 

/******************* CELL 8972 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8972 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8876]),
			.N(gen[8877]),
			.NE(gen[8878]),

			.O(gen[8971]),
			.E(gen[8973]),

			.SO(gen[8876]),
			.S(gen[8877]),
			.SE(gen[8878]),

			.SELF(gen[8972]),
			.cell_state(gen[8972])
		); 

/******************* CELL 8973 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8973 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8877]),
			.N(gen[8878]),
			.NE(gen[8879]),

			.O(gen[8972]),
			.E(gen[8974]),

			.SO(gen[8877]),
			.S(gen[8878]),
			.SE(gen[8879]),

			.SELF(gen[8973]),
			.cell_state(gen[8973])
		); 

/******************* CELL 8974 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8974 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8878]),
			.N(gen[8879]),
			.NE(gen[8880]),

			.O(gen[8973]),
			.E(gen[8975]),

			.SO(gen[8878]),
			.S(gen[8879]),
			.SE(gen[8880]),

			.SELF(gen[8974]),
			.cell_state(gen[8974])
		); 

/******************* CELL 8975 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8975 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8879]),
			.N(gen[8880]),
			.NE(gen[8881]),

			.O(gen[8974]),
			.E(gen[8976]),

			.SO(gen[8879]),
			.S(gen[8880]),
			.SE(gen[8881]),

			.SELF(gen[8975]),
			.cell_state(gen[8975])
		); 

/******************* CELL 8976 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8976 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8880]),
			.N(gen[8881]),
			.NE(gen[8882]),

			.O(gen[8975]),
			.E(gen[8977]),

			.SO(gen[8880]),
			.S(gen[8881]),
			.SE(gen[8882]),

			.SELF(gen[8976]),
			.cell_state(gen[8976])
		); 

/******************* CELL 8977 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8977 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8881]),
			.N(gen[8882]),
			.NE(gen[8883]),

			.O(gen[8976]),
			.E(gen[8978]),

			.SO(gen[8881]),
			.S(gen[8882]),
			.SE(gen[8883]),

			.SELF(gen[8977]),
			.cell_state(gen[8977])
		); 

/******************* CELL 8978 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8978 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8882]),
			.N(gen[8883]),
			.NE(gen[8884]),

			.O(gen[8977]),
			.E(gen[8979]),

			.SO(gen[8882]),
			.S(gen[8883]),
			.SE(gen[8884]),

			.SELF(gen[8978]),
			.cell_state(gen[8978])
		); 

/******************* CELL 8979 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8979 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8883]),
			.N(gen[8884]),
			.NE(gen[8885]),

			.O(gen[8978]),
			.E(gen[8980]),

			.SO(gen[8883]),
			.S(gen[8884]),
			.SE(gen[8885]),

			.SELF(gen[8979]),
			.cell_state(gen[8979])
		); 

/******************* CELL 8980 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8980 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8884]),
			.N(gen[8885]),
			.NE(gen[8886]),

			.O(gen[8979]),
			.E(gen[8981]),

			.SO(gen[8884]),
			.S(gen[8885]),
			.SE(gen[8886]),

			.SELF(gen[8980]),
			.cell_state(gen[8980])
		); 

/******************* CELL 8981 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8981 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8885]),
			.N(gen[8886]),
			.NE(gen[8887]),

			.O(gen[8980]),
			.E(gen[8982]),

			.SO(gen[8885]),
			.S(gen[8886]),
			.SE(gen[8887]),

			.SELF(gen[8981]),
			.cell_state(gen[8981])
		); 

/******************* CELL 8982 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8982 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8886]),
			.N(gen[8887]),
			.NE(gen[8888]),

			.O(gen[8981]),
			.E(gen[8983]),

			.SO(gen[8886]),
			.S(gen[8887]),
			.SE(gen[8888]),

			.SELF(gen[8982]),
			.cell_state(gen[8982])
		); 

/******************* CELL 8983 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8983 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8887]),
			.N(gen[8888]),
			.NE(gen[8889]),

			.O(gen[8982]),
			.E(gen[8984]),

			.SO(gen[8887]),
			.S(gen[8888]),
			.SE(gen[8889]),

			.SELF(gen[8983]),
			.cell_state(gen[8983])
		); 

/******************* CELL 8984 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8984 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8888]),
			.N(gen[8889]),
			.NE(gen[8890]),

			.O(gen[8983]),
			.E(gen[8985]),

			.SO(gen[8888]),
			.S(gen[8889]),
			.SE(gen[8890]),

			.SELF(gen[8984]),
			.cell_state(gen[8984])
		); 

/******************* CELL 8985 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8985 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8889]),
			.N(gen[8890]),
			.NE(gen[8891]),

			.O(gen[8984]),
			.E(gen[8986]),

			.SO(gen[8889]),
			.S(gen[8890]),
			.SE(gen[8891]),

			.SELF(gen[8985]),
			.cell_state(gen[8985])
		); 

/******************* CELL 8986 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8986 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8890]),
			.N(gen[8891]),
			.NE(gen[8892]),

			.O(gen[8985]),
			.E(gen[8987]),

			.SO(gen[8890]),
			.S(gen[8891]),
			.SE(gen[8892]),

			.SELF(gen[8986]),
			.cell_state(gen[8986])
		); 

/******************* CELL 8987 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8987 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8891]),
			.N(gen[8892]),
			.NE(gen[8893]),

			.O(gen[8986]),
			.E(gen[8988]),

			.SO(gen[8891]),
			.S(gen[8892]),
			.SE(gen[8893]),

			.SELF(gen[8987]),
			.cell_state(gen[8987])
		); 

/******************* CELL 8988 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8988 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8892]),
			.N(gen[8893]),
			.NE(gen[8894]),

			.O(gen[8987]),
			.E(gen[8989]),

			.SO(gen[8892]),
			.S(gen[8893]),
			.SE(gen[8894]),

			.SELF(gen[8988]),
			.cell_state(gen[8988])
		); 

/******************* CELL 8989 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8989 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8893]),
			.N(gen[8894]),
			.NE(gen[8895]),

			.O(gen[8988]),
			.E(gen[8990]),

			.SO(gen[8893]),
			.S(gen[8894]),
			.SE(gen[8895]),

			.SELF(gen[8989]),
			.cell_state(gen[8989])
		); 

/******************* CELL 8990 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8990 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8894]),
			.N(gen[8895]),
			.NE(gen[8896]),

			.O(gen[8989]),
			.E(gen[8991]),

			.SO(gen[8894]),
			.S(gen[8895]),
			.SE(gen[8896]),

			.SELF(gen[8990]),
			.cell_state(gen[8990])
		); 

/******************* CELL 8991 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8991 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8895]),
			.N(gen[8896]),
			.NE(gen[8897]),

			.O(gen[8990]),
			.E(gen[8992]),

			.SO(gen[8895]),
			.S(gen[8896]),
			.SE(gen[8897]),

			.SELF(gen[8991]),
			.cell_state(gen[8991])
		); 

/******************* CELL 8992 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8992 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8896]),
			.N(gen[8897]),
			.NE(gen[8898]),

			.O(gen[8991]),
			.E(gen[8993]),

			.SO(gen[8896]),
			.S(gen[8897]),
			.SE(gen[8898]),

			.SELF(gen[8992]),
			.cell_state(gen[8992])
		); 

/******************* CELL 8993 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8993 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8897]),
			.N(gen[8898]),
			.NE(gen[8899]),

			.O(gen[8992]),
			.E(gen[8994]),

			.SO(gen[8897]),
			.S(gen[8898]),
			.SE(gen[8899]),

			.SELF(gen[8993]),
			.cell_state(gen[8993])
		); 

/******************* CELL 8994 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8994 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8898]),
			.N(gen[8899]),
			.NE(gen[8900]),

			.O(gen[8993]),
			.E(gen[8995]),

			.SO(gen[8898]),
			.S(gen[8899]),
			.SE(gen[8900]),

			.SELF(gen[8994]),
			.cell_state(gen[8994])
		); 

/******************* CELL 8995 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8995 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8899]),
			.N(gen[8900]),
			.NE(gen[8901]),

			.O(gen[8994]),
			.E(gen[8996]),

			.SO(gen[8899]),
			.S(gen[8900]),
			.SE(gen[8901]),

			.SELF(gen[8995]),
			.cell_state(gen[8995])
		); 

/******************* CELL 8996 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8996 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8900]),
			.N(gen[8901]),
			.NE(gen[8902]),

			.O(gen[8995]),
			.E(gen[8997]),

			.SO(gen[8900]),
			.S(gen[8901]),
			.SE(gen[8902]),

			.SELF(gen[8996]),
			.cell_state(gen[8996])
		); 

/******************* CELL 8997 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8997 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8901]),
			.N(gen[8902]),
			.NE(gen[8903]),

			.O(gen[8996]),
			.E(gen[8998]),

			.SO(gen[8901]),
			.S(gen[8902]),
			.SE(gen[8903]),

			.SELF(gen[8997]),
			.cell_state(gen[8997])
		); 

/******************* CELL 8998 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8998 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8902]),
			.N(gen[8903]),
			.NE(gen[8904]),

			.O(gen[8997]),
			.E(gen[8999]),

			.SO(gen[8902]),
			.S(gen[8903]),
			.SE(gen[8904]),

			.SELF(gen[8998]),
			.cell_state(gen[8998])
		); 

/******************* CELL 8999 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell8999 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8903]),
			.N(gen[8904]),
			.NE(gen[8905]),

			.O(gen[8998]),
			.E(gen[9000]),

			.SO(gen[8903]),
			.S(gen[8904]),
			.SE(gen[8905]),

			.SELF(gen[8999]),
			.cell_state(gen[8999])
		); 

/******************* CELL 9000 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell9000 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8904]),
			.N(gen[8905]),
			.NE(gen[8906]),

			.O(gen[8999]),
			.E(gen[9001]),

			.SO(gen[8904]),
			.S(gen[8905]),
			.SE(gen[8906]),

			.SELF(gen[9000]),
			.cell_state(gen[9000])
		); 

/******************* CELL 9001 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell9001 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8905]),
			.N(gen[8906]),
			.NE(gen[8907]),

			.O(gen[9000]),
			.E(gen[9002]),

			.SO(gen[8905]),
			.S(gen[8906]),
			.SE(gen[8907]),

			.SELF(gen[9001]),
			.cell_state(gen[9001])
		); 

/******************* CELL 9002 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell9002 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8906]),
			.N(gen[8907]),
			.NE(gen[8908]),

			.O(gen[9001]),
			.E(gen[9003]),

			.SO(gen[8906]),
			.S(gen[8907]),
			.SE(gen[8908]),

			.SELF(gen[9002]),
			.cell_state(gen[9002])
		); 

/******************* CELL 9003 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell9003 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8907]),
			.N(gen[8908]),
			.NE(gen[8909]),

			.O(gen[9002]),
			.E(gen[9004]),

			.SO(gen[8907]),
			.S(gen[8908]),
			.SE(gen[8909]),

			.SELF(gen[9003]),
			.cell_state(gen[9003])
		); 

/******************* CELL 9004 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell9004 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8908]),
			.N(gen[8909]),
			.NE(gen[8910]),

			.O(gen[9003]),
			.E(gen[9005]),

			.SO(gen[8908]),
			.S(gen[8909]),
			.SE(gen[8910]),

			.SELF(gen[9004]),
			.cell_state(gen[9004])
		); 

/******************* CELL 9005 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell9005 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8909]),
			.N(gen[8910]),
			.NE(gen[8911]),

			.O(gen[9004]),
			.E(gen[9006]),

			.SO(gen[8909]),
			.S(gen[8910]),
			.SE(gen[8911]),

			.SELF(gen[9005]),
			.cell_state(gen[9005])
		); 

/******************* CELL 9006 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell9006 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8910]),
			.N(gen[8911]),
			.NE(gen[8912]),

			.O(gen[9005]),
			.E(gen[9007]),

			.SO(gen[8910]),
			.S(gen[8911]),
			.SE(gen[8912]),

			.SELF(gen[9006]),
			.cell_state(gen[9006])
		); 

/******************* CELL 9007 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell9007 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8911]),
			.N(gen[8912]),
			.NE(gen[8913]),

			.O(gen[9006]),
			.E(gen[9008]),

			.SO(gen[8911]),
			.S(gen[8912]),
			.SE(gen[8913]),

			.SELF(gen[9007]),
			.cell_state(gen[9007])
		); 

/******************* CELL 9008 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell9008 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8912]),
			.N(gen[8913]),
			.NE(gen[8914]),

			.O(gen[9007]),
			.E(gen[9009]),

			.SO(gen[8912]),
			.S(gen[8913]),
			.SE(gen[8914]),

			.SELF(gen[9008]),
			.cell_state(gen[9008])
		); 

/******************* CELL 9009 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell9009 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8913]),
			.N(gen[8914]),
			.NE(gen[8915]),

			.O(gen[9008]),
			.E(gen[9010]),

			.SO(gen[8913]),
			.S(gen[8914]),
			.SE(gen[8915]),

			.SELF(gen[9009]),
			.cell_state(gen[9009])
		); 

/******************* CELL 9010 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell9010 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8914]),
			.N(gen[8915]),
			.NE(gen[8916]),

			.O(gen[9009]),
			.E(gen[9011]),

			.SO(gen[8914]),
			.S(gen[8915]),
			.SE(gen[8916]),

			.SELF(gen[9010]),
			.cell_state(gen[9010])
		); 

/******************* CELL 9011 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell9011 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8915]),
			.N(gen[8916]),
			.NE(gen[8917]),

			.O(gen[9010]),
			.E(gen[9012]),

			.SO(gen[8915]),
			.S(gen[8916]),
			.SE(gen[8917]),

			.SELF(gen[9011]),
			.cell_state(gen[9011])
		); 

/******************* CELL 9012 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell9012 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8916]),
			.N(gen[8917]),
			.NE(gen[8918]),

			.O(gen[9011]),
			.E(gen[9013]),

			.SO(gen[8916]),
			.S(gen[8917]),
			.SE(gen[8918]),

			.SELF(gen[9012]),
			.cell_state(gen[9012])
		); 

/******************* CELL 9013 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell9013 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8917]),
			.N(gen[8918]),
			.NE(gen[8919]),

			.O(gen[9012]),
			.E(gen[9014]),

			.SO(gen[8917]),
			.S(gen[8918]),
			.SE(gen[8919]),

			.SELF(gen[9013]),
			.cell_state(gen[9013])
		); 

/******************* CELL 9014 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell9014 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8918]),
			.N(gen[8919]),
			.NE(gen[8920]),

			.O(gen[9013]),
			.E(gen[9015]),

			.SO(gen[8918]),
			.S(gen[8919]),
			.SE(gen[8920]),

			.SELF(gen[9014]),
			.cell_state(gen[9014])
		); 

/******************* CELL 9015 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell9015 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8919]),
			.N(gen[8920]),
			.NE(gen[8921]),

			.O(gen[9014]),
			.E(gen[9016]),

			.SO(gen[8919]),
			.S(gen[8920]),
			.SE(gen[8921]),

			.SELF(gen[9015]),
			.cell_state(gen[9015])
		); 

/******************* CELL 9016 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell9016 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8920]),
			.N(gen[8921]),
			.NE(gen[8922]),

			.O(gen[9015]),
			.E(gen[9017]),

			.SO(gen[8920]),
			.S(gen[8921]),
			.SE(gen[8922]),

			.SELF(gen[9016]),
			.cell_state(gen[9016])
		); 

/******************* CELL 9017 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell9017 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8921]),
			.N(gen[8922]),
			.NE(gen[8923]),

			.O(gen[9016]),
			.E(gen[9018]),

			.SO(gen[8921]),
			.S(gen[8922]),
			.SE(gen[8923]),

			.SELF(gen[9017]),
			.cell_state(gen[9017])
		); 

/******************* CELL 9018 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell9018 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8922]),
			.N(gen[8923]),
			.NE(gen[8924]),

			.O(gen[9017]),
			.E(gen[9019]),

			.SO(gen[8922]),
			.S(gen[8923]),
			.SE(gen[8924]),

			.SELF(gen[9018]),
			.cell_state(gen[9018])
		); 

/******************* CELL 9019 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell9019 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8923]),
			.N(gen[8924]),
			.NE(gen[8925]),

			.O(gen[9018]),
			.E(gen[9020]),

			.SO(gen[8923]),
			.S(gen[8924]),
			.SE(gen[8925]),

			.SELF(gen[9019]),
			.cell_state(gen[9019])
		); 

/******************* CELL 9020 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell9020 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8924]),
			.N(gen[8925]),
			.NE(gen[8926]),

			.O(gen[9019]),
			.E(gen[9021]),

			.SO(gen[8924]),
			.S(gen[8925]),
			.SE(gen[8926]),

			.SELF(gen[9020]),
			.cell_state(gen[9020])
		); 

/******************* CELL 9021 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell9021 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8925]),
			.N(gen[8926]),
			.NE(gen[8927]),

			.O(gen[9020]),
			.E(gen[9022]),

			.SO(gen[8925]),
			.S(gen[8926]),
			.SE(gen[8927]),

			.SELF(gen[9021]),
			.cell_state(gen[9021])
		); 

/******************* CELL 9022 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell9022 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8926]),
			.N(gen[8927]),
			.NE(gen[8928]),

			.O(gen[9021]),
			.E(gen[9023]),

			.SO(gen[8926]),
			.S(gen[8927]),
			.SE(gen[8928]),

			.SELF(gen[9022]),
			.cell_state(gen[9022])
		); 

/******************* CELL 9023 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell9023 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8927]),
			.N(gen[8928]),
			.NE(gen[8929]),

			.O(gen[9022]),
			.E(gen[9024]),

			.SO(gen[8927]),
			.S(gen[8928]),
			.SE(gen[8929]),

			.SELF(gen[9023]),
			.cell_state(gen[9023])
		); 

/******************* CELL 9024 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell9024 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8928]),
			.N(gen[8929]),
			.NE(gen[8928]),

			.O(gen[9023]),
			.E(gen[9023]),

			.SO(gen[8928]),
			.S(gen[8929]),
			.SE(gen[8928]),

			.SELF(gen[9024]),
			.cell_state(gen[9024])
		); 



 assign data_out = {7'b0, gen[9024]};

endmodule
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/10/2022 12:12:04 PM
// Design Name: 
// Module Name: GRID_SCRIPT
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module GRID_SCRIPT
    #(parameter M = 3, N = 3)

    (


    input logic clk, reset,
    
    input logic [2:0] operation,       
    
    input logic [0:0] data_in,
    
    
    
    output logic [0:0] gen [M*N -1 :0] ,
    output logic [7:0] data_out    
        
    );/******************* CELL 0 ***************/  

	CELDA   #(.ic(0), .top_row(1), .load_cell(1))

		cell0 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[61]),
			.N(gen[60]),
			.NE(gen[61]),

			.O(data_in),
			.E(gen[1]),

			.SO(gen[61]),
			.S(gen[60]),
			.SE(gen[61]),

			.SELF(gen[0]),
			.cell_state(gen[0])
		); 

/******************* CELL 1 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell1 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[60]),
			.N(gen[61]),
			.NE(gen[62]),

			.O(gen[0]),
			.E(gen[2]),

			.SO(gen[60]),
			.S(gen[61]),
			.SE(gen[62]),

			.SELF(gen[1]),
			.cell_state(gen[1])
		); 

/******************* CELL 2 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell2 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[61]),
			.N(gen[62]),
			.NE(gen[63]),

			.O(gen[1]),
			.E(gen[3]),

			.SO(gen[61]),
			.S(gen[62]),
			.SE(gen[63]),

			.SELF(gen[2]),
			.cell_state(gen[2])
		); 

/******************* CELL 3 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell3 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[62]),
			.N(gen[63]),
			.NE(gen[64]),

			.O(gen[2]),
			.E(gen[4]),

			.SO(gen[62]),
			.S(gen[63]),
			.SE(gen[64]),

			.SELF(gen[3]),
			.cell_state(gen[3])
		); 

/******************* CELL 4 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell4 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[63]),
			.N(gen[64]),
			.NE(gen[65]),

			.O(gen[3]),
			.E(gen[5]),

			.SO(gen[63]),
			.S(gen[64]),
			.SE(gen[65]),

			.SELF(gen[4]),
			.cell_state(gen[4])
		); 

/******************* CELL 5 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell5 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[64]),
			.N(gen[65]),
			.NE(gen[66]),

			.O(gen[4]),
			.E(gen[6]),

			.SO(gen[64]),
			.S(gen[65]),
			.SE(gen[66]),

			.SELF(gen[5]),
			.cell_state(gen[5])
		); 

/******************* CELL 6 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell6 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[65]),
			.N(gen[66]),
			.NE(gen[67]),

			.O(gen[5]),
			.E(gen[7]),

			.SO(gen[65]),
			.S(gen[66]),
			.SE(gen[67]),

			.SELF(gen[6]),
			.cell_state(gen[6])
		); 

/******************* CELL 7 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell7 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[66]),
			.N(gen[67]),
			.NE(gen[68]),

			.O(gen[6]),
			.E(gen[8]),

			.SO(gen[66]),
			.S(gen[67]),
			.SE(gen[68]),

			.SELF(gen[7]),
			.cell_state(gen[7])
		); 

/******************* CELL 8 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell8 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[67]),
			.N(gen[68]),
			.NE(gen[69]),

			.O(gen[7]),
			.E(gen[9]),

			.SO(gen[67]),
			.S(gen[68]),
			.SE(gen[69]),

			.SELF(gen[8]),
			.cell_state(gen[8])
		); 

/******************* CELL 9 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell9 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[68]),
			.N(gen[69]),
			.NE(gen[70]),

			.O(gen[8]),
			.E(gen[10]),

			.SO(gen[68]),
			.S(gen[69]),
			.SE(gen[70]),

			.SELF(gen[9]),
			.cell_state(gen[9])
		); 

/******************* CELL 10 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell10 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[69]),
			.N(gen[70]),
			.NE(gen[71]),

			.O(gen[9]),
			.E(gen[11]),

			.SO(gen[69]),
			.S(gen[70]),
			.SE(gen[71]),

			.SELF(gen[10]),
			.cell_state(gen[10])
		); 

/******************* CELL 11 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell11 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[70]),
			.N(gen[71]),
			.NE(gen[72]),

			.O(gen[10]),
			.E(gen[12]),

			.SO(gen[70]),
			.S(gen[71]),
			.SE(gen[72]),

			.SELF(gen[11]),
			.cell_state(gen[11])
		); 

/******************* CELL 12 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell12 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[71]),
			.N(gen[72]),
			.NE(gen[73]),

			.O(gen[11]),
			.E(gen[13]),

			.SO(gen[71]),
			.S(gen[72]),
			.SE(gen[73]),

			.SELF(gen[12]),
			.cell_state(gen[12])
		); 

/******************* CELL 13 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell13 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[72]),
			.N(gen[73]),
			.NE(gen[74]),

			.O(gen[12]),
			.E(gen[14]),

			.SO(gen[72]),
			.S(gen[73]),
			.SE(gen[74]),

			.SELF(gen[13]),
			.cell_state(gen[13])
		); 

/******************* CELL 14 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell14 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[73]),
			.N(gen[74]),
			.NE(gen[75]),

			.O(gen[13]),
			.E(gen[15]),

			.SO(gen[73]),
			.S(gen[74]),
			.SE(gen[75]),

			.SELF(gen[14]),
			.cell_state(gen[14])
		); 

/******************* CELL 15 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell15 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[74]),
			.N(gen[75]),
			.NE(gen[76]),

			.O(gen[14]),
			.E(gen[16]),

			.SO(gen[74]),
			.S(gen[75]),
			.SE(gen[76]),

			.SELF(gen[15]),
			.cell_state(gen[15])
		); 

/******************* CELL 16 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell16 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[75]),
			.N(gen[76]),
			.NE(gen[77]),

			.O(gen[15]),
			.E(gen[17]),

			.SO(gen[75]),
			.S(gen[76]),
			.SE(gen[77]),

			.SELF(gen[16]),
			.cell_state(gen[16])
		); 

/******************* CELL 17 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell17 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[76]),
			.N(gen[77]),
			.NE(gen[78]),

			.O(gen[16]),
			.E(gen[18]),

			.SO(gen[76]),
			.S(gen[77]),
			.SE(gen[78]),

			.SELF(gen[17]),
			.cell_state(gen[17])
		); 

/******************* CELL 18 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell18 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[77]),
			.N(gen[78]),
			.NE(gen[79]),

			.O(gen[17]),
			.E(gen[19]),

			.SO(gen[77]),
			.S(gen[78]),
			.SE(gen[79]),

			.SELF(gen[18]),
			.cell_state(gen[18])
		); 

/******************* CELL 19 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell19 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[78]),
			.N(gen[79]),
			.NE(gen[80]),

			.O(gen[18]),
			.E(gen[20]),

			.SO(gen[78]),
			.S(gen[79]),
			.SE(gen[80]),

			.SELF(gen[19]),
			.cell_state(gen[19])
		); 

/******************* CELL 20 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell20 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[79]),
			.N(gen[80]),
			.NE(gen[81]),

			.O(gen[19]),
			.E(gen[21]),

			.SO(gen[79]),
			.S(gen[80]),
			.SE(gen[81]),

			.SELF(gen[20]),
			.cell_state(gen[20])
		); 

/******************* CELL 21 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell21 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[80]),
			.N(gen[81]),
			.NE(gen[82]),

			.O(gen[20]),
			.E(gen[22]),

			.SO(gen[80]),
			.S(gen[81]),
			.SE(gen[82]),

			.SELF(gen[21]),
			.cell_state(gen[21])
		); 

/******************* CELL 22 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell22 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[81]),
			.N(gen[82]),
			.NE(gen[83]),

			.O(gen[21]),
			.E(gen[23]),

			.SO(gen[81]),
			.S(gen[82]),
			.SE(gen[83]),

			.SELF(gen[22]),
			.cell_state(gen[22])
		); 

/******************* CELL 23 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell23 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[82]),
			.N(gen[83]),
			.NE(gen[84]),

			.O(gen[22]),
			.E(gen[24]),

			.SO(gen[82]),
			.S(gen[83]),
			.SE(gen[84]),

			.SELF(gen[23]),
			.cell_state(gen[23])
		); 

/******************* CELL 24 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell24 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[83]),
			.N(gen[84]),
			.NE(gen[85]),

			.O(gen[23]),
			.E(gen[25]),

			.SO(gen[83]),
			.S(gen[84]),
			.SE(gen[85]),

			.SELF(gen[24]),
			.cell_state(gen[24])
		); 

/******************* CELL 25 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell25 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[84]),
			.N(gen[85]),
			.NE(gen[86]),

			.O(gen[24]),
			.E(gen[26]),

			.SO(gen[84]),
			.S(gen[85]),
			.SE(gen[86]),

			.SELF(gen[25]),
			.cell_state(gen[25])
		); 

/******************* CELL 26 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell26 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[85]),
			.N(gen[86]),
			.NE(gen[87]),

			.O(gen[25]),
			.E(gen[27]),

			.SO(gen[85]),
			.S(gen[86]),
			.SE(gen[87]),

			.SELF(gen[26]),
			.cell_state(gen[26])
		); 

/******************* CELL 27 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell27 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[86]),
			.N(gen[87]),
			.NE(gen[88]),

			.O(gen[26]),
			.E(gen[28]),

			.SO(gen[86]),
			.S(gen[87]),
			.SE(gen[88]),

			.SELF(gen[27]),
			.cell_state(gen[27])
		); 

/******************* CELL 28 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell28 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[87]),
			.N(gen[88]),
			.NE(gen[89]),

			.O(gen[27]),
			.E(gen[29]),

			.SO(gen[87]),
			.S(gen[88]),
			.SE(gen[89]),

			.SELF(gen[28]),
			.cell_state(gen[28])
		); 

/******************* CELL 29 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell29 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[88]),
			.N(gen[89]),
			.NE(gen[90]),

			.O(gen[28]),
			.E(gen[30]),

			.SO(gen[88]),
			.S(gen[89]),
			.SE(gen[90]),

			.SELF(gen[29]),
			.cell_state(gen[29])
		); 

/******************* CELL 30 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell30 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[89]),
			.N(gen[90]),
			.NE(gen[91]),

			.O(gen[29]),
			.E(gen[31]),

			.SO(gen[89]),
			.S(gen[90]),
			.SE(gen[91]),

			.SELF(gen[30]),
			.cell_state(gen[30])
		); 

/******************* CELL 31 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell31 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[90]),
			.N(gen[91]),
			.NE(gen[92]),

			.O(gen[30]),
			.E(gen[32]),

			.SO(gen[90]),
			.S(gen[91]),
			.SE(gen[92]),

			.SELF(gen[31]),
			.cell_state(gen[31])
		); 

/******************* CELL 32 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell32 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[91]),
			.N(gen[92]),
			.NE(gen[93]),

			.O(gen[31]),
			.E(gen[33]),

			.SO(gen[91]),
			.S(gen[92]),
			.SE(gen[93]),

			.SELF(gen[32]),
			.cell_state(gen[32])
		); 

/******************* CELL 33 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell33 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[92]),
			.N(gen[93]),
			.NE(gen[94]),

			.O(gen[32]),
			.E(gen[34]),

			.SO(gen[92]),
			.S(gen[93]),
			.SE(gen[94]),

			.SELF(gen[33]),
			.cell_state(gen[33])
		); 

/******************* CELL 34 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell34 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[93]),
			.N(gen[94]),
			.NE(gen[95]),

			.O(gen[33]),
			.E(gen[35]),

			.SO(gen[93]),
			.S(gen[94]),
			.SE(gen[95]),

			.SELF(gen[34]),
			.cell_state(gen[34])
		); 

/******************* CELL 35 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell35 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[94]),
			.N(gen[95]),
			.NE(gen[96]),

			.O(gen[34]),
			.E(gen[36]),

			.SO(gen[94]),
			.S(gen[95]),
			.SE(gen[96]),

			.SELF(gen[35]),
			.cell_state(gen[35])
		); 

/******************* CELL 36 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell36 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[95]),
			.N(gen[96]),
			.NE(gen[97]),

			.O(gen[35]),
			.E(gen[37]),

			.SO(gen[95]),
			.S(gen[96]),
			.SE(gen[97]),

			.SELF(gen[36]),
			.cell_state(gen[36])
		); 

/******************* CELL 37 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell37 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[96]),
			.N(gen[97]),
			.NE(gen[98]),

			.O(gen[36]),
			.E(gen[38]),

			.SO(gen[96]),
			.S(gen[97]),
			.SE(gen[98]),

			.SELF(gen[37]),
			.cell_state(gen[37])
		); 

/******************* CELL 38 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell38 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[97]),
			.N(gen[98]),
			.NE(gen[99]),

			.O(gen[37]),
			.E(gen[39]),

			.SO(gen[97]),
			.S(gen[98]),
			.SE(gen[99]),

			.SELF(gen[38]),
			.cell_state(gen[38])
		); 

/******************* CELL 39 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell39 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[98]),
			.N(gen[99]),
			.NE(gen[100]),

			.O(gen[38]),
			.E(gen[40]),

			.SO(gen[98]),
			.S(gen[99]),
			.SE(gen[100]),

			.SELF(gen[39]),
			.cell_state(gen[39])
		); 

/******************* CELL 40 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell40 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[99]),
			.N(gen[100]),
			.NE(gen[101]),

			.O(gen[39]),
			.E(gen[41]),

			.SO(gen[99]),
			.S(gen[100]),
			.SE(gen[101]),

			.SELF(gen[40]),
			.cell_state(gen[40])
		); 

/******************* CELL 41 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell41 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[100]),
			.N(gen[101]),
			.NE(gen[102]),

			.O(gen[40]),
			.E(gen[42]),

			.SO(gen[100]),
			.S(gen[101]),
			.SE(gen[102]),

			.SELF(gen[41]),
			.cell_state(gen[41])
		); 

/******************* CELL 42 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell42 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[101]),
			.N(gen[102]),
			.NE(gen[103]),

			.O(gen[41]),
			.E(gen[43]),

			.SO(gen[101]),
			.S(gen[102]),
			.SE(gen[103]),

			.SELF(gen[42]),
			.cell_state(gen[42])
		); 

/******************* CELL 43 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell43 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[102]),
			.N(gen[103]),
			.NE(gen[104]),

			.O(gen[42]),
			.E(gen[44]),

			.SO(gen[102]),
			.S(gen[103]),
			.SE(gen[104]),

			.SELF(gen[43]),
			.cell_state(gen[43])
		); 

/******************* CELL 44 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell44 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[103]),
			.N(gen[104]),
			.NE(gen[105]),

			.O(gen[43]),
			.E(gen[45]),

			.SO(gen[103]),
			.S(gen[104]),
			.SE(gen[105]),

			.SELF(gen[44]),
			.cell_state(gen[44])
		); 

/******************* CELL 45 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell45 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[104]),
			.N(gen[105]),
			.NE(gen[106]),

			.O(gen[44]),
			.E(gen[46]),

			.SO(gen[104]),
			.S(gen[105]),
			.SE(gen[106]),

			.SELF(gen[45]),
			.cell_state(gen[45])
		); 

/******************* CELL 46 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell46 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[105]),
			.N(gen[106]),
			.NE(gen[107]),

			.O(gen[45]),
			.E(gen[47]),

			.SO(gen[105]),
			.S(gen[106]),
			.SE(gen[107]),

			.SELF(gen[46]),
			.cell_state(gen[46])
		); 

/******************* CELL 47 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell47 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[106]),
			.N(gen[107]),
			.NE(gen[108]),

			.O(gen[46]),
			.E(gen[48]),

			.SO(gen[106]),
			.S(gen[107]),
			.SE(gen[108]),

			.SELF(gen[47]),
			.cell_state(gen[47])
		); 

/******************* CELL 48 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell48 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[107]),
			.N(gen[108]),
			.NE(gen[109]),

			.O(gen[47]),
			.E(gen[49]),

			.SO(gen[107]),
			.S(gen[108]),
			.SE(gen[109]),

			.SELF(gen[48]),
			.cell_state(gen[48])
		); 

/******************* CELL 49 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell49 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[108]),
			.N(gen[109]),
			.NE(gen[110]),

			.O(gen[48]),
			.E(gen[50]),

			.SO(gen[108]),
			.S(gen[109]),
			.SE(gen[110]),

			.SELF(gen[49]),
			.cell_state(gen[49])
		); 

/******************* CELL 50 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell50 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[109]),
			.N(gen[110]),
			.NE(gen[111]),

			.O(gen[49]),
			.E(gen[51]),

			.SO(gen[109]),
			.S(gen[110]),
			.SE(gen[111]),

			.SELF(gen[50]),
			.cell_state(gen[50])
		); 

/******************* CELL 51 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell51 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[110]),
			.N(gen[111]),
			.NE(gen[112]),

			.O(gen[50]),
			.E(gen[52]),

			.SO(gen[110]),
			.S(gen[111]),
			.SE(gen[112]),

			.SELF(gen[51]),
			.cell_state(gen[51])
		); 

/******************* CELL 52 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell52 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[111]),
			.N(gen[112]),
			.NE(gen[113]),

			.O(gen[51]),
			.E(gen[53]),

			.SO(gen[111]),
			.S(gen[112]),
			.SE(gen[113]),

			.SELF(gen[52]),
			.cell_state(gen[52])
		); 

/******************* CELL 53 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell53 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[112]),
			.N(gen[113]),
			.NE(gen[114]),

			.O(gen[52]),
			.E(gen[54]),

			.SO(gen[112]),
			.S(gen[113]),
			.SE(gen[114]),

			.SELF(gen[53]),
			.cell_state(gen[53])
		); 

/******************* CELL 54 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell54 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[113]),
			.N(gen[114]),
			.NE(gen[115]),

			.O(gen[53]),
			.E(gen[55]),

			.SO(gen[113]),
			.S(gen[114]),
			.SE(gen[115]),

			.SELF(gen[54]),
			.cell_state(gen[54])
		); 

/******************* CELL 55 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell55 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[114]),
			.N(gen[115]),
			.NE(gen[116]),

			.O(gen[54]),
			.E(gen[56]),

			.SO(gen[114]),
			.S(gen[115]),
			.SE(gen[116]),

			.SELF(gen[55]),
			.cell_state(gen[55])
		); 

/******************* CELL 56 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell56 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[115]),
			.N(gen[116]),
			.NE(gen[117]),

			.O(gen[55]),
			.E(gen[57]),

			.SO(gen[115]),
			.S(gen[116]),
			.SE(gen[117]),

			.SELF(gen[56]),
			.cell_state(gen[56])
		); 

/******************* CELL 57 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell57 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[116]),
			.N(gen[117]),
			.NE(gen[118]),

			.O(gen[56]),
			.E(gen[58]),

			.SO(gen[116]),
			.S(gen[117]),
			.SE(gen[118]),

			.SELF(gen[57]),
			.cell_state(gen[57])
		); 

/******************* CELL 58 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell58 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[117]),
			.N(gen[118]),
			.NE(gen[119]),

			.O(gen[57]),
			.E(gen[59]),

			.SO(gen[117]),
			.S(gen[118]),
			.SE(gen[119]),

			.SELF(gen[58]),
			.cell_state(gen[58])
		); 

/******************* CELL 59 ***************/  

	CELDA   #(.ic(0), .top_row(1), .bottom_row(0))

		cell59 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[118]),
			.N(gen[119]),
			.NE(gen[118]),

			.O(gen[58]),
			.E(gen[58]),

			.SO(gen[118]),
			.S(gen[119]),
			.SE(gen[118]),

			.SELF(gen[59]),
			.cell_state(gen[59])
		); 

/******************* CELL 60 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell60 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1]),
			.N(gen[0]),
			.NE(gen[1]),

			.O(gen[61]),
			.E(gen[61]),

			.SO(gen[121]),
			.S(gen[120]),
			.SE(gen[121]),

			.SELF(gen[60]),
			.cell_state(gen[60])
		); 

/******************* CELL 61 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell61 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[0]),
			.N(gen[1]),
			.NE(gen[2]),

			.O(gen[60]),
			.E(gen[62]),

			.SO(gen[120]),
			.S(gen[121]),
			.SE(gen[122]),

			.SELF(gen[61]),
			.cell_state(gen[61])
		); 

/******************* CELL 62 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell62 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1]),
			.N(gen[2]),
			.NE(gen[3]),

			.O(gen[61]),
			.E(gen[63]),

			.SO(gen[121]),
			.S(gen[122]),
			.SE(gen[123]),

			.SELF(gen[62]),
			.cell_state(gen[62])
		); 

/******************* CELL 63 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell63 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2]),
			.N(gen[3]),
			.NE(gen[4]),

			.O(gen[62]),
			.E(gen[64]),

			.SO(gen[122]),
			.S(gen[123]),
			.SE(gen[124]),

			.SELF(gen[63]),
			.cell_state(gen[63])
		); 

/******************* CELL 64 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell64 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3]),
			.N(gen[4]),
			.NE(gen[5]),

			.O(gen[63]),
			.E(gen[65]),

			.SO(gen[123]),
			.S(gen[124]),
			.SE(gen[125]),

			.SELF(gen[64]),
			.cell_state(gen[64])
		); 

/******************* CELL 65 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell65 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[4]),
			.N(gen[5]),
			.NE(gen[6]),

			.O(gen[64]),
			.E(gen[66]),

			.SO(gen[124]),
			.S(gen[125]),
			.SE(gen[126]),

			.SELF(gen[65]),
			.cell_state(gen[65])
		); 

/******************* CELL 66 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell66 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[5]),
			.N(gen[6]),
			.NE(gen[7]),

			.O(gen[65]),
			.E(gen[67]),

			.SO(gen[125]),
			.S(gen[126]),
			.SE(gen[127]),

			.SELF(gen[66]),
			.cell_state(gen[66])
		); 

/******************* CELL 67 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell67 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[6]),
			.N(gen[7]),
			.NE(gen[8]),

			.O(gen[66]),
			.E(gen[68]),

			.SO(gen[126]),
			.S(gen[127]),
			.SE(gen[128]),

			.SELF(gen[67]),
			.cell_state(gen[67])
		); 

/******************* CELL 68 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell68 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[7]),
			.N(gen[8]),
			.NE(gen[9]),

			.O(gen[67]),
			.E(gen[69]),

			.SO(gen[127]),
			.S(gen[128]),
			.SE(gen[129]),

			.SELF(gen[68]),
			.cell_state(gen[68])
		); 

/******************* CELL 69 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell69 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[8]),
			.N(gen[9]),
			.NE(gen[10]),

			.O(gen[68]),
			.E(gen[70]),

			.SO(gen[128]),
			.S(gen[129]),
			.SE(gen[130]),

			.SELF(gen[69]),
			.cell_state(gen[69])
		); 

/******************* CELL 70 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell70 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[9]),
			.N(gen[10]),
			.NE(gen[11]),

			.O(gen[69]),
			.E(gen[71]),

			.SO(gen[129]),
			.S(gen[130]),
			.SE(gen[131]),

			.SELF(gen[70]),
			.cell_state(gen[70])
		); 

/******************* CELL 71 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell71 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[10]),
			.N(gen[11]),
			.NE(gen[12]),

			.O(gen[70]),
			.E(gen[72]),

			.SO(gen[130]),
			.S(gen[131]),
			.SE(gen[132]),

			.SELF(gen[71]),
			.cell_state(gen[71])
		); 

/******************* CELL 72 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell72 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[11]),
			.N(gen[12]),
			.NE(gen[13]),

			.O(gen[71]),
			.E(gen[73]),

			.SO(gen[131]),
			.S(gen[132]),
			.SE(gen[133]),

			.SELF(gen[72]),
			.cell_state(gen[72])
		); 

/******************* CELL 73 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell73 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[12]),
			.N(gen[13]),
			.NE(gen[14]),

			.O(gen[72]),
			.E(gen[74]),

			.SO(gen[132]),
			.S(gen[133]),
			.SE(gen[134]),

			.SELF(gen[73]),
			.cell_state(gen[73])
		); 

/******************* CELL 74 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell74 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[13]),
			.N(gen[14]),
			.NE(gen[15]),

			.O(gen[73]),
			.E(gen[75]),

			.SO(gen[133]),
			.S(gen[134]),
			.SE(gen[135]),

			.SELF(gen[74]),
			.cell_state(gen[74])
		); 

/******************* CELL 75 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell75 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[14]),
			.N(gen[15]),
			.NE(gen[16]),

			.O(gen[74]),
			.E(gen[76]),

			.SO(gen[134]),
			.S(gen[135]),
			.SE(gen[136]),

			.SELF(gen[75]),
			.cell_state(gen[75])
		); 

/******************* CELL 76 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell76 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[15]),
			.N(gen[16]),
			.NE(gen[17]),

			.O(gen[75]),
			.E(gen[77]),

			.SO(gen[135]),
			.S(gen[136]),
			.SE(gen[137]),

			.SELF(gen[76]),
			.cell_state(gen[76])
		); 

/******************* CELL 77 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell77 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[16]),
			.N(gen[17]),
			.NE(gen[18]),

			.O(gen[76]),
			.E(gen[78]),

			.SO(gen[136]),
			.S(gen[137]),
			.SE(gen[138]),

			.SELF(gen[77]),
			.cell_state(gen[77])
		); 

/******************* CELL 78 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell78 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[17]),
			.N(gen[18]),
			.NE(gen[19]),

			.O(gen[77]),
			.E(gen[79]),

			.SO(gen[137]),
			.S(gen[138]),
			.SE(gen[139]),

			.SELF(gen[78]),
			.cell_state(gen[78])
		); 

/******************* CELL 79 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell79 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[18]),
			.N(gen[19]),
			.NE(gen[20]),

			.O(gen[78]),
			.E(gen[80]),

			.SO(gen[138]),
			.S(gen[139]),
			.SE(gen[140]),

			.SELF(gen[79]),
			.cell_state(gen[79])
		); 

/******************* CELL 80 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell80 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[19]),
			.N(gen[20]),
			.NE(gen[21]),

			.O(gen[79]),
			.E(gen[81]),

			.SO(gen[139]),
			.S(gen[140]),
			.SE(gen[141]),

			.SELF(gen[80]),
			.cell_state(gen[80])
		); 

/******************* CELL 81 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell81 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[20]),
			.N(gen[21]),
			.NE(gen[22]),

			.O(gen[80]),
			.E(gen[82]),

			.SO(gen[140]),
			.S(gen[141]),
			.SE(gen[142]),

			.SELF(gen[81]),
			.cell_state(gen[81])
		); 

/******************* CELL 82 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell82 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[21]),
			.N(gen[22]),
			.NE(gen[23]),

			.O(gen[81]),
			.E(gen[83]),

			.SO(gen[141]),
			.S(gen[142]),
			.SE(gen[143]),

			.SELF(gen[82]),
			.cell_state(gen[82])
		); 

/******************* CELL 83 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell83 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[22]),
			.N(gen[23]),
			.NE(gen[24]),

			.O(gen[82]),
			.E(gen[84]),

			.SO(gen[142]),
			.S(gen[143]),
			.SE(gen[144]),

			.SELF(gen[83]),
			.cell_state(gen[83])
		); 

/******************* CELL 84 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell84 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[23]),
			.N(gen[24]),
			.NE(gen[25]),

			.O(gen[83]),
			.E(gen[85]),

			.SO(gen[143]),
			.S(gen[144]),
			.SE(gen[145]),

			.SELF(gen[84]),
			.cell_state(gen[84])
		); 

/******************* CELL 85 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell85 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[24]),
			.N(gen[25]),
			.NE(gen[26]),

			.O(gen[84]),
			.E(gen[86]),

			.SO(gen[144]),
			.S(gen[145]),
			.SE(gen[146]),

			.SELF(gen[85]),
			.cell_state(gen[85])
		); 

/******************* CELL 86 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell86 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[25]),
			.N(gen[26]),
			.NE(gen[27]),

			.O(gen[85]),
			.E(gen[87]),

			.SO(gen[145]),
			.S(gen[146]),
			.SE(gen[147]),

			.SELF(gen[86]),
			.cell_state(gen[86])
		); 

/******************* CELL 87 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell87 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[26]),
			.N(gen[27]),
			.NE(gen[28]),

			.O(gen[86]),
			.E(gen[88]),

			.SO(gen[146]),
			.S(gen[147]),
			.SE(gen[148]),

			.SELF(gen[87]),
			.cell_state(gen[87])
		); 

/******************* CELL 88 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell88 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[27]),
			.N(gen[28]),
			.NE(gen[29]),

			.O(gen[87]),
			.E(gen[89]),

			.SO(gen[147]),
			.S(gen[148]),
			.SE(gen[149]),

			.SELF(gen[88]),
			.cell_state(gen[88])
		); 

/******************* CELL 89 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell89 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[28]),
			.N(gen[29]),
			.NE(gen[30]),

			.O(gen[88]),
			.E(gen[90]),

			.SO(gen[148]),
			.S(gen[149]),
			.SE(gen[150]),

			.SELF(gen[89]),
			.cell_state(gen[89])
		); 

/******************* CELL 90 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell90 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[29]),
			.N(gen[30]),
			.NE(gen[31]),

			.O(gen[89]),
			.E(gen[91]),

			.SO(gen[149]),
			.S(gen[150]),
			.SE(gen[151]),

			.SELF(gen[90]),
			.cell_state(gen[90])
		); 

/******************* CELL 91 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell91 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[30]),
			.N(gen[31]),
			.NE(gen[32]),

			.O(gen[90]),
			.E(gen[92]),

			.SO(gen[150]),
			.S(gen[151]),
			.SE(gen[152]),

			.SELF(gen[91]),
			.cell_state(gen[91])
		); 

/******************* CELL 92 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell92 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[31]),
			.N(gen[32]),
			.NE(gen[33]),

			.O(gen[91]),
			.E(gen[93]),

			.SO(gen[151]),
			.S(gen[152]),
			.SE(gen[153]),

			.SELF(gen[92]),
			.cell_state(gen[92])
		); 

/******************* CELL 93 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell93 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[32]),
			.N(gen[33]),
			.NE(gen[34]),

			.O(gen[92]),
			.E(gen[94]),

			.SO(gen[152]),
			.S(gen[153]),
			.SE(gen[154]),

			.SELF(gen[93]),
			.cell_state(gen[93])
		); 

/******************* CELL 94 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell94 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[33]),
			.N(gen[34]),
			.NE(gen[35]),

			.O(gen[93]),
			.E(gen[95]),

			.SO(gen[153]),
			.S(gen[154]),
			.SE(gen[155]),

			.SELF(gen[94]),
			.cell_state(gen[94])
		); 

/******************* CELL 95 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell95 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[34]),
			.N(gen[35]),
			.NE(gen[36]),

			.O(gen[94]),
			.E(gen[96]),

			.SO(gen[154]),
			.S(gen[155]),
			.SE(gen[156]),

			.SELF(gen[95]),
			.cell_state(gen[95])
		); 

/******************* CELL 96 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell96 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[35]),
			.N(gen[36]),
			.NE(gen[37]),

			.O(gen[95]),
			.E(gen[97]),

			.SO(gen[155]),
			.S(gen[156]),
			.SE(gen[157]),

			.SELF(gen[96]),
			.cell_state(gen[96])
		); 

/******************* CELL 97 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell97 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[36]),
			.N(gen[37]),
			.NE(gen[38]),

			.O(gen[96]),
			.E(gen[98]),

			.SO(gen[156]),
			.S(gen[157]),
			.SE(gen[158]),

			.SELF(gen[97]),
			.cell_state(gen[97])
		); 

/******************* CELL 98 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell98 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[37]),
			.N(gen[38]),
			.NE(gen[39]),

			.O(gen[97]),
			.E(gen[99]),

			.SO(gen[157]),
			.S(gen[158]),
			.SE(gen[159]),

			.SELF(gen[98]),
			.cell_state(gen[98])
		); 

/******************* CELL 99 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell99 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[38]),
			.N(gen[39]),
			.NE(gen[40]),

			.O(gen[98]),
			.E(gen[100]),

			.SO(gen[158]),
			.S(gen[159]),
			.SE(gen[160]),

			.SELF(gen[99]),
			.cell_state(gen[99])
		); 

/******************* CELL 100 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell100 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[39]),
			.N(gen[40]),
			.NE(gen[41]),

			.O(gen[99]),
			.E(gen[101]),

			.SO(gen[159]),
			.S(gen[160]),
			.SE(gen[161]),

			.SELF(gen[100]),
			.cell_state(gen[100])
		); 

/******************* CELL 101 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell101 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[40]),
			.N(gen[41]),
			.NE(gen[42]),

			.O(gen[100]),
			.E(gen[102]),

			.SO(gen[160]),
			.S(gen[161]),
			.SE(gen[162]),

			.SELF(gen[101]),
			.cell_state(gen[101])
		); 

/******************* CELL 102 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell102 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[41]),
			.N(gen[42]),
			.NE(gen[43]),

			.O(gen[101]),
			.E(gen[103]),

			.SO(gen[161]),
			.S(gen[162]),
			.SE(gen[163]),

			.SELF(gen[102]),
			.cell_state(gen[102])
		); 

/******************* CELL 103 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell103 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[42]),
			.N(gen[43]),
			.NE(gen[44]),

			.O(gen[102]),
			.E(gen[104]),

			.SO(gen[162]),
			.S(gen[163]),
			.SE(gen[164]),

			.SELF(gen[103]),
			.cell_state(gen[103])
		); 

/******************* CELL 104 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell104 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[43]),
			.N(gen[44]),
			.NE(gen[45]),

			.O(gen[103]),
			.E(gen[105]),

			.SO(gen[163]),
			.S(gen[164]),
			.SE(gen[165]),

			.SELF(gen[104]),
			.cell_state(gen[104])
		); 

/******************* CELL 105 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell105 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[44]),
			.N(gen[45]),
			.NE(gen[46]),

			.O(gen[104]),
			.E(gen[106]),

			.SO(gen[164]),
			.S(gen[165]),
			.SE(gen[166]),

			.SELF(gen[105]),
			.cell_state(gen[105])
		); 

/******************* CELL 106 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell106 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[45]),
			.N(gen[46]),
			.NE(gen[47]),

			.O(gen[105]),
			.E(gen[107]),

			.SO(gen[165]),
			.S(gen[166]),
			.SE(gen[167]),

			.SELF(gen[106]),
			.cell_state(gen[106])
		); 

/******************* CELL 107 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell107 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[46]),
			.N(gen[47]),
			.NE(gen[48]),

			.O(gen[106]),
			.E(gen[108]),

			.SO(gen[166]),
			.S(gen[167]),
			.SE(gen[168]),

			.SELF(gen[107]),
			.cell_state(gen[107])
		); 

/******************* CELL 108 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell108 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[47]),
			.N(gen[48]),
			.NE(gen[49]),

			.O(gen[107]),
			.E(gen[109]),

			.SO(gen[167]),
			.S(gen[168]),
			.SE(gen[169]),

			.SELF(gen[108]),
			.cell_state(gen[108])
		); 

/******************* CELL 109 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell109 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[48]),
			.N(gen[49]),
			.NE(gen[50]),

			.O(gen[108]),
			.E(gen[110]),

			.SO(gen[168]),
			.S(gen[169]),
			.SE(gen[170]),

			.SELF(gen[109]),
			.cell_state(gen[109])
		); 

/******************* CELL 110 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell110 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[49]),
			.N(gen[50]),
			.NE(gen[51]),

			.O(gen[109]),
			.E(gen[111]),

			.SO(gen[169]),
			.S(gen[170]),
			.SE(gen[171]),

			.SELF(gen[110]),
			.cell_state(gen[110])
		); 

/******************* CELL 111 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell111 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[50]),
			.N(gen[51]),
			.NE(gen[52]),

			.O(gen[110]),
			.E(gen[112]),

			.SO(gen[170]),
			.S(gen[171]),
			.SE(gen[172]),

			.SELF(gen[111]),
			.cell_state(gen[111])
		); 

/******************* CELL 112 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell112 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[51]),
			.N(gen[52]),
			.NE(gen[53]),

			.O(gen[111]),
			.E(gen[113]),

			.SO(gen[171]),
			.S(gen[172]),
			.SE(gen[173]),

			.SELF(gen[112]),
			.cell_state(gen[112])
		); 

/******************* CELL 113 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell113 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[52]),
			.N(gen[53]),
			.NE(gen[54]),

			.O(gen[112]),
			.E(gen[114]),

			.SO(gen[172]),
			.S(gen[173]),
			.SE(gen[174]),

			.SELF(gen[113]),
			.cell_state(gen[113])
		); 

/******************* CELL 114 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell114 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[53]),
			.N(gen[54]),
			.NE(gen[55]),

			.O(gen[113]),
			.E(gen[115]),

			.SO(gen[173]),
			.S(gen[174]),
			.SE(gen[175]),

			.SELF(gen[114]),
			.cell_state(gen[114])
		); 

/******************* CELL 115 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell115 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[54]),
			.N(gen[55]),
			.NE(gen[56]),

			.O(gen[114]),
			.E(gen[116]),

			.SO(gen[174]),
			.S(gen[175]),
			.SE(gen[176]),

			.SELF(gen[115]),
			.cell_state(gen[115])
		); 

/******************* CELL 116 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell116 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[55]),
			.N(gen[56]),
			.NE(gen[57]),

			.O(gen[115]),
			.E(gen[117]),

			.SO(gen[175]),
			.S(gen[176]),
			.SE(gen[177]),

			.SELF(gen[116]),
			.cell_state(gen[116])
		); 

/******************* CELL 117 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell117 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[56]),
			.N(gen[57]),
			.NE(gen[58]),

			.O(gen[116]),
			.E(gen[118]),

			.SO(gen[176]),
			.S(gen[177]),
			.SE(gen[178]),

			.SELF(gen[117]),
			.cell_state(gen[117])
		); 

/******************* CELL 118 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell118 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[57]),
			.N(gen[58]),
			.NE(gen[59]),

			.O(gen[117]),
			.E(gen[119]),

			.SO(gen[177]),
			.S(gen[178]),
			.SE(gen[179]),

			.SELF(gen[118]),
			.cell_state(gen[118])
		); 

/******************* CELL 119 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell119 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[58]),
			.N(gen[59]),
			.NE(gen[58]),

			.O(gen[118]),
			.E(gen[118]),

			.SO(gen[178]),
			.S(gen[179]),
			.SE(gen[178]),

			.SELF(gen[119]),
			.cell_state(gen[119])
		); 

/******************* CELL 120 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell120 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[61]),
			.N(gen[60]),
			.NE(gen[61]),

			.O(gen[121]),
			.E(gen[121]),

			.SO(gen[181]),
			.S(gen[180]),
			.SE(gen[181]),

			.SELF(gen[120]),
			.cell_state(gen[120])
		); 

/******************* CELL 121 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell121 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[60]),
			.N(gen[61]),
			.NE(gen[62]),

			.O(gen[120]),
			.E(gen[122]),

			.SO(gen[180]),
			.S(gen[181]),
			.SE(gen[182]),

			.SELF(gen[121]),
			.cell_state(gen[121])
		); 

/******************* CELL 122 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell122 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[61]),
			.N(gen[62]),
			.NE(gen[63]),

			.O(gen[121]),
			.E(gen[123]),

			.SO(gen[181]),
			.S(gen[182]),
			.SE(gen[183]),

			.SELF(gen[122]),
			.cell_state(gen[122])
		); 

/******************* CELL 123 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell123 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[62]),
			.N(gen[63]),
			.NE(gen[64]),

			.O(gen[122]),
			.E(gen[124]),

			.SO(gen[182]),
			.S(gen[183]),
			.SE(gen[184]),

			.SELF(gen[123]),
			.cell_state(gen[123])
		); 

/******************* CELL 124 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell124 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[63]),
			.N(gen[64]),
			.NE(gen[65]),

			.O(gen[123]),
			.E(gen[125]),

			.SO(gen[183]),
			.S(gen[184]),
			.SE(gen[185]),

			.SELF(gen[124]),
			.cell_state(gen[124])
		); 

/******************* CELL 125 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell125 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[64]),
			.N(gen[65]),
			.NE(gen[66]),

			.O(gen[124]),
			.E(gen[126]),

			.SO(gen[184]),
			.S(gen[185]),
			.SE(gen[186]),

			.SELF(gen[125]),
			.cell_state(gen[125])
		); 

/******************* CELL 126 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell126 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[65]),
			.N(gen[66]),
			.NE(gen[67]),

			.O(gen[125]),
			.E(gen[127]),

			.SO(gen[185]),
			.S(gen[186]),
			.SE(gen[187]),

			.SELF(gen[126]),
			.cell_state(gen[126])
		); 

/******************* CELL 127 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell127 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[66]),
			.N(gen[67]),
			.NE(gen[68]),

			.O(gen[126]),
			.E(gen[128]),

			.SO(gen[186]),
			.S(gen[187]),
			.SE(gen[188]),

			.SELF(gen[127]),
			.cell_state(gen[127])
		); 

/******************* CELL 128 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell128 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[67]),
			.N(gen[68]),
			.NE(gen[69]),

			.O(gen[127]),
			.E(gen[129]),

			.SO(gen[187]),
			.S(gen[188]),
			.SE(gen[189]),

			.SELF(gen[128]),
			.cell_state(gen[128])
		); 

/******************* CELL 129 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell129 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[68]),
			.N(gen[69]),
			.NE(gen[70]),

			.O(gen[128]),
			.E(gen[130]),

			.SO(gen[188]),
			.S(gen[189]),
			.SE(gen[190]),

			.SELF(gen[129]),
			.cell_state(gen[129])
		); 

/******************* CELL 130 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell130 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[69]),
			.N(gen[70]),
			.NE(gen[71]),

			.O(gen[129]),
			.E(gen[131]),

			.SO(gen[189]),
			.S(gen[190]),
			.SE(gen[191]),

			.SELF(gen[130]),
			.cell_state(gen[130])
		); 

/******************* CELL 131 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell131 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[70]),
			.N(gen[71]),
			.NE(gen[72]),

			.O(gen[130]),
			.E(gen[132]),

			.SO(gen[190]),
			.S(gen[191]),
			.SE(gen[192]),

			.SELF(gen[131]),
			.cell_state(gen[131])
		); 

/******************* CELL 132 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell132 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[71]),
			.N(gen[72]),
			.NE(gen[73]),

			.O(gen[131]),
			.E(gen[133]),

			.SO(gen[191]),
			.S(gen[192]),
			.SE(gen[193]),

			.SELF(gen[132]),
			.cell_state(gen[132])
		); 

/******************* CELL 133 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell133 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[72]),
			.N(gen[73]),
			.NE(gen[74]),

			.O(gen[132]),
			.E(gen[134]),

			.SO(gen[192]),
			.S(gen[193]),
			.SE(gen[194]),

			.SELF(gen[133]),
			.cell_state(gen[133])
		); 

/******************* CELL 134 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell134 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[73]),
			.N(gen[74]),
			.NE(gen[75]),

			.O(gen[133]),
			.E(gen[135]),

			.SO(gen[193]),
			.S(gen[194]),
			.SE(gen[195]),

			.SELF(gen[134]),
			.cell_state(gen[134])
		); 

/******************* CELL 135 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell135 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[74]),
			.N(gen[75]),
			.NE(gen[76]),

			.O(gen[134]),
			.E(gen[136]),

			.SO(gen[194]),
			.S(gen[195]),
			.SE(gen[196]),

			.SELF(gen[135]),
			.cell_state(gen[135])
		); 

/******************* CELL 136 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell136 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[75]),
			.N(gen[76]),
			.NE(gen[77]),

			.O(gen[135]),
			.E(gen[137]),

			.SO(gen[195]),
			.S(gen[196]),
			.SE(gen[197]),

			.SELF(gen[136]),
			.cell_state(gen[136])
		); 

/******************* CELL 137 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell137 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[76]),
			.N(gen[77]),
			.NE(gen[78]),

			.O(gen[136]),
			.E(gen[138]),

			.SO(gen[196]),
			.S(gen[197]),
			.SE(gen[198]),

			.SELF(gen[137]),
			.cell_state(gen[137])
		); 

/******************* CELL 138 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell138 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[77]),
			.N(gen[78]),
			.NE(gen[79]),

			.O(gen[137]),
			.E(gen[139]),

			.SO(gen[197]),
			.S(gen[198]),
			.SE(gen[199]),

			.SELF(gen[138]),
			.cell_state(gen[138])
		); 

/******************* CELL 139 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell139 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[78]),
			.N(gen[79]),
			.NE(gen[80]),

			.O(gen[138]),
			.E(gen[140]),

			.SO(gen[198]),
			.S(gen[199]),
			.SE(gen[200]),

			.SELF(gen[139]),
			.cell_state(gen[139])
		); 

/******************* CELL 140 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell140 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[79]),
			.N(gen[80]),
			.NE(gen[81]),

			.O(gen[139]),
			.E(gen[141]),

			.SO(gen[199]),
			.S(gen[200]),
			.SE(gen[201]),

			.SELF(gen[140]),
			.cell_state(gen[140])
		); 

/******************* CELL 141 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell141 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[80]),
			.N(gen[81]),
			.NE(gen[82]),

			.O(gen[140]),
			.E(gen[142]),

			.SO(gen[200]),
			.S(gen[201]),
			.SE(gen[202]),

			.SELF(gen[141]),
			.cell_state(gen[141])
		); 

/******************* CELL 142 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell142 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[81]),
			.N(gen[82]),
			.NE(gen[83]),

			.O(gen[141]),
			.E(gen[143]),

			.SO(gen[201]),
			.S(gen[202]),
			.SE(gen[203]),

			.SELF(gen[142]),
			.cell_state(gen[142])
		); 

/******************* CELL 143 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell143 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[82]),
			.N(gen[83]),
			.NE(gen[84]),

			.O(gen[142]),
			.E(gen[144]),

			.SO(gen[202]),
			.S(gen[203]),
			.SE(gen[204]),

			.SELF(gen[143]),
			.cell_state(gen[143])
		); 

/******************* CELL 144 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell144 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[83]),
			.N(gen[84]),
			.NE(gen[85]),

			.O(gen[143]),
			.E(gen[145]),

			.SO(gen[203]),
			.S(gen[204]),
			.SE(gen[205]),

			.SELF(gen[144]),
			.cell_state(gen[144])
		); 

/******************* CELL 145 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell145 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[84]),
			.N(gen[85]),
			.NE(gen[86]),

			.O(gen[144]),
			.E(gen[146]),

			.SO(gen[204]),
			.S(gen[205]),
			.SE(gen[206]),

			.SELF(gen[145]),
			.cell_state(gen[145])
		); 

/******************* CELL 146 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell146 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[85]),
			.N(gen[86]),
			.NE(gen[87]),

			.O(gen[145]),
			.E(gen[147]),

			.SO(gen[205]),
			.S(gen[206]),
			.SE(gen[207]),

			.SELF(gen[146]),
			.cell_state(gen[146])
		); 

/******************* CELL 147 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell147 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[86]),
			.N(gen[87]),
			.NE(gen[88]),

			.O(gen[146]),
			.E(gen[148]),

			.SO(gen[206]),
			.S(gen[207]),
			.SE(gen[208]),

			.SELF(gen[147]),
			.cell_state(gen[147])
		); 

/******************* CELL 148 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell148 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[87]),
			.N(gen[88]),
			.NE(gen[89]),

			.O(gen[147]),
			.E(gen[149]),

			.SO(gen[207]),
			.S(gen[208]),
			.SE(gen[209]),

			.SELF(gen[148]),
			.cell_state(gen[148])
		); 

/******************* CELL 149 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell149 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[88]),
			.N(gen[89]),
			.NE(gen[90]),

			.O(gen[148]),
			.E(gen[150]),

			.SO(gen[208]),
			.S(gen[209]),
			.SE(gen[210]),

			.SELF(gen[149]),
			.cell_state(gen[149])
		); 

/******************* CELL 150 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell150 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[89]),
			.N(gen[90]),
			.NE(gen[91]),

			.O(gen[149]),
			.E(gen[151]),

			.SO(gen[209]),
			.S(gen[210]),
			.SE(gen[211]),

			.SELF(gen[150]),
			.cell_state(gen[150])
		); 

/******************* CELL 151 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell151 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[90]),
			.N(gen[91]),
			.NE(gen[92]),

			.O(gen[150]),
			.E(gen[152]),

			.SO(gen[210]),
			.S(gen[211]),
			.SE(gen[212]),

			.SELF(gen[151]),
			.cell_state(gen[151])
		); 

/******************* CELL 152 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell152 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[91]),
			.N(gen[92]),
			.NE(gen[93]),

			.O(gen[151]),
			.E(gen[153]),

			.SO(gen[211]),
			.S(gen[212]),
			.SE(gen[213]),

			.SELF(gen[152]),
			.cell_state(gen[152])
		); 

/******************* CELL 153 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell153 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[92]),
			.N(gen[93]),
			.NE(gen[94]),

			.O(gen[152]),
			.E(gen[154]),

			.SO(gen[212]),
			.S(gen[213]),
			.SE(gen[214]),

			.SELF(gen[153]),
			.cell_state(gen[153])
		); 

/******************* CELL 154 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell154 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[93]),
			.N(gen[94]),
			.NE(gen[95]),

			.O(gen[153]),
			.E(gen[155]),

			.SO(gen[213]),
			.S(gen[214]),
			.SE(gen[215]),

			.SELF(gen[154]),
			.cell_state(gen[154])
		); 

/******************* CELL 155 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell155 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[94]),
			.N(gen[95]),
			.NE(gen[96]),

			.O(gen[154]),
			.E(gen[156]),

			.SO(gen[214]),
			.S(gen[215]),
			.SE(gen[216]),

			.SELF(gen[155]),
			.cell_state(gen[155])
		); 

/******************* CELL 156 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell156 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[95]),
			.N(gen[96]),
			.NE(gen[97]),

			.O(gen[155]),
			.E(gen[157]),

			.SO(gen[215]),
			.S(gen[216]),
			.SE(gen[217]),

			.SELF(gen[156]),
			.cell_state(gen[156])
		); 

/******************* CELL 157 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell157 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[96]),
			.N(gen[97]),
			.NE(gen[98]),

			.O(gen[156]),
			.E(gen[158]),

			.SO(gen[216]),
			.S(gen[217]),
			.SE(gen[218]),

			.SELF(gen[157]),
			.cell_state(gen[157])
		); 

/******************* CELL 158 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell158 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[97]),
			.N(gen[98]),
			.NE(gen[99]),

			.O(gen[157]),
			.E(gen[159]),

			.SO(gen[217]),
			.S(gen[218]),
			.SE(gen[219]),

			.SELF(gen[158]),
			.cell_state(gen[158])
		); 

/******************* CELL 159 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell159 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[98]),
			.N(gen[99]),
			.NE(gen[100]),

			.O(gen[158]),
			.E(gen[160]),

			.SO(gen[218]),
			.S(gen[219]),
			.SE(gen[220]),

			.SELF(gen[159]),
			.cell_state(gen[159])
		); 

/******************* CELL 160 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell160 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[99]),
			.N(gen[100]),
			.NE(gen[101]),

			.O(gen[159]),
			.E(gen[161]),

			.SO(gen[219]),
			.S(gen[220]),
			.SE(gen[221]),

			.SELF(gen[160]),
			.cell_state(gen[160])
		); 

/******************* CELL 161 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell161 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[100]),
			.N(gen[101]),
			.NE(gen[102]),

			.O(gen[160]),
			.E(gen[162]),

			.SO(gen[220]),
			.S(gen[221]),
			.SE(gen[222]),

			.SELF(gen[161]),
			.cell_state(gen[161])
		); 

/******************* CELL 162 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell162 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[101]),
			.N(gen[102]),
			.NE(gen[103]),

			.O(gen[161]),
			.E(gen[163]),

			.SO(gen[221]),
			.S(gen[222]),
			.SE(gen[223]),

			.SELF(gen[162]),
			.cell_state(gen[162])
		); 

/******************* CELL 163 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell163 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[102]),
			.N(gen[103]),
			.NE(gen[104]),

			.O(gen[162]),
			.E(gen[164]),

			.SO(gen[222]),
			.S(gen[223]),
			.SE(gen[224]),

			.SELF(gen[163]),
			.cell_state(gen[163])
		); 

/******************* CELL 164 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell164 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[103]),
			.N(gen[104]),
			.NE(gen[105]),

			.O(gen[163]),
			.E(gen[165]),

			.SO(gen[223]),
			.S(gen[224]),
			.SE(gen[225]),

			.SELF(gen[164]),
			.cell_state(gen[164])
		); 

/******************* CELL 165 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell165 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[104]),
			.N(gen[105]),
			.NE(gen[106]),

			.O(gen[164]),
			.E(gen[166]),

			.SO(gen[224]),
			.S(gen[225]),
			.SE(gen[226]),

			.SELF(gen[165]),
			.cell_state(gen[165])
		); 

/******************* CELL 166 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell166 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[105]),
			.N(gen[106]),
			.NE(gen[107]),

			.O(gen[165]),
			.E(gen[167]),

			.SO(gen[225]),
			.S(gen[226]),
			.SE(gen[227]),

			.SELF(gen[166]),
			.cell_state(gen[166])
		); 

/******************* CELL 167 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell167 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[106]),
			.N(gen[107]),
			.NE(gen[108]),

			.O(gen[166]),
			.E(gen[168]),

			.SO(gen[226]),
			.S(gen[227]),
			.SE(gen[228]),

			.SELF(gen[167]),
			.cell_state(gen[167])
		); 

/******************* CELL 168 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell168 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[107]),
			.N(gen[108]),
			.NE(gen[109]),

			.O(gen[167]),
			.E(gen[169]),

			.SO(gen[227]),
			.S(gen[228]),
			.SE(gen[229]),

			.SELF(gen[168]),
			.cell_state(gen[168])
		); 

/******************* CELL 169 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell169 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[108]),
			.N(gen[109]),
			.NE(gen[110]),

			.O(gen[168]),
			.E(gen[170]),

			.SO(gen[228]),
			.S(gen[229]),
			.SE(gen[230]),

			.SELF(gen[169]),
			.cell_state(gen[169])
		); 

/******************* CELL 170 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell170 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[109]),
			.N(gen[110]),
			.NE(gen[111]),

			.O(gen[169]),
			.E(gen[171]),

			.SO(gen[229]),
			.S(gen[230]),
			.SE(gen[231]),

			.SELF(gen[170]),
			.cell_state(gen[170])
		); 

/******************* CELL 171 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell171 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[110]),
			.N(gen[111]),
			.NE(gen[112]),

			.O(gen[170]),
			.E(gen[172]),

			.SO(gen[230]),
			.S(gen[231]),
			.SE(gen[232]),

			.SELF(gen[171]),
			.cell_state(gen[171])
		); 

/******************* CELL 172 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell172 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[111]),
			.N(gen[112]),
			.NE(gen[113]),

			.O(gen[171]),
			.E(gen[173]),

			.SO(gen[231]),
			.S(gen[232]),
			.SE(gen[233]),

			.SELF(gen[172]),
			.cell_state(gen[172])
		); 

/******************* CELL 173 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell173 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[112]),
			.N(gen[113]),
			.NE(gen[114]),

			.O(gen[172]),
			.E(gen[174]),

			.SO(gen[232]),
			.S(gen[233]),
			.SE(gen[234]),

			.SELF(gen[173]),
			.cell_state(gen[173])
		); 

/******************* CELL 174 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell174 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[113]),
			.N(gen[114]),
			.NE(gen[115]),

			.O(gen[173]),
			.E(gen[175]),

			.SO(gen[233]),
			.S(gen[234]),
			.SE(gen[235]),

			.SELF(gen[174]),
			.cell_state(gen[174])
		); 

/******************* CELL 175 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell175 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[114]),
			.N(gen[115]),
			.NE(gen[116]),

			.O(gen[174]),
			.E(gen[176]),

			.SO(gen[234]),
			.S(gen[235]),
			.SE(gen[236]),

			.SELF(gen[175]),
			.cell_state(gen[175])
		); 

/******************* CELL 176 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell176 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[115]),
			.N(gen[116]),
			.NE(gen[117]),

			.O(gen[175]),
			.E(gen[177]),

			.SO(gen[235]),
			.S(gen[236]),
			.SE(gen[237]),

			.SELF(gen[176]),
			.cell_state(gen[176])
		); 

/******************* CELL 177 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell177 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[116]),
			.N(gen[117]),
			.NE(gen[118]),

			.O(gen[176]),
			.E(gen[178]),

			.SO(gen[236]),
			.S(gen[237]),
			.SE(gen[238]),

			.SELF(gen[177]),
			.cell_state(gen[177])
		); 

/******************* CELL 178 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell178 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[117]),
			.N(gen[118]),
			.NE(gen[119]),

			.O(gen[177]),
			.E(gen[179]),

			.SO(gen[237]),
			.S(gen[238]),
			.SE(gen[239]),

			.SELF(gen[178]),
			.cell_state(gen[178])
		); 

/******************* CELL 179 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell179 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[118]),
			.N(gen[119]),
			.NE(gen[118]),

			.O(gen[178]),
			.E(gen[178]),

			.SO(gen[238]),
			.S(gen[239]),
			.SE(gen[238]),

			.SELF(gen[179]),
			.cell_state(gen[179])
		); 

/******************* CELL 180 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell180 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[121]),
			.N(gen[120]),
			.NE(gen[121]),

			.O(gen[181]),
			.E(gen[181]),

			.SO(gen[241]),
			.S(gen[240]),
			.SE(gen[241]),

			.SELF(gen[180]),
			.cell_state(gen[180])
		); 

/******************* CELL 181 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell181 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[120]),
			.N(gen[121]),
			.NE(gen[122]),

			.O(gen[180]),
			.E(gen[182]),

			.SO(gen[240]),
			.S(gen[241]),
			.SE(gen[242]),

			.SELF(gen[181]),
			.cell_state(gen[181])
		); 

/******************* CELL 182 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell182 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[121]),
			.N(gen[122]),
			.NE(gen[123]),

			.O(gen[181]),
			.E(gen[183]),

			.SO(gen[241]),
			.S(gen[242]),
			.SE(gen[243]),

			.SELF(gen[182]),
			.cell_state(gen[182])
		); 

/******************* CELL 183 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell183 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[122]),
			.N(gen[123]),
			.NE(gen[124]),

			.O(gen[182]),
			.E(gen[184]),

			.SO(gen[242]),
			.S(gen[243]),
			.SE(gen[244]),

			.SELF(gen[183]),
			.cell_state(gen[183])
		); 

/******************* CELL 184 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell184 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[123]),
			.N(gen[124]),
			.NE(gen[125]),

			.O(gen[183]),
			.E(gen[185]),

			.SO(gen[243]),
			.S(gen[244]),
			.SE(gen[245]),

			.SELF(gen[184]),
			.cell_state(gen[184])
		); 

/******************* CELL 185 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell185 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[124]),
			.N(gen[125]),
			.NE(gen[126]),

			.O(gen[184]),
			.E(gen[186]),

			.SO(gen[244]),
			.S(gen[245]),
			.SE(gen[246]),

			.SELF(gen[185]),
			.cell_state(gen[185])
		); 

/******************* CELL 186 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell186 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[125]),
			.N(gen[126]),
			.NE(gen[127]),

			.O(gen[185]),
			.E(gen[187]),

			.SO(gen[245]),
			.S(gen[246]),
			.SE(gen[247]),

			.SELF(gen[186]),
			.cell_state(gen[186])
		); 

/******************* CELL 187 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell187 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[126]),
			.N(gen[127]),
			.NE(gen[128]),

			.O(gen[186]),
			.E(gen[188]),

			.SO(gen[246]),
			.S(gen[247]),
			.SE(gen[248]),

			.SELF(gen[187]),
			.cell_state(gen[187])
		); 

/******************* CELL 188 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell188 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[127]),
			.N(gen[128]),
			.NE(gen[129]),

			.O(gen[187]),
			.E(gen[189]),

			.SO(gen[247]),
			.S(gen[248]),
			.SE(gen[249]),

			.SELF(gen[188]),
			.cell_state(gen[188])
		); 

/******************* CELL 189 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell189 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[128]),
			.N(gen[129]),
			.NE(gen[130]),

			.O(gen[188]),
			.E(gen[190]),

			.SO(gen[248]),
			.S(gen[249]),
			.SE(gen[250]),

			.SELF(gen[189]),
			.cell_state(gen[189])
		); 

/******************* CELL 190 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell190 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[129]),
			.N(gen[130]),
			.NE(gen[131]),

			.O(gen[189]),
			.E(gen[191]),

			.SO(gen[249]),
			.S(gen[250]),
			.SE(gen[251]),

			.SELF(gen[190]),
			.cell_state(gen[190])
		); 

/******************* CELL 191 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell191 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[130]),
			.N(gen[131]),
			.NE(gen[132]),

			.O(gen[190]),
			.E(gen[192]),

			.SO(gen[250]),
			.S(gen[251]),
			.SE(gen[252]),

			.SELF(gen[191]),
			.cell_state(gen[191])
		); 

/******************* CELL 192 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell192 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[131]),
			.N(gen[132]),
			.NE(gen[133]),

			.O(gen[191]),
			.E(gen[193]),

			.SO(gen[251]),
			.S(gen[252]),
			.SE(gen[253]),

			.SELF(gen[192]),
			.cell_state(gen[192])
		); 

/******************* CELL 193 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell193 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[132]),
			.N(gen[133]),
			.NE(gen[134]),

			.O(gen[192]),
			.E(gen[194]),

			.SO(gen[252]),
			.S(gen[253]),
			.SE(gen[254]),

			.SELF(gen[193]),
			.cell_state(gen[193])
		); 

/******************* CELL 194 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell194 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[133]),
			.N(gen[134]),
			.NE(gen[135]),

			.O(gen[193]),
			.E(gen[195]),

			.SO(gen[253]),
			.S(gen[254]),
			.SE(gen[255]),

			.SELF(gen[194]),
			.cell_state(gen[194])
		); 

/******************* CELL 195 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell195 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[134]),
			.N(gen[135]),
			.NE(gen[136]),

			.O(gen[194]),
			.E(gen[196]),

			.SO(gen[254]),
			.S(gen[255]),
			.SE(gen[256]),

			.SELF(gen[195]),
			.cell_state(gen[195])
		); 

/******************* CELL 196 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell196 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[135]),
			.N(gen[136]),
			.NE(gen[137]),

			.O(gen[195]),
			.E(gen[197]),

			.SO(gen[255]),
			.S(gen[256]),
			.SE(gen[257]),

			.SELF(gen[196]),
			.cell_state(gen[196])
		); 

/******************* CELL 197 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell197 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[136]),
			.N(gen[137]),
			.NE(gen[138]),

			.O(gen[196]),
			.E(gen[198]),

			.SO(gen[256]),
			.S(gen[257]),
			.SE(gen[258]),

			.SELF(gen[197]),
			.cell_state(gen[197])
		); 

/******************* CELL 198 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell198 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[137]),
			.N(gen[138]),
			.NE(gen[139]),

			.O(gen[197]),
			.E(gen[199]),

			.SO(gen[257]),
			.S(gen[258]),
			.SE(gen[259]),

			.SELF(gen[198]),
			.cell_state(gen[198])
		); 

/******************* CELL 199 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell199 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[138]),
			.N(gen[139]),
			.NE(gen[140]),

			.O(gen[198]),
			.E(gen[200]),

			.SO(gen[258]),
			.S(gen[259]),
			.SE(gen[260]),

			.SELF(gen[199]),
			.cell_state(gen[199])
		); 

/******************* CELL 200 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell200 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[139]),
			.N(gen[140]),
			.NE(gen[141]),

			.O(gen[199]),
			.E(gen[201]),

			.SO(gen[259]),
			.S(gen[260]),
			.SE(gen[261]),

			.SELF(gen[200]),
			.cell_state(gen[200])
		); 

/******************* CELL 201 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell201 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[140]),
			.N(gen[141]),
			.NE(gen[142]),

			.O(gen[200]),
			.E(gen[202]),

			.SO(gen[260]),
			.S(gen[261]),
			.SE(gen[262]),

			.SELF(gen[201]),
			.cell_state(gen[201])
		); 

/******************* CELL 202 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell202 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[141]),
			.N(gen[142]),
			.NE(gen[143]),

			.O(gen[201]),
			.E(gen[203]),

			.SO(gen[261]),
			.S(gen[262]),
			.SE(gen[263]),

			.SELF(gen[202]),
			.cell_state(gen[202])
		); 

/******************* CELL 203 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell203 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[142]),
			.N(gen[143]),
			.NE(gen[144]),

			.O(gen[202]),
			.E(gen[204]),

			.SO(gen[262]),
			.S(gen[263]),
			.SE(gen[264]),

			.SELF(gen[203]),
			.cell_state(gen[203])
		); 

/******************* CELL 204 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell204 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[143]),
			.N(gen[144]),
			.NE(gen[145]),

			.O(gen[203]),
			.E(gen[205]),

			.SO(gen[263]),
			.S(gen[264]),
			.SE(gen[265]),

			.SELF(gen[204]),
			.cell_state(gen[204])
		); 

/******************* CELL 205 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell205 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[144]),
			.N(gen[145]),
			.NE(gen[146]),

			.O(gen[204]),
			.E(gen[206]),

			.SO(gen[264]),
			.S(gen[265]),
			.SE(gen[266]),

			.SELF(gen[205]),
			.cell_state(gen[205])
		); 

/******************* CELL 206 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell206 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[145]),
			.N(gen[146]),
			.NE(gen[147]),

			.O(gen[205]),
			.E(gen[207]),

			.SO(gen[265]),
			.S(gen[266]),
			.SE(gen[267]),

			.SELF(gen[206]),
			.cell_state(gen[206])
		); 

/******************* CELL 207 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell207 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[146]),
			.N(gen[147]),
			.NE(gen[148]),

			.O(gen[206]),
			.E(gen[208]),

			.SO(gen[266]),
			.S(gen[267]),
			.SE(gen[268]),

			.SELF(gen[207]),
			.cell_state(gen[207])
		); 

/******************* CELL 208 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell208 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[147]),
			.N(gen[148]),
			.NE(gen[149]),

			.O(gen[207]),
			.E(gen[209]),

			.SO(gen[267]),
			.S(gen[268]),
			.SE(gen[269]),

			.SELF(gen[208]),
			.cell_state(gen[208])
		); 

/******************* CELL 209 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell209 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[148]),
			.N(gen[149]),
			.NE(gen[150]),

			.O(gen[208]),
			.E(gen[210]),

			.SO(gen[268]),
			.S(gen[269]),
			.SE(gen[270]),

			.SELF(gen[209]),
			.cell_state(gen[209])
		); 

/******************* CELL 210 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell210 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[149]),
			.N(gen[150]),
			.NE(gen[151]),

			.O(gen[209]),
			.E(gen[211]),

			.SO(gen[269]),
			.S(gen[270]),
			.SE(gen[271]),

			.SELF(gen[210]),
			.cell_state(gen[210])
		); 

/******************* CELL 211 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell211 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[150]),
			.N(gen[151]),
			.NE(gen[152]),

			.O(gen[210]),
			.E(gen[212]),

			.SO(gen[270]),
			.S(gen[271]),
			.SE(gen[272]),

			.SELF(gen[211]),
			.cell_state(gen[211])
		); 

/******************* CELL 212 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell212 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[151]),
			.N(gen[152]),
			.NE(gen[153]),

			.O(gen[211]),
			.E(gen[213]),

			.SO(gen[271]),
			.S(gen[272]),
			.SE(gen[273]),

			.SELF(gen[212]),
			.cell_state(gen[212])
		); 

/******************* CELL 213 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell213 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[152]),
			.N(gen[153]),
			.NE(gen[154]),

			.O(gen[212]),
			.E(gen[214]),

			.SO(gen[272]),
			.S(gen[273]),
			.SE(gen[274]),

			.SELF(gen[213]),
			.cell_state(gen[213])
		); 

/******************* CELL 214 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell214 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[153]),
			.N(gen[154]),
			.NE(gen[155]),

			.O(gen[213]),
			.E(gen[215]),

			.SO(gen[273]),
			.S(gen[274]),
			.SE(gen[275]),

			.SELF(gen[214]),
			.cell_state(gen[214])
		); 

/******************* CELL 215 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell215 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[154]),
			.N(gen[155]),
			.NE(gen[156]),

			.O(gen[214]),
			.E(gen[216]),

			.SO(gen[274]),
			.S(gen[275]),
			.SE(gen[276]),

			.SELF(gen[215]),
			.cell_state(gen[215])
		); 

/******************* CELL 216 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell216 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[155]),
			.N(gen[156]),
			.NE(gen[157]),

			.O(gen[215]),
			.E(gen[217]),

			.SO(gen[275]),
			.S(gen[276]),
			.SE(gen[277]),

			.SELF(gen[216]),
			.cell_state(gen[216])
		); 

/******************* CELL 217 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell217 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[156]),
			.N(gen[157]),
			.NE(gen[158]),

			.O(gen[216]),
			.E(gen[218]),

			.SO(gen[276]),
			.S(gen[277]),
			.SE(gen[278]),

			.SELF(gen[217]),
			.cell_state(gen[217])
		); 

/******************* CELL 218 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell218 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[157]),
			.N(gen[158]),
			.NE(gen[159]),

			.O(gen[217]),
			.E(gen[219]),

			.SO(gen[277]),
			.S(gen[278]),
			.SE(gen[279]),

			.SELF(gen[218]),
			.cell_state(gen[218])
		); 

/******************* CELL 219 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell219 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[158]),
			.N(gen[159]),
			.NE(gen[160]),

			.O(gen[218]),
			.E(gen[220]),

			.SO(gen[278]),
			.S(gen[279]),
			.SE(gen[280]),

			.SELF(gen[219]),
			.cell_state(gen[219])
		); 

/******************* CELL 220 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell220 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[159]),
			.N(gen[160]),
			.NE(gen[161]),

			.O(gen[219]),
			.E(gen[221]),

			.SO(gen[279]),
			.S(gen[280]),
			.SE(gen[281]),

			.SELF(gen[220]),
			.cell_state(gen[220])
		); 

/******************* CELL 221 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell221 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[160]),
			.N(gen[161]),
			.NE(gen[162]),

			.O(gen[220]),
			.E(gen[222]),

			.SO(gen[280]),
			.S(gen[281]),
			.SE(gen[282]),

			.SELF(gen[221]),
			.cell_state(gen[221])
		); 

/******************* CELL 222 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell222 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[161]),
			.N(gen[162]),
			.NE(gen[163]),

			.O(gen[221]),
			.E(gen[223]),

			.SO(gen[281]),
			.S(gen[282]),
			.SE(gen[283]),

			.SELF(gen[222]),
			.cell_state(gen[222])
		); 

/******************* CELL 223 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell223 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[162]),
			.N(gen[163]),
			.NE(gen[164]),

			.O(gen[222]),
			.E(gen[224]),

			.SO(gen[282]),
			.S(gen[283]),
			.SE(gen[284]),

			.SELF(gen[223]),
			.cell_state(gen[223])
		); 

/******************* CELL 224 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell224 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[163]),
			.N(gen[164]),
			.NE(gen[165]),

			.O(gen[223]),
			.E(gen[225]),

			.SO(gen[283]),
			.S(gen[284]),
			.SE(gen[285]),

			.SELF(gen[224]),
			.cell_state(gen[224])
		); 

/******************* CELL 225 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell225 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[164]),
			.N(gen[165]),
			.NE(gen[166]),

			.O(gen[224]),
			.E(gen[226]),

			.SO(gen[284]),
			.S(gen[285]),
			.SE(gen[286]),

			.SELF(gen[225]),
			.cell_state(gen[225])
		); 

/******************* CELL 226 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell226 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[165]),
			.N(gen[166]),
			.NE(gen[167]),

			.O(gen[225]),
			.E(gen[227]),

			.SO(gen[285]),
			.S(gen[286]),
			.SE(gen[287]),

			.SELF(gen[226]),
			.cell_state(gen[226])
		); 

/******************* CELL 227 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell227 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[166]),
			.N(gen[167]),
			.NE(gen[168]),

			.O(gen[226]),
			.E(gen[228]),

			.SO(gen[286]),
			.S(gen[287]),
			.SE(gen[288]),

			.SELF(gen[227]),
			.cell_state(gen[227])
		); 

/******************* CELL 228 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell228 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[167]),
			.N(gen[168]),
			.NE(gen[169]),

			.O(gen[227]),
			.E(gen[229]),

			.SO(gen[287]),
			.S(gen[288]),
			.SE(gen[289]),

			.SELF(gen[228]),
			.cell_state(gen[228])
		); 

/******************* CELL 229 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell229 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[168]),
			.N(gen[169]),
			.NE(gen[170]),

			.O(gen[228]),
			.E(gen[230]),

			.SO(gen[288]),
			.S(gen[289]),
			.SE(gen[290]),

			.SELF(gen[229]),
			.cell_state(gen[229])
		); 

/******************* CELL 230 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell230 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[169]),
			.N(gen[170]),
			.NE(gen[171]),

			.O(gen[229]),
			.E(gen[231]),

			.SO(gen[289]),
			.S(gen[290]),
			.SE(gen[291]),

			.SELF(gen[230]),
			.cell_state(gen[230])
		); 

/******************* CELL 231 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell231 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[170]),
			.N(gen[171]),
			.NE(gen[172]),

			.O(gen[230]),
			.E(gen[232]),

			.SO(gen[290]),
			.S(gen[291]),
			.SE(gen[292]),

			.SELF(gen[231]),
			.cell_state(gen[231])
		); 

/******************* CELL 232 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell232 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[171]),
			.N(gen[172]),
			.NE(gen[173]),

			.O(gen[231]),
			.E(gen[233]),

			.SO(gen[291]),
			.S(gen[292]),
			.SE(gen[293]),

			.SELF(gen[232]),
			.cell_state(gen[232])
		); 

/******************* CELL 233 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell233 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[172]),
			.N(gen[173]),
			.NE(gen[174]),

			.O(gen[232]),
			.E(gen[234]),

			.SO(gen[292]),
			.S(gen[293]),
			.SE(gen[294]),

			.SELF(gen[233]),
			.cell_state(gen[233])
		); 

/******************* CELL 234 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell234 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[173]),
			.N(gen[174]),
			.NE(gen[175]),

			.O(gen[233]),
			.E(gen[235]),

			.SO(gen[293]),
			.S(gen[294]),
			.SE(gen[295]),

			.SELF(gen[234]),
			.cell_state(gen[234])
		); 

/******************* CELL 235 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell235 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[174]),
			.N(gen[175]),
			.NE(gen[176]),

			.O(gen[234]),
			.E(gen[236]),

			.SO(gen[294]),
			.S(gen[295]),
			.SE(gen[296]),

			.SELF(gen[235]),
			.cell_state(gen[235])
		); 

/******************* CELL 236 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell236 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[175]),
			.N(gen[176]),
			.NE(gen[177]),

			.O(gen[235]),
			.E(gen[237]),

			.SO(gen[295]),
			.S(gen[296]),
			.SE(gen[297]),

			.SELF(gen[236]),
			.cell_state(gen[236])
		); 

/******************* CELL 237 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell237 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[176]),
			.N(gen[177]),
			.NE(gen[178]),

			.O(gen[236]),
			.E(gen[238]),

			.SO(gen[296]),
			.S(gen[297]),
			.SE(gen[298]),

			.SELF(gen[237]),
			.cell_state(gen[237])
		); 

/******************* CELL 238 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell238 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[177]),
			.N(gen[178]),
			.NE(gen[179]),

			.O(gen[237]),
			.E(gen[239]),

			.SO(gen[297]),
			.S(gen[298]),
			.SE(gen[299]),

			.SELF(gen[238]),
			.cell_state(gen[238])
		); 

/******************* CELL 239 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell239 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[178]),
			.N(gen[179]),
			.NE(gen[178]),

			.O(gen[238]),
			.E(gen[238]),

			.SO(gen[298]),
			.S(gen[299]),
			.SE(gen[298]),

			.SELF(gen[239]),
			.cell_state(gen[239])
		); 

/******************* CELL 240 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell240 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[181]),
			.N(gen[180]),
			.NE(gen[181]),

			.O(gen[241]),
			.E(gen[241]),

			.SO(gen[301]),
			.S(gen[300]),
			.SE(gen[301]),

			.SELF(gen[240]),
			.cell_state(gen[240])
		); 

/******************* CELL 241 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell241 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[180]),
			.N(gen[181]),
			.NE(gen[182]),

			.O(gen[240]),
			.E(gen[242]),

			.SO(gen[300]),
			.S(gen[301]),
			.SE(gen[302]),

			.SELF(gen[241]),
			.cell_state(gen[241])
		); 

/******************* CELL 242 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell242 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[181]),
			.N(gen[182]),
			.NE(gen[183]),

			.O(gen[241]),
			.E(gen[243]),

			.SO(gen[301]),
			.S(gen[302]),
			.SE(gen[303]),

			.SELF(gen[242]),
			.cell_state(gen[242])
		); 

/******************* CELL 243 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell243 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[182]),
			.N(gen[183]),
			.NE(gen[184]),

			.O(gen[242]),
			.E(gen[244]),

			.SO(gen[302]),
			.S(gen[303]),
			.SE(gen[304]),

			.SELF(gen[243]),
			.cell_state(gen[243])
		); 

/******************* CELL 244 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell244 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[183]),
			.N(gen[184]),
			.NE(gen[185]),

			.O(gen[243]),
			.E(gen[245]),

			.SO(gen[303]),
			.S(gen[304]),
			.SE(gen[305]),

			.SELF(gen[244]),
			.cell_state(gen[244])
		); 

/******************* CELL 245 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell245 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[184]),
			.N(gen[185]),
			.NE(gen[186]),

			.O(gen[244]),
			.E(gen[246]),

			.SO(gen[304]),
			.S(gen[305]),
			.SE(gen[306]),

			.SELF(gen[245]),
			.cell_state(gen[245])
		); 

/******************* CELL 246 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell246 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[185]),
			.N(gen[186]),
			.NE(gen[187]),

			.O(gen[245]),
			.E(gen[247]),

			.SO(gen[305]),
			.S(gen[306]),
			.SE(gen[307]),

			.SELF(gen[246]),
			.cell_state(gen[246])
		); 

/******************* CELL 247 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell247 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[186]),
			.N(gen[187]),
			.NE(gen[188]),

			.O(gen[246]),
			.E(gen[248]),

			.SO(gen[306]),
			.S(gen[307]),
			.SE(gen[308]),

			.SELF(gen[247]),
			.cell_state(gen[247])
		); 

/******************* CELL 248 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell248 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[187]),
			.N(gen[188]),
			.NE(gen[189]),

			.O(gen[247]),
			.E(gen[249]),

			.SO(gen[307]),
			.S(gen[308]),
			.SE(gen[309]),

			.SELF(gen[248]),
			.cell_state(gen[248])
		); 

/******************* CELL 249 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell249 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[188]),
			.N(gen[189]),
			.NE(gen[190]),

			.O(gen[248]),
			.E(gen[250]),

			.SO(gen[308]),
			.S(gen[309]),
			.SE(gen[310]),

			.SELF(gen[249]),
			.cell_state(gen[249])
		); 

/******************* CELL 250 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell250 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[189]),
			.N(gen[190]),
			.NE(gen[191]),

			.O(gen[249]),
			.E(gen[251]),

			.SO(gen[309]),
			.S(gen[310]),
			.SE(gen[311]),

			.SELF(gen[250]),
			.cell_state(gen[250])
		); 

/******************* CELL 251 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell251 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[190]),
			.N(gen[191]),
			.NE(gen[192]),

			.O(gen[250]),
			.E(gen[252]),

			.SO(gen[310]),
			.S(gen[311]),
			.SE(gen[312]),

			.SELF(gen[251]),
			.cell_state(gen[251])
		); 

/******************* CELL 252 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell252 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[191]),
			.N(gen[192]),
			.NE(gen[193]),

			.O(gen[251]),
			.E(gen[253]),

			.SO(gen[311]),
			.S(gen[312]),
			.SE(gen[313]),

			.SELF(gen[252]),
			.cell_state(gen[252])
		); 

/******************* CELL 253 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell253 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[192]),
			.N(gen[193]),
			.NE(gen[194]),

			.O(gen[252]),
			.E(gen[254]),

			.SO(gen[312]),
			.S(gen[313]),
			.SE(gen[314]),

			.SELF(gen[253]),
			.cell_state(gen[253])
		); 

/******************* CELL 254 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell254 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[193]),
			.N(gen[194]),
			.NE(gen[195]),

			.O(gen[253]),
			.E(gen[255]),

			.SO(gen[313]),
			.S(gen[314]),
			.SE(gen[315]),

			.SELF(gen[254]),
			.cell_state(gen[254])
		); 

/******************* CELL 255 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell255 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[194]),
			.N(gen[195]),
			.NE(gen[196]),

			.O(gen[254]),
			.E(gen[256]),

			.SO(gen[314]),
			.S(gen[315]),
			.SE(gen[316]),

			.SELF(gen[255]),
			.cell_state(gen[255])
		); 

/******************* CELL 256 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell256 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[195]),
			.N(gen[196]),
			.NE(gen[197]),

			.O(gen[255]),
			.E(gen[257]),

			.SO(gen[315]),
			.S(gen[316]),
			.SE(gen[317]),

			.SELF(gen[256]),
			.cell_state(gen[256])
		); 

/******************* CELL 257 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell257 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[196]),
			.N(gen[197]),
			.NE(gen[198]),

			.O(gen[256]),
			.E(gen[258]),

			.SO(gen[316]),
			.S(gen[317]),
			.SE(gen[318]),

			.SELF(gen[257]),
			.cell_state(gen[257])
		); 

/******************* CELL 258 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell258 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[197]),
			.N(gen[198]),
			.NE(gen[199]),

			.O(gen[257]),
			.E(gen[259]),

			.SO(gen[317]),
			.S(gen[318]),
			.SE(gen[319]),

			.SELF(gen[258]),
			.cell_state(gen[258])
		); 

/******************* CELL 259 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell259 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[198]),
			.N(gen[199]),
			.NE(gen[200]),

			.O(gen[258]),
			.E(gen[260]),

			.SO(gen[318]),
			.S(gen[319]),
			.SE(gen[320]),

			.SELF(gen[259]),
			.cell_state(gen[259])
		); 

/******************* CELL 260 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell260 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[199]),
			.N(gen[200]),
			.NE(gen[201]),

			.O(gen[259]),
			.E(gen[261]),

			.SO(gen[319]),
			.S(gen[320]),
			.SE(gen[321]),

			.SELF(gen[260]),
			.cell_state(gen[260])
		); 

/******************* CELL 261 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell261 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[200]),
			.N(gen[201]),
			.NE(gen[202]),

			.O(gen[260]),
			.E(gen[262]),

			.SO(gen[320]),
			.S(gen[321]),
			.SE(gen[322]),

			.SELF(gen[261]),
			.cell_state(gen[261])
		); 

/******************* CELL 262 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell262 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[201]),
			.N(gen[202]),
			.NE(gen[203]),

			.O(gen[261]),
			.E(gen[263]),

			.SO(gen[321]),
			.S(gen[322]),
			.SE(gen[323]),

			.SELF(gen[262]),
			.cell_state(gen[262])
		); 

/******************* CELL 263 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell263 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[202]),
			.N(gen[203]),
			.NE(gen[204]),

			.O(gen[262]),
			.E(gen[264]),

			.SO(gen[322]),
			.S(gen[323]),
			.SE(gen[324]),

			.SELF(gen[263]),
			.cell_state(gen[263])
		); 

/******************* CELL 264 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell264 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[203]),
			.N(gen[204]),
			.NE(gen[205]),

			.O(gen[263]),
			.E(gen[265]),

			.SO(gen[323]),
			.S(gen[324]),
			.SE(gen[325]),

			.SELF(gen[264]),
			.cell_state(gen[264])
		); 

/******************* CELL 265 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell265 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[204]),
			.N(gen[205]),
			.NE(gen[206]),

			.O(gen[264]),
			.E(gen[266]),

			.SO(gen[324]),
			.S(gen[325]),
			.SE(gen[326]),

			.SELF(gen[265]),
			.cell_state(gen[265])
		); 

/******************* CELL 266 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell266 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[205]),
			.N(gen[206]),
			.NE(gen[207]),

			.O(gen[265]),
			.E(gen[267]),

			.SO(gen[325]),
			.S(gen[326]),
			.SE(gen[327]),

			.SELF(gen[266]),
			.cell_state(gen[266])
		); 

/******************* CELL 267 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell267 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[206]),
			.N(gen[207]),
			.NE(gen[208]),

			.O(gen[266]),
			.E(gen[268]),

			.SO(gen[326]),
			.S(gen[327]),
			.SE(gen[328]),

			.SELF(gen[267]),
			.cell_state(gen[267])
		); 

/******************* CELL 268 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell268 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[207]),
			.N(gen[208]),
			.NE(gen[209]),

			.O(gen[267]),
			.E(gen[269]),

			.SO(gen[327]),
			.S(gen[328]),
			.SE(gen[329]),

			.SELF(gen[268]),
			.cell_state(gen[268])
		); 

/******************* CELL 269 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell269 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[208]),
			.N(gen[209]),
			.NE(gen[210]),

			.O(gen[268]),
			.E(gen[270]),

			.SO(gen[328]),
			.S(gen[329]),
			.SE(gen[330]),

			.SELF(gen[269]),
			.cell_state(gen[269])
		); 

/******************* CELL 270 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell270 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[209]),
			.N(gen[210]),
			.NE(gen[211]),

			.O(gen[269]),
			.E(gen[271]),

			.SO(gen[329]),
			.S(gen[330]),
			.SE(gen[331]),

			.SELF(gen[270]),
			.cell_state(gen[270])
		); 

/******************* CELL 271 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell271 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[210]),
			.N(gen[211]),
			.NE(gen[212]),

			.O(gen[270]),
			.E(gen[272]),

			.SO(gen[330]),
			.S(gen[331]),
			.SE(gen[332]),

			.SELF(gen[271]),
			.cell_state(gen[271])
		); 

/******************* CELL 272 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell272 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[211]),
			.N(gen[212]),
			.NE(gen[213]),

			.O(gen[271]),
			.E(gen[273]),

			.SO(gen[331]),
			.S(gen[332]),
			.SE(gen[333]),

			.SELF(gen[272]),
			.cell_state(gen[272])
		); 

/******************* CELL 273 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell273 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[212]),
			.N(gen[213]),
			.NE(gen[214]),

			.O(gen[272]),
			.E(gen[274]),

			.SO(gen[332]),
			.S(gen[333]),
			.SE(gen[334]),

			.SELF(gen[273]),
			.cell_state(gen[273])
		); 

/******************* CELL 274 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell274 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[213]),
			.N(gen[214]),
			.NE(gen[215]),

			.O(gen[273]),
			.E(gen[275]),

			.SO(gen[333]),
			.S(gen[334]),
			.SE(gen[335]),

			.SELF(gen[274]),
			.cell_state(gen[274])
		); 

/******************* CELL 275 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell275 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[214]),
			.N(gen[215]),
			.NE(gen[216]),

			.O(gen[274]),
			.E(gen[276]),

			.SO(gen[334]),
			.S(gen[335]),
			.SE(gen[336]),

			.SELF(gen[275]),
			.cell_state(gen[275])
		); 

/******************* CELL 276 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell276 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[215]),
			.N(gen[216]),
			.NE(gen[217]),

			.O(gen[275]),
			.E(gen[277]),

			.SO(gen[335]),
			.S(gen[336]),
			.SE(gen[337]),

			.SELF(gen[276]),
			.cell_state(gen[276])
		); 

/******************* CELL 277 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell277 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[216]),
			.N(gen[217]),
			.NE(gen[218]),

			.O(gen[276]),
			.E(gen[278]),

			.SO(gen[336]),
			.S(gen[337]),
			.SE(gen[338]),

			.SELF(gen[277]),
			.cell_state(gen[277])
		); 

/******************* CELL 278 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell278 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[217]),
			.N(gen[218]),
			.NE(gen[219]),

			.O(gen[277]),
			.E(gen[279]),

			.SO(gen[337]),
			.S(gen[338]),
			.SE(gen[339]),

			.SELF(gen[278]),
			.cell_state(gen[278])
		); 

/******************* CELL 279 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell279 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[218]),
			.N(gen[219]),
			.NE(gen[220]),

			.O(gen[278]),
			.E(gen[280]),

			.SO(gen[338]),
			.S(gen[339]),
			.SE(gen[340]),

			.SELF(gen[279]),
			.cell_state(gen[279])
		); 

/******************* CELL 280 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell280 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[219]),
			.N(gen[220]),
			.NE(gen[221]),

			.O(gen[279]),
			.E(gen[281]),

			.SO(gen[339]),
			.S(gen[340]),
			.SE(gen[341]),

			.SELF(gen[280]),
			.cell_state(gen[280])
		); 

/******************* CELL 281 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell281 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[220]),
			.N(gen[221]),
			.NE(gen[222]),

			.O(gen[280]),
			.E(gen[282]),

			.SO(gen[340]),
			.S(gen[341]),
			.SE(gen[342]),

			.SELF(gen[281]),
			.cell_state(gen[281])
		); 

/******************* CELL 282 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell282 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[221]),
			.N(gen[222]),
			.NE(gen[223]),

			.O(gen[281]),
			.E(gen[283]),

			.SO(gen[341]),
			.S(gen[342]),
			.SE(gen[343]),

			.SELF(gen[282]),
			.cell_state(gen[282])
		); 

/******************* CELL 283 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell283 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[222]),
			.N(gen[223]),
			.NE(gen[224]),

			.O(gen[282]),
			.E(gen[284]),

			.SO(gen[342]),
			.S(gen[343]),
			.SE(gen[344]),

			.SELF(gen[283]),
			.cell_state(gen[283])
		); 

/******************* CELL 284 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell284 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[223]),
			.N(gen[224]),
			.NE(gen[225]),

			.O(gen[283]),
			.E(gen[285]),

			.SO(gen[343]),
			.S(gen[344]),
			.SE(gen[345]),

			.SELF(gen[284]),
			.cell_state(gen[284])
		); 

/******************* CELL 285 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell285 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[224]),
			.N(gen[225]),
			.NE(gen[226]),

			.O(gen[284]),
			.E(gen[286]),

			.SO(gen[344]),
			.S(gen[345]),
			.SE(gen[346]),

			.SELF(gen[285]),
			.cell_state(gen[285])
		); 

/******************* CELL 286 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell286 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[225]),
			.N(gen[226]),
			.NE(gen[227]),

			.O(gen[285]),
			.E(gen[287]),

			.SO(gen[345]),
			.S(gen[346]),
			.SE(gen[347]),

			.SELF(gen[286]),
			.cell_state(gen[286])
		); 

/******************* CELL 287 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell287 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[226]),
			.N(gen[227]),
			.NE(gen[228]),

			.O(gen[286]),
			.E(gen[288]),

			.SO(gen[346]),
			.S(gen[347]),
			.SE(gen[348]),

			.SELF(gen[287]),
			.cell_state(gen[287])
		); 

/******************* CELL 288 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell288 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[227]),
			.N(gen[228]),
			.NE(gen[229]),

			.O(gen[287]),
			.E(gen[289]),

			.SO(gen[347]),
			.S(gen[348]),
			.SE(gen[349]),

			.SELF(gen[288]),
			.cell_state(gen[288])
		); 

/******************* CELL 289 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell289 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[228]),
			.N(gen[229]),
			.NE(gen[230]),

			.O(gen[288]),
			.E(gen[290]),

			.SO(gen[348]),
			.S(gen[349]),
			.SE(gen[350]),

			.SELF(gen[289]),
			.cell_state(gen[289])
		); 

/******************* CELL 290 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell290 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[229]),
			.N(gen[230]),
			.NE(gen[231]),

			.O(gen[289]),
			.E(gen[291]),

			.SO(gen[349]),
			.S(gen[350]),
			.SE(gen[351]),

			.SELF(gen[290]),
			.cell_state(gen[290])
		); 

/******************* CELL 291 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell291 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[230]),
			.N(gen[231]),
			.NE(gen[232]),

			.O(gen[290]),
			.E(gen[292]),

			.SO(gen[350]),
			.S(gen[351]),
			.SE(gen[352]),

			.SELF(gen[291]),
			.cell_state(gen[291])
		); 

/******************* CELL 292 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell292 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[231]),
			.N(gen[232]),
			.NE(gen[233]),

			.O(gen[291]),
			.E(gen[293]),

			.SO(gen[351]),
			.S(gen[352]),
			.SE(gen[353]),

			.SELF(gen[292]),
			.cell_state(gen[292])
		); 

/******************* CELL 293 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell293 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[232]),
			.N(gen[233]),
			.NE(gen[234]),

			.O(gen[292]),
			.E(gen[294]),

			.SO(gen[352]),
			.S(gen[353]),
			.SE(gen[354]),

			.SELF(gen[293]),
			.cell_state(gen[293])
		); 

/******************* CELL 294 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell294 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[233]),
			.N(gen[234]),
			.NE(gen[235]),

			.O(gen[293]),
			.E(gen[295]),

			.SO(gen[353]),
			.S(gen[354]),
			.SE(gen[355]),

			.SELF(gen[294]),
			.cell_state(gen[294])
		); 

/******************* CELL 295 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell295 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[234]),
			.N(gen[235]),
			.NE(gen[236]),

			.O(gen[294]),
			.E(gen[296]),

			.SO(gen[354]),
			.S(gen[355]),
			.SE(gen[356]),

			.SELF(gen[295]),
			.cell_state(gen[295])
		); 

/******************* CELL 296 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell296 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[235]),
			.N(gen[236]),
			.NE(gen[237]),

			.O(gen[295]),
			.E(gen[297]),

			.SO(gen[355]),
			.S(gen[356]),
			.SE(gen[357]),

			.SELF(gen[296]),
			.cell_state(gen[296])
		); 

/******************* CELL 297 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell297 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[236]),
			.N(gen[237]),
			.NE(gen[238]),

			.O(gen[296]),
			.E(gen[298]),

			.SO(gen[356]),
			.S(gen[357]),
			.SE(gen[358]),

			.SELF(gen[297]),
			.cell_state(gen[297])
		); 

/******************* CELL 298 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell298 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[237]),
			.N(gen[238]),
			.NE(gen[239]),

			.O(gen[297]),
			.E(gen[299]),

			.SO(gen[357]),
			.S(gen[358]),
			.SE(gen[359]),

			.SELF(gen[298]),
			.cell_state(gen[298])
		); 

/******************* CELL 299 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell299 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[238]),
			.N(gen[239]),
			.NE(gen[238]),

			.O(gen[298]),
			.E(gen[298]),

			.SO(gen[358]),
			.S(gen[359]),
			.SE(gen[358]),

			.SELF(gen[299]),
			.cell_state(gen[299])
		); 

/******************* CELL 300 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell300 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[241]),
			.N(gen[240]),
			.NE(gen[241]),

			.O(gen[301]),
			.E(gen[301]),

			.SO(gen[361]),
			.S(gen[360]),
			.SE(gen[361]),

			.SELF(gen[300]),
			.cell_state(gen[300])
		); 

/******************* CELL 301 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell301 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[240]),
			.N(gen[241]),
			.NE(gen[242]),

			.O(gen[300]),
			.E(gen[302]),

			.SO(gen[360]),
			.S(gen[361]),
			.SE(gen[362]),

			.SELF(gen[301]),
			.cell_state(gen[301])
		); 

/******************* CELL 302 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell302 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[241]),
			.N(gen[242]),
			.NE(gen[243]),

			.O(gen[301]),
			.E(gen[303]),

			.SO(gen[361]),
			.S(gen[362]),
			.SE(gen[363]),

			.SELF(gen[302]),
			.cell_state(gen[302])
		); 

/******************* CELL 303 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell303 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[242]),
			.N(gen[243]),
			.NE(gen[244]),

			.O(gen[302]),
			.E(gen[304]),

			.SO(gen[362]),
			.S(gen[363]),
			.SE(gen[364]),

			.SELF(gen[303]),
			.cell_state(gen[303])
		); 

/******************* CELL 304 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell304 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[243]),
			.N(gen[244]),
			.NE(gen[245]),

			.O(gen[303]),
			.E(gen[305]),

			.SO(gen[363]),
			.S(gen[364]),
			.SE(gen[365]),

			.SELF(gen[304]),
			.cell_state(gen[304])
		); 

/******************* CELL 305 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell305 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[244]),
			.N(gen[245]),
			.NE(gen[246]),

			.O(gen[304]),
			.E(gen[306]),

			.SO(gen[364]),
			.S(gen[365]),
			.SE(gen[366]),

			.SELF(gen[305]),
			.cell_state(gen[305])
		); 

/******************* CELL 306 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell306 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[245]),
			.N(gen[246]),
			.NE(gen[247]),

			.O(gen[305]),
			.E(gen[307]),

			.SO(gen[365]),
			.S(gen[366]),
			.SE(gen[367]),

			.SELF(gen[306]),
			.cell_state(gen[306])
		); 

/******************* CELL 307 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell307 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[246]),
			.N(gen[247]),
			.NE(gen[248]),

			.O(gen[306]),
			.E(gen[308]),

			.SO(gen[366]),
			.S(gen[367]),
			.SE(gen[368]),

			.SELF(gen[307]),
			.cell_state(gen[307])
		); 

/******************* CELL 308 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell308 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[247]),
			.N(gen[248]),
			.NE(gen[249]),

			.O(gen[307]),
			.E(gen[309]),

			.SO(gen[367]),
			.S(gen[368]),
			.SE(gen[369]),

			.SELF(gen[308]),
			.cell_state(gen[308])
		); 

/******************* CELL 309 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell309 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[248]),
			.N(gen[249]),
			.NE(gen[250]),

			.O(gen[308]),
			.E(gen[310]),

			.SO(gen[368]),
			.S(gen[369]),
			.SE(gen[370]),

			.SELF(gen[309]),
			.cell_state(gen[309])
		); 

/******************* CELL 310 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell310 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[249]),
			.N(gen[250]),
			.NE(gen[251]),

			.O(gen[309]),
			.E(gen[311]),

			.SO(gen[369]),
			.S(gen[370]),
			.SE(gen[371]),

			.SELF(gen[310]),
			.cell_state(gen[310])
		); 

/******************* CELL 311 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell311 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[250]),
			.N(gen[251]),
			.NE(gen[252]),

			.O(gen[310]),
			.E(gen[312]),

			.SO(gen[370]),
			.S(gen[371]),
			.SE(gen[372]),

			.SELF(gen[311]),
			.cell_state(gen[311])
		); 

/******************* CELL 312 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell312 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[251]),
			.N(gen[252]),
			.NE(gen[253]),

			.O(gen[311]),
			.E(gen[313]),

			.SO(gen[371]),
			.S(gen[372]),
			.SE(gen[373]),

			.SELF(gen[312]),
			.cell_state(gen[312])
		); 

/******************* CELL 313 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell313 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[252]),
			.N(gen[253]),
			.NE(gen[254]),

			.O(gen[312]),
			.E(gen[314]),

			.SO(gen[372]),
			.S(gen[373]),
			.SE(gen[374]),

			.SELF(gen[313]),
			.cell_state(gen[313])
		); 

/******************* CELL 314 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell314 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[253]),
			.N(gen[254]),
			.NE(gen[255]),

			.O(gen[313]),
			.E(gen[315]),

			.SO(gen[373]),
			.S(gen[374]),
			.SE(gen[375]),

			.SELF(gen[314]),
			.cell_state(gen[314])
		); 

/******************* CELL 315 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell315 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[254]),
			.N(gen[255]),
			.NE(gen[256]),

			.O(gen[314]),
			.E(gen[316]),

			.SO(gen[374]),
			.S(gen[375]),
			.SE(gen[376]),

			.SELF(gen[315]),
			.cell_state(gen[315])
		); 

/******************* CELL 316 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell316 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[255]),
			.N(gen[256]),
			.NE(gen[257]),

			.O(gen[315]),
			.E(gen[317]),

			.SO(gen[375]),
			.S(gen[376]),
			.SE(gen[377]),

			.SELF(gen[316]),
			.cell_state(gen[316])
		); 

/******************* CELL 317 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell317 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[256]),
			.N(gen[257]),
			.NE(gen[258]),

			.O(gen[316]),
			.E(gen[318]),

			.SO(gen[376]),
			.S(gen[377]),
			.SE(gen[378]),

			.SELF(gen[317]),
			.cell_state(gen[317])
		); 

/******************* CELL 318 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell318 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[257]),
			.N(gen[258]),
			.NE(gen[259]),

			.O(gen[317]),
			.E(gen[319]),

			.SO(gen[377]),
			.S(gen[378]),
			.SE(gen[379]),

			.SELF(gen[318]),
			.cell_state(gen[318])
		); 

/******************* CELL 319 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell319 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[258]),
			.N(gen[259]),
			.NE(gen[260]),

			.O(gen[318]),
			.E(gen[320]),

			.SO(gen[378]),
			.S(gen[379]),
			.SE(gen[380]),

			.SELF(gen[319]),
			.cell_state(gen[319])
		); 

/******************* CELL 320 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell320 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[259]),
			.N(gen[260]),
			.NE(gen[261]),

			.O(gen[319]),
			.E(gen[321]),

			.SO(gen[379]),
			.S(gen[380]),
			.SE(gen[381]),

			.SELF(gen[320]),
			.cell_state(gen[320])
		); 

/******************* CELL 321 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell321 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[260]),
			.N(gen[261]),
			.NE(gen[262]),

			.O(gen[320]),
			.E(gen[322]),

			.SO(gen[380]),
			.S(gen[381]),
			.SE(gen[382]),

			.SELF(gen[321]),
			.cell_state(gen[321])
		); 

/******************* CELL 322 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell322 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[261]),
			.N(gen[262]),
			.NE(gen[263]),

			.O(gen[321]),
			.E(gen[323]),

			.SO(gen[381]),
			.S(gen[382]),
			.SE(gen[383]),

			.SELF(gen[322]),
			.cell_state(gen[322])
		); 

/******************* CELL 323 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell323 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[262]),
			.N(gen[263]),
			.NE(gen[264]),

			.O(gen[322]),
			.E(gen[324]),

			.SO(gen[382]),
			.S(gen[383]),
			.SE(gen[384]),

			.SELF(gen[323]),
			.cell_state(gen[323])
		); 

/******************* CELL 324 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell324 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[263]),
			.N(gen[264]),
			.NE(gen[265]),

			.O(gen[323]),
			.E(gen[325]),

			.SO(gen[383]),
			.S(gen[384]),
			.SE(gen[385]),

			.SELF(gen[324]),
			.cell_state(gen[324])
		); 

/******************* CELL 325 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell325 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[264]),
			.N(gen[265]),
			.NE(gen[266]),

			.O(gen[324]),
			.E(gen[326]),

			.SO(gen[384]),
			.S(gen[385]),
			.SE(gen[386]),

			.SELF(gen[325]),
			.cell_state(gen[325])
		); 

/******************* CELL 326 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell326 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[265]),
			.N(gen[266]),
			.NE(gen[267]),

			.O(gen[325]),
			.E(gen[327]),

			.SO(gen[385]),
			.S(gen[386]),
			.SE(gen[387]),

			.SELF(gen[326]),
			.cell_state(gen[326])
		); 

/******************* CELL 327 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell327 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[266]),
			.N(gen[267]),
			.NE(gen[268]),

			.O(gen[326]),
			.E(gen[328]),

			.SO(gen[386]),
			.S(gen[387]),
			.SE(gen[388]),

			.SELF(gen[327]),
			.cell_state(gen[327])
		); 

/******************* CELL 328 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell328 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[267]),
			.N(gen[268]),
			.NE(gen[269]),

			.O(gen[327]),
			.E(gen[329]),

			.SO(gen[387]),
			.S(gen[388]),
			.SE(gen[389]),

			.SELF(gen[328]),
			.cell_state(gen[328])
		); 

/******************* CELL 329 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell329 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[268]),
			.N(gen[269]),
			.NE(gen[270]),

			.O(gen[328]),
			.E(gen[330]),

			.SO(gen[388]),
			.S(gen[389]),
			.SE(gen[390]),

			.SELF(gen[329]),
			.cell_state(gen[329])
		); 

/******************* CELL 330 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell330 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[269]),
			.N(gen[270]),
			.NE(gen[271]),

			.O(gen[329]),
			.E(gen[331]),

			.SO(gen[389]),
			.S(gen[390]),
			.SE(gen[391]),

			.SELF(gen[330]),
			.cell_state(gen[330])
		); 

/******************* CELL 331 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell331 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[270]),
			.N(gen[271]),
			.NE(gen[272]),

			.O(gen[330]),
			.E(gen[332]),

			.SO(gen[390]),
			.S(gen[391]),
			.SE(gen[392]),

			.SELF(gen[331]),
			.cell_state(gen[331])
		); 

/******************* CELL 332 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell332 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[271]),
			.N(gen[272]),
			.NE(gen[273]),

			.O(gen[331]),
			.E(gen[333]),

			.SO(gen[391]),
			.S(gen[392]),
			.SE(gen[393]),

			.SELF(gen[332]),
			.cell_state(gen[332])
		); 

/******************* CELL 333 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell333 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[272]),
			.N(gen[273]),
			.NE(gen[274]),

			.O(gen[332]),
			.E(gen[334]),

			.SO(gen[392]),
			.S(gen[393]),
			.SE(gen[394]),

			.SELF(gen[333]),
			.cell_state(gen[333])
		); 

/******************* CELL 334 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell334 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[273]),
			.N(gen[274]),
			.NE(gen[275]),

			.O(gen[333]),
			.E(gen[335]),

			.SO(gen[393]),
			.S(gen[394]),
			.SE(gen[395]),

			.SELF(gen[334]),
			.cell_state(gen[334])
		); 

/******************* CELL 335 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell335 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[274]),
			.N(gen[275]),
			.NE(gen[276]),

			.O(gen[334]),
			.E(gen[336]),

			.SO(gen[394]),
			.S(gen[395]),
			.SE(gen[396]),

			.SELF(gen[335]),
			.cell_state(gen[335])
		); 

/******************* CELL 336 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell336 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[275]),
			.N(gen[276]),
			.NE(gen[277]),

			.O(gen[335]),
			.E(gen[337]),

			.SO(gen[395]),
			.S(gen[396]),
			.SE(gen[397]),

			.SELF(gen[336]),
			.cell_state(gen[336])
		); 

/******************* CELL 337 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell337 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[276]),
			.N(gen[277]),
			.NE(gen[278]),

			.O(gen[336]),
			.E(gen[338]),

			.SO(gen[396]),
			.S(gen[397]),
			.SE(gen[398]),

			.SELF(gen[337]),
			.cell_state(gen[337])
		); 

/******************* CELL 338 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell338 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[277]),
			.N(gen[278]),
			.NE(gen[279]),

			.O(gen[337]),
			.E(gen[339]),

			.SO(gen[397]),
			.S(gen[398]),
			.SE(gen[399]),

			.SELF(gen[338]),
			.cell_state(gen[338])
		); 

/******************* CELL 339 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell339 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[278]),
			.N(gen[279]),
			.NE(gen[280]),

			.O(gen[338]),
			.E(gen[340]),

			.SO(gen[398]),
			.S(gen[399]),
			.SE(gen[400]),

			.SELF(gen[339]),
			.cell_state(gen[339])
		); 

/******************* CELL 340 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell340 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[279]),
			.N(gen[280]),
			.NE(gen[281]),

			.O(gen[339]),
			.E(gen[341]),

			.SO(gen[399]),
			.S(gen[400]),
			.SE(gen[401]),

			.SELF(gen[340]),
			.cell_state(gen[340])
		); 

/******************* CELL 341 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell341 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[280]),
			.N(gen[281]),
			.NE(gen[282]),

			.O(gen[340]),
			.E(gen[342]),

			.SO(gen[400]),
			.S(gen[401]),
			.SE(gen[402]),

			.SELF(gen[341]),
			.cell_state(gen[341])
		); 

/******************* CELL 342 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell342 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[281]),
			.N(gen[282]),
			.NE(gen[283]),

			.O(gen[341]),
			.E(gen[343]),

			.SO(gen[401]),
			.S(gen[402]),
			.SE(gen[403]),

			.SELF(gen[342]),
			.cell_state(gen[342])
		); 

/******************* CELL 343 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell343 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[282]),
			.N(gen[283]),
			.NE(gen[284]),

			.O(gen[342]),
			.E(gen[344]),

			.SO(gen[402]),
			.S(gen[403]),
			.SE(gen[404]),

			.SELF(gen[343]),
			.cell_state(gen[343])
		); 

/******************* CELL 344 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell344 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[283]),
			.N(gen[284]),
			.NE(gen[285]),

			.O(gen[343]),
			.E(gen[345]),

			.SO(gen[403]),
			.S(gen[404]),
			.SE(gen[405]),

			.SELF(gen[344]),
			.cell_state(gen[344])
		); 

/******************* CELL 345 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell345 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[284]),
			.N(gen[285]),
			.NE(gen[286]),

			.O(gen[344]),
			.E(gen[346]),

			.SO(gen[404]),
			.S(gen[405]),
			.SE(gen[406]),

			.SELF(gen[345]),
			.cell_state(gen[345])
		); 

/******************* CELL 346 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell346 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[285]),
			.N(gen[286]),
			.NE(gen[287]),

			.O(gen[345]),
			.E(gen[347]),

			.SO(gen[405]),
			.S(gen[406]),
			.SE(gen[407]),

			.SELF(gen[346]),
			.cell_state(gen[346])
		); 

/******************* CELL 347 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell347 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[286]),
			.N(gen[287]),
			.NE(gen[288]),

			.O(gen[346]),
			.E(gen[348]),

			.SO(gen[406]),
			.S(gen[407]),
			.SE(gen[408]),

			.SELF(gen[347]),
			.cell_state(gen[347])
		); 

/******************* CELL 348 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell348 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[287]),
			.N(gen[288]),
			.NE(gen[289]),

			.O(gen[347]),
			.E(gen[349]),

			.SO(gen[407]),
			.S(gen[408]),
			.SE(gen[409]),

			.SELF(gen[348]),
			.cell_state(gen[348])
		); 

/******************* CELL 349 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell349 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[288]),
			.N(gen[289]),
			.NE(gen[290]),

			.O(gen[348]),
			.E(gen[350]),

			.SO(gen[408]),
			.S(gen[409]),
			.SE(gen[410]),

			.SELF(gen[349]),
			.cell_state(gen[349])
		); 

/******************* CELL 350 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell350 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[289]),
			.N(gen[290]),
			.NE(gen[291]),

			.O(gen[349]),
			.E(gen[351]),

			.SO(gen[409]),
			.S(gen[410]),
			.SE(gen[411]),

			.SELF(gen[350]),
			.cell_state(gen[350])
		); 

/******************* CELL 351 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell351 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[290]),
			.N(gen[291]),
			.NE(gen[292]),

			.O(gen[350]),
			.E(gen[352]),

			.SO(gen[410]),
			.S(gen[411]),
			.SE(gen[412]),

			.SELF(gen[351]),
			.cell_state(gen[351])
		); 

/******************* CELL 352 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell352 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[291]),
			.N(gen[292]),
			.NE(gen[293]),

			.O(gen[351]),
			.E(gen[353]),

			.SO(gen[411]),
			.S(gen[412]),
			.SE(gen[413]),

			.SELF(gen[352]),
			.cell_state(gen[352])
		); 

/******************* CELL 353 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell353 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[292]),
			.N(gen[293]),
			.NE(gen[294]),

			.O(gen[352]),
			.E(gen[354]),

			.SO(gen[412]),
			.S(gen[413]),
			.SE(gen[414]),

			.SELF(gen[353]),
			.cell_state(gen[353])
		); 

/******************* CELL 354 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell354 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[293]),
			.N(gen[294]),
			.NE(gen[295]),

			.O(gen[353]),
			.E(gen[355]),

			.SO(gen[413]),
			.S(gen[414]),
			.SE(gen[415]),

			.SELF(gen[354]),
			.cell_state(gen[354])
		); 

/******************* CELL 355 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell355 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[294]),
			.N(gen[295]),
			.NE(gen[296]),

			.O(gen[354]),
			.E(gen[356]),

			.SO(gen[414]),
			.S(gen[415]),
			.SE(gen[416]),

			.SELF(gen[355]),
			.cell_state(gen[355])
		); 

/******************* CELL 356 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell356 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[295]),
			.N(gen[296]),
			.NE(gen[297]),

			.O(gen[355]),
			.E(gen[357]),

			.SO(gen[415]),
			.S(gen[416]),
			.SE(gen[417]),

			.SELF(gen[356]),
			.cell_state(gen[356])
		); 

/******************* CELL 357 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell357 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[296]),
			.N(gen[297]),
			.NE(gen[298]),

			.O(gen[356]),
			.E(gen[358]),

			.SO(gen[416]),
			.S(gen[417]),
			.SE(gen[418]),

			.SELF(gen[357]),
			.cell_state(gen[357])
		); 

/******************* CELL 358 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell358 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[297]),
			.N(gen[298]),
			.NE(gen[299]),

			.O(gen[357]),
			.E(gen[359]),

			.SO(gen[417]),
			.S(gen[418]),
			.SE(gen[419]),

			.SELF(gen[358]),
			.cell_state(gen[358])
		); 

/******************* CELL 359 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell359 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[298]),
			.N(gen[299]),
			.NE(gen[298]),

			.O(gen[358]),
			.E(gen[358]),

			.SO(gen[418]),
			.S(gen[419]),
			.SE(gen[418]),

			.SELF(gen[359]),
			.cell_state(gen[359])
		); 

/******************* CELL 360 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell360 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[301]),
			.N(gen[300]),
			.NE(gen[301]),

			.O(gen[361]),
			.E(gen[361]),

			.SO(gen[421]),
			.S(gen[420]),
			.SE(gen[421]),

			.SELF(gen[360]),
			.cell_state(gen[360])
		); 

/******************* CELL 361 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell361 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[300]),
			.N(gen[301]),
			.NE(gen[302]),

			.O(gen[360]),
			.E(gen[362]),

			.SO(gen[420]),
			.S(gen[421]),
			.SE(gen[422]),

			.SELF(gen[361]),
			.cell_state(gen[361])
		); 

/******************* CELL 362 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell362 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[301]),
			.N(gen[302]),
			.NE(gen[303]),

			.O(gen[361]),
			.E(gen[363]),

			.SO(gen[421]),
			.S(gen[422]),
			.SE(gen[423]),

			.SELF(gen[362]),
			.cell_state(gen[362])
		); 

/******************* CELL 363 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell363 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[302]),
			.N(gen[303]),
			.NE(gen[304]),

			.O(gen[362]),
			.E(gen[364]),

			.SO(gen[422]),
			.S(gen[423]),
			.SE(gen[424]),

			.SELF(gen[363]),
			.cell_state(gen[363])
		); 

/******************* CELL 364 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell364 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[303]),
			.N(gen[304]),
			.NE(gen[305]),

			.O(gen[363]),
			.E(gen[365]),

			.SO(gen[423]),
			.S(gen[424]),
			.SE(gen[425]),

			.SELF(gen[364]),
			.cell_state(gen[364])
		); 

/******************* CELL 365 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell365 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[304]),
			.N(gen[305]),
			.NE(gen[306]),

			.O(gen[364]),
			.E(gen[366]),

			.SO(gen[424]),
			.S(gen[425]),
			.SE(gen[426]),

			.SELF(gen[365]),
			.cell_state(gen[365])
		); 

/******************* CELL 366 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell366 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[305]),
			.N(gen[306]),
			.NE(gen[307]),

			.O(gen[365]),
			.E(gen[367]),

			.SO(gen[425]),
			.S(gen[426]),
			.SE(gen[427]),

			.SELF(gen[366]),
			.cell_state(gen[366])
		); 

/******************* CELL 367 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell367 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[306]),
			.N(gen[307]),
			.NE(gen[308]),

			.O(gen[366]),
			.E(gen[368]),

			.SO(gen[426]),
			.S(gen[427]),
			.SE(gen[428]),

			.SELF(gen[367]),
			.cell_state(gen[367])
		); 

/******************* CELL 368 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell368 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[307]),
			.N(gen[308]),
			.NE(gen[309]),

			.O(gen[367]),
			.E(gen[369]),

			.SO(gen[427]),
			.S(gen[428]),
			.SE(gen[429]),

			.SELF(gen[368]),
			.cell_state(gen[368])
		); 

/******************* CELL 369 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell369 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[308]),
			.N(gen[309]),
			.NE(gen[310]),

			.O(gen[368]),
			.E(gen[370]),

			.SO(gen[428]),
			.S(gen[429]),
			.SE(gen[430]),

			.SELF(gen[369]),
			.cell_state(gen[369])
		); 

/******************* CELL 370 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell370 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[309]),
			.N(gen[310]),
			.NE(gen[311]),

			.O(gen[369]),
			.E(gen[371]),

			.SO(gen[429]),
			.S(gen[430]),
			.SE(gen[431]),

			.SELF(gen[370]),
			.cell_state(gen[370])
		); 

/******************* CELL 371 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell371 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[310]),
			.N(gen[311]),
			.NE(gen[312]),

			.O(gen[370]),
			.E(gen[372]),

			.SO(gen[430]),
			.S(gen[431]),
			.SE(gen[432]),

			.SELF(gen[371]),
			.cell_state(gen[371])
		); 

/******************* CELL 372 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell372 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[311]),
			.N(gen[312]),
			.NE(gen[313]),

			.O(gen[371]),
			.E(gen[373]),

			.SO(gen[431]),
			.S(gen[432]),
			.SE(gen[433]),

			.SELF(gen[372]),
			.cell_state(gen[372])
		); 

/******************* CELL 373 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell373 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[312]),
			.N(gen[313]),
			.NE(gen[314]),

			.O(gen[372]),
			.E(gen[374]),

			.SO(gen[432]),
			.S(gen[433]),
			.SE(gen[434]),

			.SELF(gen[373]),
			.cell_state(gen[373])
		); 

/******************* CELL 374 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell374 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[313]),
			.N(gen[314]),
			.NE(gen[315]),

			.O(gen[373]),
			.E(gen[375]),

			.SO(gen[433]),
			.S(gen[434]),
			.SE(gen[435]),

			.SELF(gen[374]),
			.cell_state(gen[374])
		); 

/******************* CELL 375 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell375 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[314]),
			.N(gen[315]),
			.NE(gen[316]),

			.O(gen[374]),
			.E(gen[376]),

			.SO(gen[434]),
			.S(gen[435]),
			.SE(gen[436]),

			.SELF(gen[375]),
			.cell_state(gen[375])
		); 

/******************* CELL 376 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell376 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[315]),
			.N(gen[316]),
			.NE(gen[317]),

			.O(gen[375]),
			.E(gen[377]),

			.SO(gen[435]),
			.S(gen[436]),
			.SE(gen[437]),

			.SELF(gen[376]),
			.cell_state(gen[376])
		); 

/******************* CELL 377 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell377 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[316]),
			.N(gen[317]),
			.NE(gen[318]),

			.O(gen[376]),
			.E(gen[378]),

			.SO(gen[436]),
			.S(gen[437]),
			.SE(gen[438]),

			.SELF(gen[377]),
			.cell_state(gen[377])
		); 

/******************* CELL 378 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell378 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[317]),
			.N(gen[318]),
			.NE(gen[319]),

			.O(gen[377]),
			.E(gen[379]),

			.SO(gen[437]),
			.S(gen[438]),
			.SE(gen[439]),

			.SELF(gen[378]),
			.cell_state(gen[378])
		); 

/******************* CELL 379 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell379 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[318]),
			.N(gen[319]),
			.NE(gen[320]),

			.O(gen[378]),
			.E(gen[380]),

			.SO(gen[438]),
			.S(gen[439]),
			.SE(gen[440]),

			.SELF(gen[379]),
			.cell_state(gen[379])
		); 

/******************* CELL 380 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell380 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[319]),
			.N(gen[320]),
			.NE(gen[321]),

			.O(gen[379]),
			.E(gen[381]),

			.SO(gen[439]),
			.S(gen[440]),
			.SE(gen[441]),

			.SELF(gen[380]),
			.cell_state(gen[380])
		); 

/******************* CELL 381 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell381 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[320]),
			.N(gen[321]),
			.NE(gen[322]),

			.O(gen[380]),
			.E(gen[382]),

			.SO(gen[440]),
			.S(gen[441]),
			.SE(gen[442]),

			.SELF(gen[381]),
			.cell_state(gen[381])
		); 

/******************* CELL 382 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell382 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[321]),
			.N(gen[322]),
			.NE(gen[323]),

			.O(gen[381]),
			.E(gen[383]),

			.SO(gen[441]),
			.S(gen[442]),
			.SE(gen[443]),

			.SELF(gen[382]),
			.cell_state(gen[382])
		); 

/******************* CELL 383 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell383 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[322]),
			.N(gen[323]),
			.NE(gen[324]),

			.O(gen[382]),
			.E(gen[384]),

			.SO(gen[442]),
			.S(gen[443]),
			.SE(gen[444]),

			.SELF(gen[383]),
			.cell_state(gen[383])
		); 

/******************* CELL 384 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell384 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[323]),
			.N(gen[324]),
			.NE(gen[325]),

			.O(gen[383]),
			.E(gen[385]),

			.SO(gen[443]),
			.S(gen[444]),
			.SE(gen[445]),

			.SELF(gen[384]),
			.cell_state(gen[384])
		); 

/******************* CELL 385 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell385 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[324]),
			.N(gen[325]),
			.NE(gen[326]),

			.O(gen[384]),
			.E(gen[386]),

			.SO(gen[444]),
			.S(gen[445]),
			.SE(gen[446]),

			.SELF(gen[385]),
			.cell_state(gen[385])
		); 

/******************* CELL 386 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell386 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[325]),
			.N(gen[326]),
			.NE(gen[327]),

			.O(gen[385]),
			.E(gen[387]),

			.SO(gen[445]),
			.S(gen[446]),
			.SE(gen[447]),

			.SELF(gen[386]),
			.cell_state(gen[386])
		); 

/******************* CELL 387 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell387 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[326]),
			.N(gen[327]),
			.NE(gen[328]),

			.O(gen[386]),
			.E(gen[388]),

			.SO(gen[446]),
			.S(gen[447]),
			.SE(gen[448]),

			.SELF(gen[387]),
			.cell_state(gen[387])
		); 

/******************* CELL 388 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell388 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[327]),
			.N(gen[328]),
			.NE(gen[329]),

			.O(gen[387]),
			.E(gen[389]),

			.SO(gen[447]),
			.S(gen[448]),
			.SE(gen[449]),

			.SELF(gen[388]),
			.cell_state(gen[388])
		); 

/******************* CELL 389 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell389 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[328]),
			.N(gen[329]),
			.NE(gen[330]),

			.O(gen[388]),
			.E(gen[390]),

			.SO(gen[448]),
			.S(gen[449]),
			.SE(gen[450]),

			.SELF(gen[389]),
			.cell_state(gen[389])
		); 

/******************* CELL 390 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell390 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[329]),
			.N(gen[330]),
			.NE(gen[331]),

			.O(gen[389]),
			.E(gen[391]),

			.SO(gen[449]),
			.S(gen[450]),
			.SE(gen[451]),

			.SELF(gen[390]),
			.cell_state(gen[390])
		); 

/******************* CELL 391 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell391 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[330]),
			.N(gen[331]),
			.NE(gen[332]),

			.O(gen[390]),
			.E(gen[392]),

			.SO(gen[450]),
			.S(gen[451]),
			.SE(gen[452]),

			.SELF(gen[391]),
			.cell_state(gen[391])
		); 

/******************* CELL 392 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell392 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[331]),
			.N(gen[332]),
			.NE(gen[333]),

			.O(gen[391]),
			.E(gen[393]),

			.SO(gen[451]),
			.S(gen[452]),
			.SE(gen[453]),

			.SELF(gen[392]),
			.cell_state(gen[392])
		); 

/******************* CELL 393 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell393 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[332]),
			.N(gen[333]),
			.NE(gen[334]),

			.O(gen[392]),
			.E(gen[394]),

			.SO(gen[452]),
			.S(gen[453]),
			.SE(gen[454]),

			.SELF(gen[393]),
			.cell_state(gen[393])
		); 

/******************* CELL 394 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell394 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[333]),
			.N(gen[334]),
			.NE(gen[335]),

			.O(gen[393]),
			.E(gen[395]),

			.SO(gen[453]),
			.S(gen[454]),
			.SE(gen[455]),

			.SELF(gen[394]),
			.cell_state(gen[394])
		); 

/******************* CELL 395 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell395 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[334]),
			.N(gen[335]),
			.NE(gen[336]),

			.O(gen[394]),
			.E(gen[396]),

			.SO(gen[454]),
			.S(gen[455]),
			.SE(gen[456]),

			.SELF(gen[395]),
			.cell_state(gen[395])
		); 

/******************* CELL 396 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell396 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[335]),
			.N(gen[336]),
			.NE(gen[337]),

			.O(gen[395]),
			.E(gen[397]),

			.SO(gen[455]),
			.S(gen[456]),
			.SE(gen[457]),

			.SELF(gen[396]),
			.cell_state(gen[396])
		); 

/******************* CELL 397 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell397 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[336]),
			.N(gen[337]),
			.NE(gen[338]),

			.O(gen[396]),
			.E(gen[398]),

			.SO(gen[456]),
			.S(gen[457]),
			.SE(gen[458]),

			.SELF(gen[397]),
			.cell_state(gen[397])
		); 

/******************* CELL 398 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell398 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[337]),
			.N(gen[338]),
			.NE(gen[339]),

			.O(gen[397]),
			.E(gen[399]),

			.SO(gen[457]),
			.S(gen[458]),
			.SE(gen[459]),

			.SELF(gen[398]),
			.cell_state(gen[398])
		); 

/******************* CELL 399 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell399 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[338]),
			.N(gen[339]),
			.NE(gen[340]),

			.O(gen[398]),
			.E(gen[400]),

			.SO(gen[458]),
			.S(gen[459]),
			.SE(gen[460]),

			.SELF(gen[399]),
			.cell_state(gen[399])
		); 

/******************* CELL 400 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell400 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[339]),
			.N(gen[340]),
			.NE(gen[341]),

			.O(gen[399]),
			.E(gen[401]),

			.SO(gen[459]),
			.S(gen[460]),
			.SE(gen[461]),

			.SELF(gen[400]),
			.cell_state(gen[400])
		); 

/******************* CELL 401 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell401 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[340]),
			.N(gen[341]),
			.NE(gen[342]),

			.O(gen[400]),
			.E(gen[402]),

			.SO(gen[460]),
			.S(gen[461]),
			.SE(gen[462]),

			.SELF(gen[401]),
			.cell_state(gen[401])
		); 

/******************* CELL 402 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell402 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[341]),
			.N(gen[342]),
			.NE(gen[343]),

			.O(gen[401]),
			.E(gen[403]),

			.SO(gen[461]),
			.S(gen[462]),
			.SE(gen[463]),

			.SELF(gen[402]),
			.cell_state(gen[402])
		); 

/******************* CELL 403 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell403 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[342]),
			.N(gen[343]),
			.NE(gen[344]),

			.O(gen[402]),
			.E(gen[404]),

			.SO(gen[462]),
			.S(gen[463]),
			.SE(gen[464]),

			.SELF(gen[403]),
			.cell_state(gen[403])
		); 

/******************* CELL 404 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell404 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[343]),
			.N(gen[344]),
			.NE(gen[345]),

			.O(gen[403]),
			.E(gen[405]),

			.SO(gen[463]),
			.S(gen[464]),
			.SE(gen[465]),

			.SELF(gen[404]),
			.cell_state(gen[404])
		); 

/******************* CELL 405 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell405 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[344]),
			.N(gen[345]),
			.NE(gen[346]),

			.O(gen[404]),
			.E(gen[406]),

			.SO(gen[464]),
			.S(gen[465]),
			.SE(gen[466]),

			.SELF(gen[405]),
			.cell_state(gen[405])
		); 

/******************* CELL 406 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell406 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[345]),
			.N(gen[346]),
			.NE(gen[347]),

			.O(gen[405]),
			.E(gen[407]),

			.SO(gen[465]),
			.S(gen[466]),
			.SE(gen[467]),

			.SELF(gen[406]),
			.cell_state(gen[406])
		); 

/******************* CELL 407 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell407 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[346]),
			.N(gen[347]),
			.NE(gen[348]),

			.O(gen[406]),
			.E(gen[408]),

			.SO(gen[466]),
			.S(gen[467]),
			.SE(gen[468]),

			.SELF(gen[407]),
			.cell_state(gen[407])
		); 

/******************* CELL 408 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell408 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[347]),
			.N(gen[348]),
			.NE(gen[349]),

			.O(gen[407]),
			.E(gen[409]),

			.SO(gen[467]),
			.S(gen[468]),
			.SE(gen[469]),

			.SELF(gen[408]),
			.cell_state(gen[408])
		); 

/******************* CELL 409 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell409 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[348]),
			.N(gen[349]),
			.NE(gen[350]),

			.O(gen[408]),
			.E(gen[410]),

			.SO(gen[468]),
			.S(gen[469]),
			.SE(gen[470]),

			.SELF(gen[409]),
			.cell_state(gen[409])
		); 

/******************* CELL 410 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell410 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[349]),
			.N(gen[350]),
			.NE(gen[351]),

			.O(gen[409]),
			.E(gen[411]),

			.SO(gen[469]),
			.S(gen[470]),
			.SE(gen[471]),

			.SELF(gen[410]),
			.cell_state(gen[410])
		); 

/******************* CELL 411 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell411 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[350]),
			.N(gen[351]),
			.NE(gen[352]),

			.O(gen[410]),
			.E(gen[412]),

			.SO(gen[470]),
			.S(gen[471]),
			.SE(gen[472]),

			.SELF(gen[411]),
			.cell_state(gen[411])
		); 

/******************* CELL 412 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell412 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[351]),
			.N(gen[352]),
			.NE(gen[353]),

			.O(gen[411]),
			.E(gen[413]),

			.SO(gen[471]),
			.S(gen[472]),
			.SE(gen[473]),

			.SELF(gen[412]),
			.cell_state(gen[412])
		); 

/******************* CELL 413 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell413 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[352]),
			.N(gen[353]),
			.NE(gen[354]),

			.O(gen[412]),
			.E(gen[414]),

			.SO(gen[472]),
			.S(gen[473]),
			.SE(gen[474]),

			.SELF(gen[413]),
			.cell_state(gen[413])
		); 

/******************* CELL 414 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell414 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[353]),
			.N(gen[354]),
			.NE(gen[355]),

			.O(gen[413]),
			.E(gen[415]),

			.SO(gen[473]),
			.S(gen[474]),
			.SE(gen[475]),

			.SELF(gen[414]),
			.cell_state(gen[414])
		); 

/******************* CELL 415 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell415 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[354]),
			.N(gen[355]),
			.NE(gen[356]),

			.O(gen[414]),
			.E(gen[416]),

			.SO(gen[474]),
			.S(gen[475]),
			.SE(gen[476]),

			.SELF(gen[415]),
			.cell_state(gen[415])
		); 

/******************* CELL 416 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell416 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[355]),
			.N(gen[356]),
			.NE(gen[357]),

			.O(gen[415]),
			.E(gen[417]),

			.SO(gen[475]),
			.S(gen[476]),
			.SE(gen[477]),

			.SELF(gen[416]),
			.cell_state(gen[416])
		); 

/******************* CELL 417 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell417 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[356]),
			.N(gen[357]),
			.NE(gen[358]),

			.O(gen[416]),
			.E(gen[418]),

			.SO(gen[476]),
			.S(gen[477]),
			.SE(gen[478]),

			.SELF(gen[417]),
			.cell_state(gen[417])
		); 

/******************* CELL 418 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell418 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[357]),
			.N(gen[358]),
			.NE(gen[359]),

			.O(gen[417]),
			.E(gen[419]),

			.SO(gen[477]),
			.S(gen[478]),
			.SE(gen[479]),

			.SELF(gen[418]),
			.cell_state(gen[418])
		); 

/******************* CELL 419 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell419 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[358]),
			.N(gen[359]),
			.NE(gen[358]),

			.O(gen[418]),
			.E(gen[418]),

			.SO(gen[478]),
			.S(gen[479]),
			.SE(gen[478]),

			.SELF(gen[419]),
			.cell_state(gen[419])
		); 

/******************* CELL 420 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell420 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[361]),
			.N(gen[360]),
			.NE(gen[361]),

			.O(gen[421]),
			.E(gen[421]),

			.SO(gen[481]),
			.S(gen[480]),
			.SE(gen[481]),

			.SELF(gen[420]),
			.cell_state(gen[420])
		); 

/******************* CELL 421 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell421 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[360]),
			.N(gen[361]),
			.NE(gen[362]),

			.O(gen[420]),
			.E(gen[422]),

			.SO(gen[480]),
			.S(gen[481]),
			.SE(gen[482]),

			.SELF(gen[421]),
			.cell_state(gen[421])
		); 

/******************* CELL 422 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell422 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[361]),
			.N(gen[362]),
			.NE(gen[363]),

			.O(gen[421]),
			.E(gen[423]),

			.SO(gen[481]),
			.S(gen[482]),
			.SE(gen[483]),

			.SELF(gen[422]),
			.cell_state(gen[422])
		); 

/******************* CELL 423 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell423 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[362]),
			.N(gen[363]),
			.NE(gen[364]),

			.O(gen[422]),
			.E(gen[424]),

			.SO(gen[482]),
			.S(gen[483]),
			.SE(gen[484]),

			.SELF(gen[423]),
			.cell_state(gen[423])
		); 

/******************* CELL 424 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell424 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[363]),
			.N(gen[364]),
			.NE(gen[365]),

			.O(gen[423]),
			.E(gen[425]),

			.SO(gen[483]),
			.S(gen[484]),
			.SE(gen[485]),

			.SELF(gen[424]),
			.cell_state(gen[424])
		); 

/******************* CELL 425 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell425 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[364]),
			.N(gen[365]),
			.NE(gen[366]),

			.O(gen[424]),
			.E(gen[426]),

			.SO(gen[484]),
			.S(gen[485]),
			.SE(gen[486]),

			.SELF(gen[425]),
			.cell_state(gen[425])
		); 

/******************* CELL 426 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell426 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[365]),
			.N(gen[366]),
			.NE(gen[367]),

			.O(gen[425]),
			.E(gen[427]),

			.SO(gen[485]),
			.S(gen[486]),
			.SE(gen[487]),

			.SELF(gen[426]),
			.cell_state(gen[426])
		); 

/******************* CELL 427 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell427 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[366]),
			.N(gen[367]),
			.NE(gen[368]),

			.O(gen[426]),
			.E(gen[428]),

			.SO(gen[486]),
			.S(gen[487]),
			.SE(gen[488]),

			.SELF(gen[427]),
			.cell_state(gen[427])
		); 

/******************* CELL 428 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell428 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[367]),
			.N(gen[368]),
			.NE(gen[369]),

			.O(gen[427]),
			.E(gen[429]),

			.SO(gen[487]),
			.S(gen[488]),
			.SE(gen[489]),

			.SELF(gen[428]),
			.cell_state(gen[428])
		); 

/******************* CELL 429 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell429 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[368]),
			.N(gen[369]),
			.NE(gen[370]),

			.O(gen[428]),
			.E(gen[430]),

			.SO(gen[488]),
			.S(gen[489]),
			.SE(gen[490]),

			.SELF(gen[429]),
			.cell_state(gen[429])
		); 

/******************* CELL 430 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell430 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[369]),
			.N(gen[370]),
			.NE(gen[371]),

			.O(gen[429]),
			.E(gen[431]),

			.SO(gen[489]),
			.S(gen[490]),
			.SE(gen[491]),

			.SELF(gen[430]),
			.cell_state(gen[430])
		); 

/******************* CELL 431 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell431 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[370]),
			.N(gen[371]),
			.NE(gen[372]),

			.O(gen[430]),
			.E(gen[432]),

			.SO(gen[490]),
			.S(gen[491]),
			.SE(gen[492]),

			.SELF(gen[431]),
			.cell_state(gen[431])
		); 

/******************* CELL 432 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell432 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[371]),
			.N(gen[372]),
			.NE(gen[373]),

			.O(gen[431]),
			.E(gen[433]),

			.SO(gen[491]),
			.S(gen[492]),
			.SE(gen[493]),

			.SELF(gen[432]),
			.cell_state(gen[432])
		); 

/******************* CELL 433 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell433 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[372]),
			.N(gen[373]),
			.NE(gen[374]),

			.O(gen[432]),
			.E(gen[434]),

			.SO(gen[492]),
			.S(gen[493]),
			.SE(gen[494]),

			.SELF(gen[433]),
			.cell_state(gen[433])
		); 

/******************* CELL 434 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell434 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[373]),
			.N(gen[374]),
			.NE(gen[375]),

			.O(gen[433]),
			.E(gen[435]),

			.SO(gen[493]),
			.S(gen[494]),
			.SE(gen[495]),

			.SELF(gen[434]),
			.cell_state(gen[434])
		); 

/******************* CELL 435 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell435 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[374]),
			.N(gen[375]),
			.NE(gen[376]),

			.O(gen[434]),
			.E(gen[436]),

			.SO(gen[494]),
			.S(gen[495]),
			.SE(gen[496]),

			.SELF(gen[435]),
			.cell_state(gen[435])
		); 

/******************* CELL 436 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell436 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[375]),
			.N(gen[376]),
			.NE(gen[377]),

			.O(gen[435]),
			.E(gen[437]),

			.SO(gen[495]),
			.S(gen[496]),
			.SE(gen[497]),

			.SELF(gen[436]),
			.cell_state(gen[436])
		); 

/******************* CELL 437 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell437 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[376]),
			.N(gen[377]),
			.NE(gen[378]),

			.O(gen[436]),
			.E(gen[438]),

			.SO(gen[496]),
			.S(gen[497]),
			.SE(gen[498]),

			.SELF(gen[437]),
			.cell_state(gen[437])
		); 

/******************* CELL 438 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell438 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[377]),
			.N(gen[378]),
			.NE(gen[379]),

			.O(gen[437]),
			.E(gen[439]),

			.SO(gen[497]),
			.S(gen[498]),
			.SE(gen[499]),

			.SELF(gen[438]),
			.cell_state(gen[438])
		); 

/******************* CELL 439 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell439 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[378]),
			.N(gen[379]),
			.NE(gen[380]),

			.O(gen[438]),
			.E(gen[440]),

			.SO(gen[498]),
			.S(gen[499]),
			.SE(gen[500]),

			.SELF(gen[439]),
			.cell_state(gen[439])
		); 

/******************* CELL 440 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell440 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[379]),
			.N(gen[380]),
			.NE(gen[381]),

			.O(gen[439]),
			.E(gen[441]),

			.SO(gen[499]),
			.S(gen[500]),
			.SE(gen[501]),

			.SELF(gen[440]),
			.cell_state(gen[440])
		); 

/******************* CELL 441 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell441 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[380]),
			.N(gen[381]),
			.NE(gen[382]),

			.O(gen[440]),
			.E(gen[442]),

			.SO(gen[500]),
			.S(gen[501]),
			.SE(gen[502]),

			.SELF(gen[441]),
			.cell_state(gen[441])
		); 

/******************* CELL 442 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell442 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[381]),
			.N(gen[382]),
			.NE(gen[383]),

			.O(gen[441]),
			.E(gen[443]),

			.SO(gen[501]),
			.S(gen[502]),
			.SE(gen[503]),

			.SELF(gen[442]),
			.cell_state(gen[442])
		); 

/******************* CELL 443 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell443 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[382]),
			.N(gen[383]),
			.NE(gen[384]),

			.O(gen[442]),
			.E(gen[444]),

			.SO(gen[502]),
			.S(gen[503]),
			.SE(gen[504]),

			.SELF(gen[443]),
			.cell_state(gen[443])
		); 

/******************* CELL 444 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell444 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[383]),
			.N(gen[384]),
			.NE(gen[385]),

			.O(gen[443]),
			.E(gen[445]),

			.SO(gen[503]),
			.S(gen[504]),
			.SE(gen[505]),

			.SELF(gen[444]),
			.cell_state(gen[444])
		); 

/******************* CELL 445 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell445 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[384]),
			.N(gen[385]),
			.NE(gen[386]),

			.O(gen[444]),
			.E(gen[446]),

			.SO(gen[504]),
			.S(gen[505]),
			.SE(gen[506]),

			.SELF(gen[445]),
			.cell_state(gen[445])
		); 

/******************* CELL 446 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell446 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[385]),
			.N(gen[386]),
			.NE(gen[387]),

			.O(gen[445]),
			.E(gen[447]),

			.SO(gen[505]),
			.S(gen[506]),
			.SE(gen[507]),

			.SELF(gen[446]),
			.cell_state(gen[446])
		); 

/******************* CELL 447 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell447 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[386]),
			.N(gen[387]),
			.NE(gen[388]),

			.O(gen[446]),
			.E(gen[448]),

			.SO(gen[506]),
			.S(gen[507]),
			.SE(gen[508]),

			.SELF(gen[447]),
			.cell_state(gen[447])
		); 

/******************* CELL 448 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell448 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[387]),
			.N(gen[388]),
			.NE(gen[389]),

			.O(gen[447]),
			.E(gen[449]),

			.SO(gen[507]),
			.S(gen[508]),
			.SE(gen[509]),

			.SELF(gen[448]),
			.cell_state(gen[448])
		); 

/******************* CELL 449 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell449 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[388]),
			.N(gen[389]),
			.NE(gen[390]),

			.O(gen[448]),
			.E(gen[450]),

			.SO(gen[508]),
			.S(gen[509]),
			.SE(gen[510]),

			.SELF(gen[449]),
			.cell_state(gen[449])
		); 

/******************* CELL 450 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell450 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[389]),
			.N(gen[390]),
			.NE(gen[391]),

			.O(gen[449]),
			.E(gen[451]),

			.SO(gen[509]),
			.S(gen[510]),
			.SE(gen[511]),

			.SELF(gen[450]),
			.cell_state(gen[450])
		); 

/******************* CELL 451 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell451 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[390]),
			.N(gen[391]),
			.NE(gen[392]),

			.O(gen[450]),
			.E(gen[452]),

			.SO(gen[510]),
			.S(gen[511]),
			.SE(gen[512]),

			.SELF(gen[451]),
			.cell_state(gen[451])
		); 

/******************* CELL 452 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell452 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[391]),
			.N(gen[392]),
			.NE(gen[393]),

			.O(gen[451]),
			.E(gen[453]),

			.SO(gen[511]),
			.S(gen[512]),
			.SE(gen[513]),

			.SELF(gen[452]),
			.cell_state(gen[452])
		); 

/******************* CELL 453 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell453 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[392]),
			.N(gen[393]),
			.NE(gen[394]),

			.O(gen[452]),
			.E(gen[454]),

			.SO(gen[512]),
			.S(gen[513]),
			.SE(gen[514]),

			.SELF(gen[453]),
			.cell_state(gen[453])
		); 

/******************* CELL 454 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell454 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[393]),
			.N(gen[394]),
			.NE(gen[395]),

			.O(gen[453]),
			.E(gen[455]),

			.SO(gen[513]),
			.S(gen[514]),
			.SE(gen[515]),

			.SELF(gen[454]),
			.cell_state(gen[454])
		); 

/******************* CELL 455 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell455 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[394]),
			.N(gen[395]),
			.NE(gen[396]),

			.O(gen[454]),
			.E(gen[456]),

			.SO(gen[514]),
			.S(gen[515]),
			.SE(gen[516]),

			.SELF(gen[455]),
			.cell_state(gen[455])
		); 

/******************* CELL 456 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell456 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[395]),
			.N(gen[396]),
			.NE(gen[397]),

			.O(gen[455]),
			.E(gen[457]),

			.SO(gen[515]),
			.S(gen[516]),
			.SE(gen[517]),

			.SELF(gen[456]),
			.cell_state(gen[456])
		); 

/******************* CELL 457 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell457 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[396]),
			.N(gen[397]),
			.NE(gen[398]),

			.O(gen[456]),
			.E(gen[458]),

			.SO(gen[516]),
			.S(gen[517]),
			.SE(gen[518]),

			.SELF(gen[457]),
			.cell_state(gen[457])
		); 

/******************* CELL 458 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell458 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[397]),
			.N(gen[398]),
			.NE(gen[399]),

			.O(gen[457]),
			.E(gen[459]),

			.SO(gen[517]),
			.S(gen[518]),
			.SE(gen[519]),

			.SELF(gen[458]),
			.cell_state(gen[458])
		); 

/******************* CELL 459 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell459 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[398]),
			.N(gen[399]),
			.NE(gen[400]),

			.O(gen[458]),
			.E(gen[460]),

			.SO(gen[518]),
			.S(gen[519]),
			.SE(gen[520]),

			.SELF(gen[459]),
			.cell_state(gen[459])
		); 

/******************* CELL 460 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell460 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[399]),
			.N(gen[400]),
			.NE(gen[401]),

			.O(gen[459]),
			.E(gen[461]),

			.SO(gen[519]),
			.S(gen[520]),
			.SE(gen[521]),

			.SELF(gen[460]),
			.cell_state(gen[460])
		); 

/******************* CELL 461 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell461 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[400]),
			.N(gen[401]),
			.NE(gen[402]),

			.O(gen[460]),
			.E(gen[462]),

			.SO(gen[520]),
			.S(gen[521]),
			.SE(gen[522]),

			.SELF(gen[461]),
			.cell_state(gen[461])
		); 

/******************* CELL 462 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell462 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[401]),
			.N(gen[402]),
			.NE(gen[403]),

			.O(gen[461]),
			.E(gen[463]),

			.SO(gen[521]),
			.S(gen[522]),
			.SE(gen[523]),

			.SELF(gen[462]),
			.cell_state(gen[462])
		); 

/******************* CELL 463 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell463 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[402]),
			.N(gen[403]),
			.NE(gen[404]),

			.O(gen[462]),
			.E(gen[464]),

			.SO(gen[522]),
			.S(gen[523]),
			.SE(gen[524]),

			.SELF(gen[463]),
			.cell_state(gen[463])
		); 

/******************* CELL 464 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell464 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[403]),
			.N(gen[404]),
			.NE(gen[405]),

			.O(gen[463]),
			.E(gen[465]),

			.SO(gen[523]),
			.S(gen[524]),
			.SE(gen[525]),

			.SELF(gen[464]),
			.cell_state(gen[464])
		); 

/******************* CELL 465 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell465 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[404]),
			.N(gen[405]),
			.NE(gen[406]),

			.O(gen[464]),
			.E(gen[466]),

			.SO(gen[524]),
			.S(gen[525]),
			.SE(gen[526]),

			.SELF(gen[465]),
			.cell_state(gen[465])
		); 

/******************* CELL 466 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell466 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[405]),
			.N(gen[406]),
			.NE(gen[407]),

			.O(gen[465]),
			.E(gen[467]),

			.SO(gen[525]),
			.S(gen[526]),
			.SE(gen[527]),

			.SELF(gen[466]),
			.cell_state(gen[466])
		); 

/******************* CELL 467 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell467 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[406]),
			.N(gen[407]),
			.NE(gen[408]),

			.O(gen[466]),
			.E(gen[468]),

			.SO(gen[526]),
			.S(gen[527]),
			.SE(gen[528]),

			.SELF(gen[467]),
			.cell_state(gen[467])
		); 

/******************* CELL 468 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell468 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[407]),
			.N(gen[408]),
			.NE(gen[409]),

			.O(gen[467]),
			.E(gen[469]),

			.SO(gen[527]),
			.S(gen[528]),
			.SE(gen[529]),

			.SELF(gen[468]),
			.cell_state(gen[468])
		); 

/******************* CELL 469 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell469 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[408]),
			.N(gen[409]),
			.NE(gen[410]),

			.O(gen[468]),
			.E(gen[470]),

			.SO(gen[528]),
			.S(gen[529]),
			.SE(gen[530]),

			.SELF(gen[469]),
			.cell_state(gen[469])
		); 

/******************* CELL 470 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell470 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[409]),
			.N(gen[410]),
			.NE(gen[411]),

			.O(gen[469]),
			.E(gen[471]),

			.SO(gen[529]),
			.S(gen[530]),
			.SE(gen[531]),

			.SELF(gen[470]),
			.cell_state(gen[470])
		); 

/******************* CELL 471 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell471 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[410]),
			.N(gen[411]),
			.NE(gen[412]),

			.O(gen[470]),
			.E(gen[472]),

			.SO(gen[530]),
			.S(gen[531]),
			.SE(gen[532]),

			.SELF(gen[471]),
			.cell_state(gen[471])
		); 

/******************* CELL 472 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell472 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[411]),
			.N(gen[412]),
			.NE(gen[413]),

			.O(gen[471]),
			.E(gen[473]),

			.SO(gen[531]),
			.S(gen[532]),
			.SE(gen[533]),

			.SELF(gen[472]),
			.cell_state(gen[472])
		); 

/******************* CELL 473 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell473 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[412]),
			.N(gen[413]),
			.NE(gen[414]),

			.O(gen[472]),
			.E(gen[474]),

			.SO(gen[532]),
			.S(gen[533]),
			.SE(gen[534]),

			.SELF(gen[473]),
			.cell_state(gen[473])
		); 

/******************* CELL 474 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell474 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[413]),
			.N(gen[414]),
			.NE(gen[415]),

			.O(gen[473]),
			.E(gen[475]),

			.SO(gen[533]),
			.S(gen[534]),
			.SE(gen[535]),

			.SELF(gen[474]),
			.cell_state(gen[474])
		); 

/******************* CELL 475 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell475 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[414]),
			.N(gen[415]),
			.NE(gen[416]),

			.O(gen[474]),
			.E(gen[476]),

			.SO(gen[534]),
			.S(gen[535]),
			.SE(gen[536]),

			.SELF(gen[475]),
			.cell_state(gen[475])
		); 

/******************* CELL 476 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell476 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[415]),
			.N(gen[416]),
			.NE(gen[417]),

			.O(gen[475]),
			.E(gen[477]),

			.SO(gen[535]),
			.S(gen[536]),
			.SE(gen[537]),

			.SELF(gen[476]),
			.cell_state(gen[476])
		); 

/******************* CELL 477 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell477 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[416]),
			.N(gen[417]),
			.NE(gen[418]),

			.O(gen[476]),
			.E(gen[478]),

			.SO(gen[536]),
			.S(gen[537]),
			.SE(gen[538]),

			.SELF(gen[477]),
			.cell_state(gen[477])
		); 

/******************* CELL 478 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell478 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[417]),
			.N(gen[418]),
			.NE(gen[419]),

			.O(gen[477]),
			.E(gen[479]),

			.SO(gen[537]),
			.S(gen[538]),
			.SE(gen[539]),

			.SELF(gen[478]),
			.cell_state(gen[478])
		); 

/******************* CELL 479 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell479 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[418]),
			.N(gen[419]),
			.NE(gen[418]),

			.O(gen[478]),
			.E(gen[478]),

			.SO(gen[538]),
			.S(gen[539]),
			.SE(gen[538]),

			.SELF(gen[479]),
			.cell_state(gen[479])
		); 

/******************* CELL 480 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell480 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[421]),
			.N(gen[420]),
			.NE(gen[421]),

			.O(gen[481]),
			.E(gen[481]),

			.SO(gen[541]),
			.S(gen[540]),
			.SE(gen[541]),

			.SELF(gen[480]),
			.cell_state(gen[480])
		); 

/******************* CELL 481 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell481 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[420]),
			.N(gen[421]),
			.NE(gen[422]),

			.O(gen[480]),
			.E(gen[482]),

			.SO(gen[540]),
			.S(gen[541]),
			.SE(gen[542]),

			.SELF(gen[481]),
			.cell_state(gen[481])
		); 

/******************* CELL 482 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell482 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[421]),
			.N(gen[422]),
			.NE(gen[423]),

			.O(gen[481]),
			.E(gen[483]),

			.SO(gen[541]),
			.S(gen[542]),
			.SE(gen[543]),

			.SELF(gen[482]),
			.cell_state(gen[482])
		); 

/******************* CELL 483 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell483 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[422]),
			.N(gen[423]),
			.NE(gen[424]),

			.O(gen[482]),
			.E(gen[484]),

			.SO(gen[542]),
			.S(gen[543]),
			.SE(gen[544]),

			.SELF(gen[483]),
			.cell_state(gen[483])
		); 

/******************* CELL 484 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell484 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[423]),
			.N(gen[424]),
			.NE(gen[425]),

			.O(gen[483]),
			.E(gen[485]),

			.SO(gen[543]),
			.S(gen[544]),
			.SE(gen[545]),

			.SELF(gen[484]),
			.cell_state(gen[484])
		); 

/******************* CELL 485 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell485 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[424]),
			.N(gen[425]),
			.NE(gen[426]),

			.O(gen[484]),
			.E(gen[486]),

			.SO(gen[544]),
			.S(gen[545]),
			.SE(gen[546]),

			.SELF(gen[485]),
			.cell_state(gen[485])
		); 

/******************* CELL 486 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell486 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[425]),
			.N(gen[426]),
			.NE(gen[427]),

			.O(gen[485]),
			.E(gen[487]),

			.SO(gen[545]),
			.S(gen[546]),
			.SE(gen[547]),

			.SELF(gen[486]),
			.cell_state(gen[486])
		); 

/******************* CELL 487 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell487 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[426]),
			.N(gen[427]),
			.NE(gen[428]),

			.O(gen[486]),
			.E(gen[488]),

			.SO(gen[546]),
			.S(gen[547]),
			.SE(gen[548]),

			.SELF(gen[487]),
			.cell_state(gen[487])
		); 

/******************* CELL 488 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell488 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[427]),
			.N(gen[428]),
			.NE(gen[429]),

			.O(gen[487]),
			.E(gen[489]),

			.SO(gen[547]),
			.S(gen[548]),
			.SE(gen[549]),

			.SELF(gen[488]),
			.cell_state(gen[488])
		); 

/******************* CELL 489 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell489 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[428]),
			.N(gen[429]),
			.NE(gen[430]),

			.O(gen[488]),
			.E(gen[490]),

			.SO(gen[548]),
			.S(gen[549]),
			.SE(gen[550]),

			.SELF(gen[489]),
			.cell_state(gen[489])
		); 

/******************* CELL 490 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell490 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[429]),
			.N(gen[430]),
			.NE(gen[431]),

			.O(gen[489]),
			.E(gen[491]),

			.SO(gen[549]),
			.S(gen[550]),
			.SE(gen[551]),

			.SELF(gen[490]),
			.cell_state(gen[490])
		); 

/******************* CELL 491 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell491 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[430]),
			.N(gen[431]),
			.NE(gen[432]),

			.O(gen[490]),
			.E(gen[492]),

			.SO(gen[550]),
			.S(gen[551]),
			.SE(gen[552]),

			.SELF(gen[491]),
			.cell_state(gen[491])
		); 

/******************* CELL 492 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell492 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[431]),
			.N(gen[432]),
			.NE(gen[433]),

			.O(gen[491]),
			.E(gen[493]),

			.SO(gen[551]),
			.S(gen[552]),
			.SE(gen[553]),

			.SELF(gen[492]),
			.cell_state(gen[492])
		); 

/******************* CELL 493 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell493 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[432]),
			.N(gen[433]),
			.NE(gen[434]),

			.O(gen[492]),
			.E(gen[494]),

			.SO(gen[552]),
			.S(gen[553]),
			.SE(gen[554]),

			.SELF(gen[493]),
			.cell_state(gen[493])
		); 

/******************* CELL 494 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell494 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[433]),
			.N(gen[434]),
			.NE(gen[435]),

			.O(gen[493]),
			.E(gen[495]),

			.SO(gen[553]),
			.S(gen[554]),
			.SE(gen[555]),

			.SELF(gen[494]),
			.cell_state(gen[494])
		); 

/******************* CELL 495 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell495 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[434]),
			.N(gen[435]),
			.NE(gen[436]),

			.O(gen[494]),
			.E(gen[496]),

			.SO(gen[554]),
			.S(gen[555]),
			.SE(gen[556]),

			.SELF(gen[495]),
			.cell_state(gen[495])
		); 

/******************* CELL 496 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell496 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[435]),
			.N(gen[436]),
			.NE(gen[437]),

			.O(gen[495]),
			.E(gen[497]),

			.SO(gen[555]),
			.S(gen[556]),
			.SE(gen[557]),

			.SELF(gen[496]),
			.cell_state(gen[496])
		); 

/******************* CELL 497 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell497 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[436]),
			.N(gen[437]),
			.NE(gen[438]),

			.O(gen[496]),
			.E(gen[498]),

			.SO(gen[556]),
			.S(gen[557]),
			.SE(gen[558]),

			.SELF(gen[497]),
			.cell_state(gen[497])
		); 

/******************* CELL 498 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell498 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[437]),
			.N(gen[438]),
			.NE(gen[439]),

			.O(gen[497]),
			.E(gen[499]),

			.SO(gen[557]),
			.S(gen[558]),
			.SE(gen[559]),

			.SELF(gen[498]),
			.cell_state(gen[498])
		); 

/******************* CELL 499 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell499 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[438]),
			.N(gen[439]),
			.NE(gen[440]),

			.O(gen[498]),
			.E(gen[500]),

			.SO(gen[558]),
			.S(gen[559]),
			.SE(gen[560]),

			.SELF(gen[499]),
			.cell_state(gen[499])
		); 

/******************* CELL 500 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell500 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[439]),
			.N(gen[440]),
			.NE(gen[441]),

			.O(gen[499]),
			.E(gen[501]),

			.SO(gen[559]),
			.S(gen[560]),
			.SE(gen[561]),

			.SELF(gen[500]),
			.cell_state(gen[500])
		); 

/******************* CELL 501 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell501 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[440]),
			.N(gen[441]),
			.NE(gen[442]),

			.O(gen[500]),
			.E(gen[502]),

			.SO(gen[560]),
			.S(gen[561]),
			.SE(gen[562]),

			.SELF(gen[501]),
			.cell_state(gen[501])
		); 

/******************* CELL 502 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell502 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[441]),
			.N(gen[442]),
			.NE(gen[443]),

			.O(gen[501]),
			.E(gen[503]),

			.SO(gen[561]),
			.S(gen[562]),
			.SE(gen[563]),

			.SELF(gen[502]),
			.cell_state(gen[502])
		); 

/******************* CELL 503 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell503 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[442]),
			.N(gen[443]),
			.NE(gen[444]),

			.O(gen[502]),
			.E(gen[504]),

			.SO(gen[562]),
			.S(gen[563]),
			.SE(gen[564]),

			.SELF(gen[503]),
			.cell_state(gen[503])
		); 

/******************* CELL 504 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell504 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[443]),
			.N(gen[444]),
			.NE(gen[445]),

			.O(gen[503]),
			.E(gen[505]),

			.SO(gen[563]),
			.S(gen[564]),
			.SE(gen[565]),

			.SELF(gen[504]),
			.cell_state(gen[504])
		); 

/******************* CELL 505 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell505 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[444]),
			.N(gen[445]),
			.NE(gen[446]),

			.O(gen[504]),
			.E(gen[506]),

			.SO(gen[564]),
			.S(gen[565]),
			.SE(gen[566]),

			.SELF(gen[505]),
			.cell_state(gen[505])
		); 

/******************* CELL 506 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell506 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[445]),
			.N(gen[446]),
			.NE(gen[447]),

			.O(gen[505]),
			.E(gen[507]),

			.SO(gen[565]),
			.S(gen[566]),
			.SE(gen[567]),

			.SELF(gen[506]),
			.cell_state(gen[506])
		); 

/******************* CELL 507 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell507 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[446]),
			.N(gen[447]),
			.NE(gen[448]),

			.O(gen[506]),
			.E(gen[508]),

			.SO(gen[566]),
			.S(gen[567]),
			.SE(gen[568]),

			.SELF(gen[507]),
			.cell_state(gen[507])
		); 

/******************* CELL 508 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell508 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[447]),
			.N(gen[448]),
			.NE(gen[449]),

			.O(gen[507]),
			.E(gen[509]),

			.SO(gen[567]),
			.S(gen[568]),
			.SE(gen[569]),

			.SELF(gen[508]),
			.cell_state(gen[508])
		); 

/******************* CELL 509 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell509 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[448]),
			.N(gen[449]),
			.NE(gen[450]),

			.O(gen[508]),
			.E(gen[510]),

			.SO(gen[568]),
			.S(gen[569]),
			.SE(gen[570]),

			.SELF(gen[509]),
			.cell_state(gen[509])
		); 

/******************* CELL 510 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell510 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[449]),
			.N(gen[450]),
			.NE(gen[451]),

			.O(gen[509]),
			.E(gen[511]),

			.SO(gen[569]),
			.S(gen[570]),
			.SE(gen[571]),

			.SELF(gen[510]),
			.cell_state(gen[510])
		); 

/******************* CELL 511 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell511 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[450]),
			.N(gen[451]),
			.NE(gen[452]),

			.O(gen[510]),
			.E(gen[512]),

			.SO(gen[570]),
			.S(gen[571]),
			.SE(gen[572]),

			.SELF(gen[511]),
			.cell_state(gen[511])
		); 

/******************* CELL 512 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell512 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[451]),
			.N(gen[452]),
			.NE(gen[453]),

			.O(gen[511]),
			.E(gen[513]),

			.SO(gen[571]),
			.S(gen[572]),
			.SE(gen[573]),

			.SELF(gen[512]),
			.cell_state(gen[512])
		); 

/******************* CELL 513 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell513 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[452]),
			.N(gen[453]),
			.NE(gen[454]),

			.O(gen[512]),
			.E(gen[514]),

			.SO(gen[572]),
			.S(gen[573]),
			.SE(gen[574]),

			.SELF(gen[513]),
			.cell_state(gen[513])
		); 

/******************* CELL 514 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell514 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[453]),
			.N(gen[454]),
			.NE(gen[455]),

			.O(gen[513]),
			.E(gen[515]),

			.SO(gen[573]),
			.S(gen[574]),
			.SE(gen[575]),

			.SELF(gen[514]),
			.cell_state(gen[514])
		); 

/******************* CELL 515 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell515 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[454]),
			.N(gen[455]),
			.NE(gen[456]),

			.O(gen[514]),
			.E(gen[516]),

			.SO(gen[574]),
			.S(gen[575]),
			.SE(gen[576]),

			.SELF(gen[515]),
			.cell_state(gen[515])
		); 

/******************* CELL 516 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell516 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[455]),
			.N(gen[456]),
			.NE(gen[457]),

			.O(gen[515]),
			.E(gen[517]),

			.SO(gen[575]),
			.S(gen[576]),
			.SE(gen[577]),

			.SELF(gen[516]),
			.cell_state(gen[516])
		); 

/******************* CELL 517 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell517 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[456]),
			.N(gen[457]),
			.NE(gen[458]),

			.O(gen[516]),
			.E(gen[518]),

			.SO(gen[576]),
			.S(gen[577]),
			.SE(gen[578]),

			.SELF(gen[517]),
			.cell_state(gen[517])
		); 

/******************* CELL 518 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell518 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[457]),
			.N(gen[458]),
			.NE(gen[459]),

			.O(gen[517]),
			.E(gen[519]),

			.SO(gen[577]),
			.S(gen[578]),
			.SE(gen[579]),

			.SELF(gen[518]),
			.cell_state(gen[518])
		); 

/******************* CELL 519 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell519 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[458]),
			.N(gen[459]),
			.NE(gen[460]),

			.O(gen[518]),
			.E(gen[520]),

			.SO(gen[578]),
			.S(gen[579]),
			.SE(gen[580]),

			.SELF(gen[519]),
			.cell_state(gen[519])
		); 

/******************* CELL 520 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell520 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[459]),
			.N(gen[460]),
			.NE(gen[461]),

			.O(gen[519]),
			.E(gen[521]),

			.SO(gen[579]),
			.S(gen[580]),
			.SE(gen[581]),

			.SELF(gen[520]),
			.cell_state(gen[520])
		); 

/******************* CELL 521 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell521 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[460]),
			.N(gen[461]),
			.NE(gen[462]),

			.O(gen[520]),
			.E(gen[522]),

			.SO(gen[580]),
			.S(gen[581]),
			.SE(gen[582]),

			.SELF(gen[521]),
			.cell_state(gen[521])
		); 

/******************* CELL 522 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell522 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[461]),
			.N(gen[462]),
			.NE(gen[463]),

			.O(gen[521]),
			.E(gen[523]),

			.SO(gen[581]),
			.S(gen[582]),
			.SE(gen[583]),

			.SELF(gen[522]),
			.cell_state(gen[522])
		); 

/******************* CELL 523 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell523 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[462]),
			.N(gen[463]),
			.NE(gen[464]),

			.O(gen[522]),
			.E(gen[524]),

			.SO(gen[582]),
			.S(gen[583]),
			.SE(gen[584]),

			.SELF(gen[523]),
			.cell_state(gen[523])
		); 

/******************* CELL 524 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell524 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[463]),
			.N(gen[464]),
			.NE(gen[465]),

			.O(gen[523]),
			.E(gen[525]),

			.SO(gen[583]),
			.S(gen[584]),
			.SE(gen[585]),

			.SELF(gen[524]),
			.cell_state(gen[524])
		); 

/******************* CELL 525 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell525 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[464]),
			.N(gen[465]),
			.NE(gen[466]),

			.O(gen[524]),
			.E(gen[526]),

			.SO(gen[584]),
			.S(gen[585]),
			.SE(gen[586]),

			.SELF(gen[525]),
			.cell_state(gen[525])
		); 

/******************* CELL 526 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell526 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[465]),
			.N(gen[466]),
			.NE(gen[467]),

			.O(gen[525]),
			.E(gen[527]),

			.SO(gen[585]),
			.S(gen[586]),
			.SE(gen[587]),

			.SELF(gen[526]),
			.cell_state(gen[526])
		); 

/******************* CELL 527 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell527 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[466]),
			.N(gen[467]),
			.NE(gen[468]),

			.O(gen[526]),
			.E(gen[528]),

			.SO(gen[586]),
			.S(gen[587]),
			.SE(gen[588]),

			.SELF(gen[527]),
			.cell_state(gen[527])
		); 

/******************* CELL 528 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell528 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[467]),
			.N(gen[468]),
			.NE(gen[469]),

			.O(gen[527]),
			.E(gen[529]),

			.SO(gen[587]),
			.S(gen[588]),
			.SE(gen[589]),

			.SELF(gen[528]),
			.cell_state(gen[528])
		); 

/******************* CELL 529 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell529 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[468]),
			.N(gen[469]),
			.NE(gen[470]),

			.O(gen[528]),
			.E(gen[530]),

			.SO(gen[588]),
			.S(gen[589]),
			.SE(gen[590]),

			.SELF(gen[529]),
			.cell_state(gen[529])
		); 

/******************* CELL 530 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell530 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[469]),
			.N(gen[470]),
			.NE(gen[471]),

			.O(gen[529]),
			.E(gen[531]),

			.SO(gen[589]),
			.S(gen[590]),
			.SE(gen[591]),

			.SELF(gen[530]),
			.cell_state(gen[530])
		); 

/******************* CELL 531 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell531 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[470]),
			.N(gen[471]),
			.NE(gen[472]),

			.O(gen[530]),
			.E(gen[532]),

			.SO(gen[590]),
			.S(gen[591]),
			.SE(gen[592]),

			.SELF(gen[531]),
			.cell_state(gen[531])
		); 

/******************* CELL 532 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell532 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[471]),
			.N(gen[472]),
			.NE(gen[473]),

			.O(gen[531]),
			.E(gen[533]),

			.SO(gen[591]),
			.S(gen[592]),
			.SE(gen[593]),

			.SELF(gen[532]),
			.cell_state(gen[532])
		); 

/******************* CELL 533 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell533 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[472]),
			.N(gen[473]),
			.NE(gen[474]),

			.O(gen[532]),
			.E(gen[534]),

			.SO(gen[592]),
			.S(gen[593]),
			.SE(gen[594]),

			.SELF(gen[533]),
			.cell_state(gen[533])
		); 

/******************* CELL 534 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell534 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[473]),
			.N(gen[474]),
			.NE(gen[475]),

			.O(gen[533]),
			.E(gen[535]),

			.SO(gen[593]),
			.S(gen[594]),
			.SE(gen[595]),

			.SELF(gen[534]),
			.cell_state(gen[534])
		); 

/******************* CELL 535 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell535 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[474]),
			.N(gen[475]),
			.NE(gen[476]),

			.O(gen[534]),
			.E(gen[536]),

			.SO(gen[594]),
			.S(gen[595]),
			.SE(gen[596]),

			.SELF(gen[535]),
			.cell_state(gen[535])
		); 

/******************* CELL 536 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell536 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[475]),
			.N(gen[476]),
			.NE(gen[477]),

			.O(gen[535]),
			.E(gen[537]),

			.SO(gen[595]),
			.S(gen[596]),
			.SE(gen[597]),

			.SELF(gen[536]),
			.cell_state(gen[536])
		); 

/******************* CELL 537 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell537 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[476]),
			.N(gen[477]),
			.NE(gen[478]),

			.O(gen[536]),
			.E(gen[538]),

			.SO(gen[596]),
			.S(gen[597]),
			.SE(gen[598]),

			.SELF(gen[537]),
			.cell_state(gen[537])
		); 

/******************* CELL 538 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell538 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[477]),
			.N(gen[478]),
			.NE(gen[479]),

			.O(gen[537]),
			.E(gen[539]),

			.SO(gen[597]),
			.S(gen[598]),
			.SE(gen[599]),

			.SELF(gen[538]),
			.cell_state(gen[538])
		); 

/******************* CELL 539 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell539 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[478]),
			.N(gen[479]),
			.NE(gen[478]),

			.O(gen[538]),
			.E(gen[538]),

			.SO(gen[598]),
			.S(gen[599]),
			.SE(gen[598]),

			.SELF(gen[539]),
			.cell_state(gen[539])
		); 

/******************* CELL 540 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell540 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[481]),
			.N(gen[480]),
			.NE(gen[481]),

			.O(gen[541]),
			.E(gen[541]),

			.SO(gen[601]),
			.S(gen[600]),
			.SE(gen[601]),

			.SELF(gen[540]),
			.cell_state(gen[540])
		); 

/******************* CELL 541 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell541 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[480]),
			.N(gen[481]),
			.NE(gen[482]),

			.O(gen[540]),
			.E(gen[542]),

			.SO(gen[600]),
			.S(gen[601]),
			.SE(gen[602]),

			.SELF(gen[541]),
			.cell_state(gen[541])
		); 

/******************* CELL 542 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell542 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[481]),
			.N(gen[482]),
			.NE(gen[483]),

			.O(gen[541]),
			.E(gen[543]),

			.SO(gen[601]),
			.S(gen[602]),
			.SE(gen[603]),

			.SELF(gen[542]),
			.cell_state(gen[542])
		); 

/******************* CELL 543 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell543 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[482]),
			.N(gen[483]),
			.NE(gen[484]),

			.O(gen[542]),
			.E(gen[544]),

			.SO(gen[602]),
			.S(gen[603]),
			.SE(gen[604]),

			.SELF(gen[543]),
			.cell_state(gen[543])
		); 

/******************* CELL 544 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell544 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[483]),
			.N(gen[484]),
			.NE(gen[485]),

			.O(gen[543]),
			.E(gen[545]),

			.SO(gen[603]),
			.S(gen[604]),
			.SE(gen[605]),

			.SELF(gen[544]),
			.cell_state(gen[544])
		); 

/******************* CELL 545 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell545 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[484]),
			.N(gen[485]),
			.NE(gen[486]),

			.O(gen[544]),
			.E(gen[546]),

			.SO(gen[604]),
			.S(gen[605]),
			.SE(gen[606]),

			.SELF(gen[545]),
			.cell_state(gen[545])
		); 

/******************* CELL 546 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell546 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[485]),
			.N(gen[486]),
			.NE(gen[487]),

			.O(gen[545]),
			.E(gen[547]),

			.SO(gen[605]),
			.S(gen[606]),
			.SE(gen[607]),

			.SELF(gen[546]),
			.cell_state(gen[546])
		); 

/******************* CELL 547 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell547 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[486]),
			.N(gen[487]),
			.NE(gen[488]),

			.O(gen[546]),
			.E(gen[548]),

			.SO(gen[606]),
			.S(gen[607]),
			.SE(gen[608]),

			.SELF(gen[547]),
			.cell_state(gen[547])
		); 

/******************* CELL 548 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell548 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[487]),
			.N(gen[488]),
			.NE(gen[489]),

			.O(gen[547]),
			.E(gen[549]),

			.SO(gen[607]),
			.S(gen[608]),
			.SE(gen[609]),

			.SELF(gen[548]),
			.cell_state(gen[548])
		); 

/******************* CELL 549 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell549 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[488]),
			.N(gen[489]),
			.NE(gen[490]),

			.O(gen[548]),
			.E(gen[550]),

			.SO(gen[608]),
			.S(gen[609]),
			.SE(gen[610]),

			.SELF(gen[549]),
			.cell_state(gen[549])
		); 

/******************* CELL 550 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell550 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[489]),
			.N(gen[490]),
			.NE(gen[491]),

			.O(gen[549]),
			.E(gen[551]),

			.SO(gen[609]),
			.S(gen[610]),
			.SE(gen[611]),

			.SELF(gen[550]),
			.cell_state(gen[550])
		); 

/******************* CELL 551 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell551 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[490]),
			.N(gen[491]),
			.NE(gen[492]),

			.O(gen[550]),
			.E(gen[552]),

			.SO(gen[610]),
			.S(gen[611]),
			.SE(gen[612]),

			.SELF(gen[551]),
			.cell_state(gen[551])
		); 

/******************* CELL 552 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell552 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[491]),
			.N(gen[492]),
			.NE(gen[493]),

			.O(gen[551]),
			.E(gen[553]),

			.SO(gen[611]),
			.S(gen[612]),
			.SE(gen[613]),

			.SELF(gen[552]),
			.cell_state(gen[552])
		); 

/******************* CELL 553 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell553 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[492]),
			.N(gen[493]),
			.NE(gen[494]),

			.O(gen[552]),
			.E(gen[554]),

			.SO(gen[612]),
			.S(gen[613]),
			.SE(gen[614]),

			.SELF(gen[553]),
			.cell_state(gen[553])
		); 

/******************* CELL 554 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell554 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[493]),
			.N(gen[494]),
			.NE(gen[495]),

			.O(gen[553]),
			.E(gen[555]),

			.SO(gen[613]),
			.S(gen[614]),
			.SE(gen[615]),

			.SELF(gen[554]),
			.cell_state(gen[554])
		); 

/******************* CELL 555 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell555 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[494]),
			.N(gen[495]),
			.NE(gen[496]),

			.O(gen[554]),
			.E(gen[556]),

			.SO(gen[614]),
			.S(gen[615]),
			.SE(gen[616]),

			.SELF(gen[555]),
			.cell_state(gen[555])
		); 

/******************* CELL 556 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell556 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[495]),
			.N(gen[496]),
			.NE(gen[497]),

			.O(gen[555]),
			.E(gen[557]),

			.SO(gen[615]),
			.S(gen[616]),
			.SE(gen[617]),

			.SELF(gen[556]),
			.cell_state(gen[556])
		); 

/******************* CELL 557 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell557 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[496]),
			.N(gen[497]),
			.NE(gen[498]),

			.O(gen[556]),
			.E(gen[558]),

			.SO(gen[616]),
			.S(gen[617]),
			.SE(gen[618]),

			.SELF(gen[557]),
			.cell_state(gen[557])
		); 

/******************* CELL 558 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell558 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[497]),
			.N(gen[498]),
			.NE(gen[499]),

			.O(gen[557]),
			.E(gen[559]),

			.SO(gen[617]),
			.S(gen[618]),
			.SE(gen[619]),

			.SELF(gen[558]),
			.cell_state(gen[558])
		); 

/******************* CELL 559 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell559 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[498]),
			.N(gen[499]),
			.NE(gen[500]),

			.O(gen[558]),
			.E(gen[560]),

			.SO(gen[618]),
			.S(gen[619]),
			.SE(gen[620]),

			.SELF(gen[559]),
			.cell_state(gen[559])
		); 

/******************* CELL 560 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell560 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[499]),
			.N(gen[500]),
			.NE(gen[501]),

			.O(gen[559]),
			.E(gen[561]),

			.SO(gen[619]),
			.S(gen[620]),
			.SE(gen[621]),

			.SELF(gen[560]),
			.cell_state(gen[560])
		); 

/******************* CELL 561 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell561 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[500]),
			.N(gen[501]),
			.NE(gen[502]),

			.O(gen[560]),
			.E(gen[562]),

			.SO(gen[620]),
			.S(gen[621]),
			.SE(gen[622]),

			.SELF(gen[561]),
			.cell_state(gen[561])
		); 

/******************* CELL 562 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell562 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[501]),
			.N(gen[502]),
			.NE(gen[503]),

			.O(gen[561]),
			.E(gen[563]),

			.SO(gen[621]),
			.S(gen[622]),
			.SE(gen[623]),

			.SELF(gen[562]),
			.cell_state(gen[562])
		); 

/******************* CELL 563 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell563 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[502]),
			.N(gen[503]),
			.NE(gen[504]),

			.O(gen[562]),
			.E(gen[564]),

			.SO(gen[622]),
			.S(gen[623]),
			.SE(gen[624]),

			.SELF(gen[563]),
			.cell_state(gen[563])
		); 

/******************* CELL 564 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell564 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[503]),
			.N(gen[504]),
			.NE(gen[505]),

			.O(gen[563]),
			.E(gen[565]),

			.SO(gen[623]),
			.S(gen[624]),
			.SE(gen[625]),

			.SELF(gen[564]),
			.cell_state(gen[564])
		); 

/******************* CELL 565 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell565 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[504]),
			.N(gen[505]),
			.NE(gen[506]),

			.O(gen[564]),
			.E(gen[566]),

			.SO(gen[624]),
			.S(gen[625]),
			.SE(gen[626]),

			.SELF(gen[565]),
			.cell_state(gen[565])
		); 

/******************* CELL 566 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell566 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[505]),
			.N(gen[506]),
			.NE(gen[507]),

			.O(gen[565]),
			.E(gen[567]),

			.SO(gen[625]),
			.S(gen[626]),
			.SE(gen[627]),

			.SELF(gen[566]),
			.cell_state(gen[566])
		); 

/******************* CELL 567 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell567 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[506]),
			.N(gen[507]),
			.NE(gen[508]),

			.O(gen[566]),
			.E(gen[568]),

			.SO(gen[626]),
			.S(gen[627]),
			.SE(gen[628]),

			.SELF(gen[567]),
			.cell_state(gen[567])
		); 

/******************* CELL 568 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell568 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[507]),
			.N(gen[508]),
			.NE(gen[509]),

			.O(gen[567]),
			.E(gen[569]),

			.SO(gen[627]),
			.S(gen[628]),
			.SE(gen[629]),

			.SELF(gen[568]),
			.cell_state(gen[568])
		); 

/******************* CELL 569 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell569 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[508]),
			.N(gen[509]),
			.NE(gen[510]),

			.O(gen[568]),
			.E(gen[570]),

			.SO(gen[628]),
			.S(gen[629]),
			.SE(gen[630]),

			.SELF(gen[569]),
			.cell_state(gen[569])
		); 

/******************* CELL 570 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell570 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[509]),
			.N(gen[510]),
			.NE(gen[511]),

			.O(gen[569]),
			.E(gen[571]),

			.SO(gen[629]),
			.S(gen[630]),
			.SE(gen[631]),

			.SELF(gen[570]),
			.cell_state(gen[570])
		); 

/******************* CELL 571 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell571 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[510]),
			.N(gen[511]),
			.NE(gen[512]),

			.O(gen[570]),
			.E(gen[572]),

			.SO(gen[630]),
			.S(gen[631]),
			.SE(gen[632]),

			.SELF(gen[571]),
			.cell_state(gen[571])
		); 

/******************* CELL 572 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell572 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[511]),
			.N(gen[512]),
			.NE(gen[513]),

			.O(gen[571]),
			.E(gen[573]),

			.SO(gen[631]),
			.S(gen[632]),
			.SE(gen[633]),

			.SELF(gen[572]),
			.cell_state(gen[572])
		); 

/******************* CELL 573 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell573 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[512]),
			.N(gen[513]),
			.NE(gen[514]),

			.O(gen[572]),
			.E(gen[574]),

			.SO(gen[632]),
			.S(gen[633]),
			.SE(gen[634]),

			.SELF(gen[573]),
			.cell_state(gen[573])
		); 

/******************* CELL 574 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell574 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[513]),
			.N(gen[514]),
			.NE(gen[515]),

			.O(gen[573]),
			.E(gen[575]),

			.SO(gen[633]),
			.S(gen[634]),
			.SE(gen[635]),

			.SELF(gen[574]),
			.cell_state(gen[574])
		); 

/******************* CELL 575 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell575 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[514]),
			.N(gen[515]),
			.NE(gen[516]),

			.O(gen[574]),
			.E(gen[576]),

			.SO(gen[634]),
			.S(gen[635]),
			.SE(gen[636]),

			.SELF(gen[575]),
			.cell_state(gen[575])
		); 

/******************* CELL 576 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell576 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[515]),
			.N(gen[516]),
			.NE(gen[517]),

			.O(gen[575]),
			.E(gen[577]),

			.SO(gen[635]),
			.S(gen[636]),
			.SE(gen[637]),

			.SELF(gen[576]),
			.cell_state(gen[576])
		); 

/******************* CELL 577 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell577 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[516]),
			.N(gen[517]),
			.NE(gen[518]),

			.O(gen[576]),
			.E(gen[578]),

			.SO(gen[636]),
			.S(gen[637]),
			.SE(gen[638]),

			.SELF(gen[577]),
			.cell_state(gen[577])
		); 

/******************* CELL 578 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell578 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[517]),
			.N(gen[518]),
			.NE(gen[519]),

			.O(gen[577]),
			.E(gen[579]),

			.SO(gen[637]),
			.S(gen[638]),
			.SE(gen[639]),

			.SELF(gen[578]),
			.cell_state(gen[578])
		); 

/******************* CELL 579 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell579 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[518]),
			.N(gen[519]),
			.NE(gen[520]),

			.O(gen[578]),
			.E(gen[580]),

			.SO(gen[638]),
			.S(gen[639]),
			.SE(gen[640]),

			.SELF(gen[579]),
			.cell_state(gen[579])
		); 

/******************* CELL 580 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell580 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[519]),
			.N(gen[520]),
			.NE(gen[521]),

			.O(gen[579]),
			.E(gen[581]),

			.SO(gen[639]),
			.S(gen[640]),
			.SE(gen[641]),

			.SELF(gen[580]),
			.cell_state(gen[580])
		); 

/******************* CELL 581 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell581 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[520]),
			.N(gen[521]),
			.NE(gen[522]),

			.O(gen[580]),
			.E(gen[582]),

			.SO(gen[640]),
			.S(gen[641]),
			.SE(gen[642]),

			.SELF(gen[581]),
			.cell_state(gen[581])
		); 

/******************* CELL 582 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell582 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[521]),
			.N(gen[522]),
			.NE(gen[523]),

			.O(gen[581]),
			.E(gen[583]),

			.SO(gen[641]),
			.S(gen[642]),
			.SE(gen[643]),

			.SELF(gen[582]),
			.cell_state(gen[582])
		); 

/******************* CELL 583 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell583 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[522]),
			.N(gen[523]),
			.NE(gen[524]),

			.O(gen[582]),
			.E(gen[584]),

			.SO(gen[642]),
			.S(gen[643]),
			.SE(gen[644]),

			.SELF(gen[583]),
			.cell_state(gen[583])
		); 

/******************* CELL 584 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell584 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[523]),
			.N(gen[524]),
			.NE(gen[525]),

			.O(gen[583]),
			.E(gen[585]),

			.SO(gen[643]),
			.S(gen[644]),
			.SE(gen[645]),

			.SELF(gen[584]),
			.cell_state(gen[584])
		); 

/******************* CELL 585 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell585 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[524]),
			.N(gen[525]),
			.NE(gen[526]),

			.O(gen[584]),
			.E(gen[586]),

			.SO(gen[644]),
			.S(gen[645]),
			.SE(gen[646]),

			.SELF(gen[585]),
			.cell_state(gen[585])
		); 

/******************* CELL 586 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell586 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[525]),
			.N(gen[526]),
			.NE(gen[527]),

			.O(gen[585]),
			.E(gen[587]),

			.SO(gen[645]),
			.S(gen[646]),
			.SE(gen[647]),

			.SELF(gen[586]),
			.cell_state(gen[586])
		); 

/******************* CELL 587 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell587 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[526]),
			.N(gen[527]),
			.NE(gen[528]),

			.O(gen[586]),
			.E(gen[588]),

			.SO(gen[646]),
			.S(gen[647]),
			.SE(gen[648]),

			.SELF(gen[587]),
			.cell_state(gen[587])
		); 

/******************* CELL 588 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell588 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[527]),
			.N(gen[528]),
			.NE(gen[529]),

			.O(gen[587]),
			.E(gen[589]),

			.SO(gen[647]),
			.S(gen[648]),
			.SE(gen[649]),

			.SELF(gen[588]),
			.cell_state(gen[588])
		); 

/******************* CELL 589 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell589 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[528]),
			.N(gen[529]),
			.NE(gen[530]),

			.O(gen[588]),
			.E(gen[590]),

			.SO(gen[648]),
			.S(gen[649]),
			.SE(gen[650]),

			.SELF(gen[589]),
			.cell_state(gen[589])
		); 

/******************* CELL 590 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell590 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[529]),
			.N(gen[530]),
			.NE(gen[531]),

			.O(gen[589]),
			.E(gen[591]),

			.SO(gen[649]),
			.S(gen[650]),
			.SE(gen[651]),

			.SELF(gen[590]),
			.cell_state(gen[590])
		); 

/******************* CELL 591 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell591 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[530]),
			.N(gen[531]),
			.NE(gen[532]),

			.O(gen[590]),
			.E(gen[592]),

			.SO(gen[650]),
			.S(gen[651]),
			.SE(gen[652]),

			.SELF(gen[591]),
			.cell_state(gen[591])
		); 

/******************* CELL 592 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell592 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[531]),
			.N(gen[532]),
			.NE(gen[533]),

			.O(gen[591]),
			.E(gen[593]),

			.SO(gen[651]),
			.S(gen[652]),
			.SE(gen[653]),

			.SELF(gen[592]),
			.cell_state(gen[592])
		); 

/******************* CELL 593 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell593 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[532]),
			.N(gen[533]),
			.NE(gen[534]),

			.O(gen[592]),
			.E(gen[594]),

			.SO(gen[652]),
			.S(gen[653]),
			.SE(gen[654]),

			.SELF(gen[593]),
			.cell_state(gen[593])
		); 

/******************* CELL 594 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell594 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[533]),
			.N(gen[534]),
			.NE(gen[535]),

			.O(gen[593]),
			.E(gen[595]),

			.SO(gen[653]),
			.S(gen[654]),
			.SE(gen[655]),

			.SELF(gen[594]),
			.cell_state(gen[594])
		); 

/******************* CELL 595 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell595 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[534]),
			.N(gen[535]),
			.NE(gen[536]),

			.O(gen[594]),
			.E(gen[596]),

			.SO(gen[654]),
			.S(gen[655]),
			.SE(gen[656]),

			.SELF(gen[595]),
			.cell_state(gen[595])
		); 

/******************* CELL 596 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell596 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[535]),
			.N(gen[536]),
			.NE(gen[537]),

			.O(gen[595]),
			.E(gen[597]),

			.SO(gen[655]),
			.S(gen[656]),
			.SE(gen[657]),

			.SELF(gen[596]),
			.cell_state(gen[596])
		); 

/******************* CELL 597 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell597 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[536]),
			.N(gen[537]),
			.NE(gen[538]),

			.O(gen[596]),
			.E(gen[598]),

			.SO(gen[656]),
			.S(gen[657]),
			.SE(gen[658]),

			.SELF(gen[597]),
			.cell_state(gen[597])
		); 

/******************* CELL 598 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell598 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[537]),
			.N(gen[538]),
			.NE(gen[539]),

			.O(gen[597]),
			.E(gen[599]),

			.SO(gen[657]),
			.S(gen[658]),
			.SE(gen[659]),

			.SELF(gen[598]),
			.cell_state(gen[598])
		); 

/******************* CELL 599 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell599 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[538]),
			.N(gen[539]),
			.NE(gen[538]),

			.O(gen[598]),
			.E(gen[598]),

			.SO(gen[658]),
			.S(gen[659]),
			.SE(gen[658]),

			.SELF(gen[599]),
			.cell_state(gen[599])
		); 

/******************* CELL 600 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell600 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[541]),
			.N(gen[540]),
			.NE(gen[541]),

			.O(gen[601]),
			.E(gen[601]),

			.SO(gen[661]),
			.S(gen[660]),
			.SE(gen[661]),

			.SELF(gen[600]),
			.cell_state(gen[600])
		); 

/******************* CELL 601 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell601 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[540]),
			.N(gen[541]),
			.NE(gen[542]),

			.O(gen[600]),
			.E(gen[602]),

			.SO(gen[660]),
			.S(gen[661]),
			.SE(gen[662]),

			.SELF(gen[601]),
			.cell_state(gen[601])
		); 

/******************* CELL 602 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell602 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[541]),
			.N(gen[542]),
			.NE(gen[543]),

			.O(gen[601]),
			.E(gen[603]),

			.SO(gen[661]),
			.S(gen[662]),
			.SE(gen[663]),

			.SELF(gen[602]),
			.cell_state(gen[602])
		); 

/******************* CELL 603 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell603 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[542]),
			.N(gen[543]),
			.NE(gen[544]),

			.O(gen[602]),
			.E(gen[604]),

			.SO(gen[662]),
			.S(gen[663]),
			.SE(gen[664]),

			.SELF(gen[603]),
			.cell_state(gen[603])
		); 

/******************* CELL 604 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell604 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[543]),
			.N(gen[544]),
			.NE(gen[545]),

			.O(gen[603]),
			.E(gen[605]),

			.SO(gen[663]),
			.S(gen[664]),
			.SE(gen[665]),

			.SELF(gen[604]),
			.cell_state(gen[604])
		); 

/******************* CELL 605 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell605 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[544]),
			.N(gen[545]),
			.NE(gen[546]),

			.O(gen[604]),
			.E(gen[606]),

			.SO(gen[664]),
			.S(gen[665]),
			.SE(gen[666]),

			.SELF(gen[605]),
			.cell_state(gen[605])
		); 

/******************* CELL 606 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell606 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[545]),
			.N(gen[546]),
			.NE(gen[547]),

			.O(gen[605]),
			.E(gen[607]),

			.SO(gen[665]),
			.S(gen[666]),
			.SE(gen[667]),

			.SELF(gen[606]),
			.cell_state(gen[606])
		); 

/******************* CELL 607 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell607 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[546]),
			.N(gen[547]),
			.NE(gen[548]),

			.O(gen[606]),
			.E(gen[608]),

			.SO(gen[666]),
			.S(gen[667]),
			.SE(gen[668]),

			.SELF(gen[607]),
			.cell_state(gen[607])
		); 

/******************* CELL 608 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell608 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[547]),
			.N(gen[548]),
			.NE(gen[549]),

			.O(gen[607]),
			.E(gen[609]),

			.SO(gen[667]),
			.S(gen[668]),
			.SE(gen[669]),

			.SELF(gen[608]),
			.cell_state(gen[608])
		); 

/******************* CELL 609 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell609 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[548]),
			.N(gen[549]),
			.NE(gen[550]),

			.O(gen[608]),
			.E(gen[610]),

			.SO(gen[668]),
			.S(gen[669]),
			.SE(gen[670]),

			.SELF(gen[609]),
			.cell_state(gen[609])
		); 

/******************* CELL 610 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell610 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[549]),
			.N(gen[550]),
			.NE(gen[551]),

			.O(gen[609]),
			.E(gen[611]),

			.SO(gen[669]),
			.S(gen[670]),
			.SE(gen[671]),

			.SELF(gen[610]),
			.cell_state(gen[610])
		); 

/******************* CELL 611 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell611 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[550]),
			.N(gen[551]),
			.NE(gen[552]),

			.O(gen[610]),
			.E(gen[612]),

			.SO(gen[670]),
			.S(gen[671]),
			.SE(gen[672]),

			.SELF(gen[611]),
			.cell_state(gen[611])
		); 

/******************* CELL 612 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell612 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[551]),
			.N(gen[552]),
			.NE(gen[553]),

			.O(gen[611]),
			.E(gen[613]),

			.SO(gen[671]),
			.S(gen[672]),
			.SE(gen[673]),

			.SELF(gen[612]),
			.cell_state(gen[612])
		); 

/******************* CELL 613 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell613 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[552]),
			.N(gen[553]),
			.NE(gen[554]),

			.O(gen[612]),
			.E(gen[614]),

			.SO(gen[672]),
			.S(gen[673]),
			.SE(gen[674]),

			.SELF(gen[613]),
			.cell_state(gen[613])
		); 

/******************* CELL 614 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell614 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[553]),
			.N(gen[554]),
			.NE(gen[555]),

			.O(gen[613]),
			.E(gen[615]),

			.SO(gen[673]),
			.S(gen[674]),
			.SE(gen[675]),

			.SELF(gen[614]),
			.cell_state(gen[614])
		); 

/******************* CELL 615 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell615 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[554]),
			.N(gen[555]),
			.NE(gen[556]),

			.O(gen[614]),
			.E(gen[616]),

			.SO(gen[674]),
			.S(gen[675]),
			.SE(gen[676]),

			.SELF(gen[615]),
			.cell_state(gen[615])
		); 

/******************* CELL 616 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell616 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[555]),
			.N(gen[556]),
			.NE(gen[557]),

			.O(gen[615]),
			.E(gen[617]),

			.SO(gen[675]),
			.S(gen[676]),
			.SE(gen[677]),

			.SELF(gen[616]),
			.cell_state(gen[616])
		); 

/******************* CELL 617 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell617 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[556]),
			.N(gen[557]),
			.NE(gen[558]),

			.O(gen[616]),
			.E(gen[618]),

			.SO(gen[676]),
			.S(gen[677]),
			.SE(gen[678]),

			.SELF(gen[617]),
			.cell_state(gen[617])
		); 

/******************* CELL 618 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell618 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[557]),
			.N(gen[558]),
			.NE(gen[559]),

			.O(gen[617]),
			.E(gen[619]),

			.SO(gen[677]),
			.S(gen[678]),
			.SE(gen[679]),

			.SELF(gen[618]),
			.cell_state(gen[618])
		); 

/******************* CELL 619 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell619 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[558]),
			.N(gen[559]),
			.NE(gen[560]),

			.O(gen[618]),
			.E(gen[620]),

			.SO(gen[678]),
			.S(gen[679]),
			.SE(gen[680]),

			.SELF(gen[619]),
			.cell_state(gen[619])
		); 

/******************* CELL 620 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell620 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[559]),
			.N(gen[560]),
			.NE(gen[561]),

			.O(gen[619]),
			.E(gen[621]),

			.SO(gen[679]),
			.S(gen[680]),
			.SE(gen[681]),

			.SELF(gen[620]),
			.cell_state(gen[620])
		); 

/******************* CELL 621 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell621 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[560]),
			.N(gen[561]),
			.NE(gen[562]),

			.O(gen[620]),
			.E(gen[622]),

			.SO(gen[680]),
			.S(gen[681]),
			.SE(gen[682]),

			.SELF(gen[621]),
			.cell_state(gen[621])
		); 

/******************* CELL 622 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell622 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[561]),
			.N(gen[562]),
			.NE(gen[563]),

			.O(gen[621]),
			.E(gen[623]),

			.SO(gen[681]),
			.S(gen[682]),
			.SE(gen[683]),

			.SELF(gen[622]),
			.cell_state(gen[622])
		); 

/******************* CELL 623 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell623 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[562]),
			.N(gen[563]),
			.NE(gen[564]),

			.O(gen[622]),
			.E(gen[624]),

			.SO(gen[682]),
			.S(gen[683]),
			.SE(gen[684]),

			.SELF(gen[623]),
			.cell_state(gen[623])
		); 

/******************* CELL 624 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell624 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[563]),
			.N(gen[564]),
			.NE(gen[565]),

			.O(gen[623]),
			.E(gen[625]),

			.SO(gen[683]),
			.S(gen[684]),
			.SE(gen[685]),

			.SELF(gen[624]),
			.cell_state(gen[624])
		); 

/******************* CELL 625 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell625 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[564]),
			.N(gen[565]),
			.NE(gen[566]),

			.O(gen[624]),
			.E(gen[626]),

			.SO(gen[684]),
			.S(gen[685]),
			.SE(gen[686]),

			.SELF(gen[625]),
			.cell_state(gen[625])
		); 

/******************* CELL 626 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell626 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[565]),
			.N(gen[566]),
			.NE(gen[567]),

			.O(gen[625]),
			.E(gen[627]),

			.SO(gen[685]),
			.S(gen[686]),
			.SE(gen[687]),

			.SELF(gen[626]),
			.cell_state(gen[626])
		); 

/******************* CELL 627 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell627 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[566]),
			.N(gen[567]),
			.NE(gen[568]),

			.O(gen[626]),
			.E(gen[628]),

			.SO(gen[686]),
			.S(gen[687]),
			.SE(gen[688]),

			.SELF(gen[627]),
			.cell_state(gen[627])
		); 

/******************* CELL 628 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell628 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[567]),
			.N(gen[568]),
			.NE(gen[569]),

			.O(gen[627]),
			.E(gen[629]),

			.SO(gen[687]),
			.S(gen[688]),
			.SE(gen[689]),

			.SELF(gen[628]),
			.cell_state(gen[628])
		); 

/******************* CELL 629 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell629 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[568]),
			.N(gen[569]),
			.NE(gen[570]),

			.O(gen[628]),
			.E(gen[630]),

			.SO(gen[688]),
			.S(gen[689]),
			.SE(gen[690]),

			.SELF(gen[629]),
			.cell_state(gen[629])
		); 

/******************* CELL 630 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell630 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[569]),
			.N(gen[570]),
			.NE(gen[571]),

			.O(gen[629]),
			.E(gen[631]),

			.SO(gen[689]),
			.S(gen[690]),
			.SE(gen[691]),

			.SELF(gen[630]),
			.cell_state(gen[630])
		); 

/******************* CELL 631 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell631 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[570]),
			.N(gen[571]),
			.NE(gen[572]),

			.O(gen[630]),
			.E(gen[632]),

			.SO(gen[690]),
			.S(gen[691]),
			.SE(gen[692]),

			.SELF(gen[631]),
			.cell_state(gen[631])
		); 

/******************* CELL 632 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell632 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[571]),
			.N(gen[572]),
			.NE(gen[573]),

			.O(gen[631]),
			.E(gen[633]),

			.SO(gen[691]),
			.S(gen[692]),
			.SE(gen[693]),

			.SELF(gen[632]),
			.cell_state(gen[632])
		); 

/******************* CELL 633 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell633 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[572]),
			.N(gen[573]),
			.NE(gen[574]),

			.O(gen[632]),
			.E(gen[634]),

			.SO(gen[692]),
			.S(gen[693]),
			.SE(gen[694]),

			.SELF(gen[633]),
			.cell_state(gen[633])
		); 

/******************* CELL 634 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell634 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[573]),
			.N(gen[574]),
			.NE(gen[575]),

			.O(gen[633]),
			.E(gen[635]),

			.SO(gen[693]),
			.S(gen[694]),
			.SE(gen[695]),

			.SELF(gen[634]),
			.cell_state(gen[634])
		); 

/******************* CELL 635 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell635 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[574]),
			.N(gen[575]),
			.NE(gen[576]),

			.O(gen[634]),
			.E(gen[636]),

			.SO(gen[694]),
			.S(gen[695]),
			.SE(gen[696]),

			.SELF(gen[635]),
			.cell_state(gen[635])
		); 

/******************* CELL 636 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell636 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[575]),
			.N(gen[576]),
			.NE(gen[577]),

			.O(gen[635]),
			.E(gen[637]),

			.SO(gen[695]),
			.S(gen[696]),
			.SE(gen[697]),

			.SELF(gen[636]),
			.cell_state(gen[636])
		); 

/******************* CELL 637 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell637 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[576]),
			.N(gen[577]),
			.NE(gen[578]),

			.O(gen[636]),
			.E(gen[638]),

			.SO(gen[696]),
			.S(gen[697]),
			.SE(gen[698]),

			.SELF(gen[637]),
			.cell_state(gen[637])
		); 

/******************* CELL 638 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell638 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[577]),
			.N(gen[578]),
			.NE(gen[579]),

			.O(gen[637]),
			.E(gen[639]),

			.SO(gen[697]),
			.S(gen[698]),
			.SE(gen[699]),

			.SELF(gen[638]),
			.cell_state(gen[638])
		); 

/******************* CELL 639 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell639 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[578]),
			.N(gen[579]),
			.NE(gen[580]),

			.O(gen[638]),
			.E(gen[640]),

			.SO(gen[698]),
			.S(gen[699]),
			.SE(gen[700]),

			.SELF(gen[639]),
			.cell_state(gen[639])
		); 

/******************* CELL 640 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell640 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[579]),
			.N(gen[580]),
			.NE(gen[581]),

			.O(gen[639]),
			.E(gen[641]),

			.SO(gen[699]),
			.S(gen[700]),
			.SE(gen[701]),

			.SELF(gen[640]),
			.cell_state(gen[640])
		); 

/******************* CELL 641 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell641 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[580]),
			.N(gen[581]),
			.NE(gen[582]),

			.O(gen[640]),
			.E(gen[642]),

			.SO(gen[700]),
			.S(gen[701]),
			.SE(gen[702]),

			.SELF(gen[641]),
			.cell_state(gen[641])
		); 

/******************* CELL 642 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell642 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[581]),
			.N(gen[582]),
			.NE(gen[583]),

			.O(gen[641]),
			.E(gen[643]),

			.SO(gen[701]),
			.S(gen[702]),
			.SE(gen[703]),

			.SELF(gen[642]),
			.cell_state(gen[642])
		); 

/******************* CELL 643 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell643 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[582]),
			.N(gen[583]),
			.NE(gen[584]),

			.O(gen[642]),
			.E(gen[644]),

			.SO(gen[702]),
			.S(gen[703]),
			.SE(gen[704]),

			.SELF(gen[643]),
			.cell_state(gen[643])
		); 

/******************* CELL 644 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell644 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[583]),
			.N(gen[584]),
			.NE(gen[585]),

			.O(gen[643]),
			.E(gen[645]),

			.SO(gen[703]),
			.S(gen[704]),
			.SE(gen[705]),

			.SELF(gen[644]),
			.cell_state(gen[644])
		); 

/******************* CELL 645 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell645 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[584]),
			.N(gen[585]),
			.NE(gen[586]),

			.O(gen[644]),
			.E(gen[646]),

			.SO(gen[704]),
			.S(gen[705]),
			.SE(gen[706]),

			.SELF(gen[645]),
			.cell_state(gen[645])
		); 

/******************* CELL 646 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell646 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[585]),
			.N(gen[586]),
			.NE(gen[587]),

			.O(gen[645]),
			.E(gen[647]),

			.SO(gen[705]),
			.S(gen[706]),
			.SE(gen[707]),

			.SELF(gen[646]),
			.cell_state(gen[646])
		); 

/******************* CELL 647 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell647 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[586]),
			.N(gen[587]),
			.NE(gen[588]),

			.O(gen[646]),
			.E(gen[648]),

			.SO(gen[706]),
			.S(gen[707]),
			.SE(gen[708]),

			.SELF(gen[647]),
			.cell_state(gen[647])
		); 

/******************* CELL 648 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell648 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[587]),
			.N(gen[588]),
			.NE(gen[589]),

			.O(gen[647]),
			.E(gen[649]),

			.SO(gen[707]),
			.S(gen[708]),
			.SE(gen[709]),

			.SELF(gen[648]),
			.cell_state(gen[648])
		); 

/******************* CELL 649 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell649 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[588]),
			.N(gen[589]),
			.NE(gen[590]),

			.O(gen[648]),
			.E(gen[650]),

			.SO(gen[708]),
			.S(gen[709]),
			.SE(gen[710]),

			.SELF(gen[649]),
			.cell_state(gen[649])
		); 

/******************* CELL 650 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell650 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[589]),
			.N(gen[590]),
			.NE(gen[591]),

			.O(gen[649]),
			.E(gen[651]),

			.SO(gen[709]),
			.S(gen[710]),
			.SE(gen[711]),

			.SELF(gen[650]),
			.cell_state(gen[650])
		); 

/******************* CELL 651 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell651 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[590]),
			.N(gen[591]),
			.NE(gen[592]),

			.O(gen[650]),
			.E(gen[652]),

			.SO(gen[710]),
			.S(gen[711]),
			.SE(gen[712]),

			.SELF(gen[651]),
			.cell_state(gen[651])
		); 

/******************* CELL 652 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell652 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[591]),
			.N(gen[592]),
			.NE(gen[593]),

			.O(gen[651]),
			.E(gen[653]),

			.SO(gen[711]),
			.S(gen[712]),
			.SE(gen[713]),

			.SELF(gen[652]),
			.cell_state(gen[652])
		); 

/******************* CELL 653 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell653 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[592]),
			.N(gen[593]),
			.NE(gen[594]),

			.O(gen[652]),
			.E(gen[654]),

			.SO(gen[712]),
			.S(gen[713]),
			.SE(gen[714]),

			.SELF(gen[653]),
			.cell_state(gen[653])
		); 

/******************* CELL 654 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell654 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[593]),
			.N(gen[594]),
			.NE(gen[595]),

			.O(gen[653]),
			.E(gen[655]),

			.SO(gen[713]),
			.S(gen[714]),
			.SE(gen[715]),

			.SELF(gen[654]),
			.cell_state(gen[654])
		); 

/******************* CELL 655 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell655 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[594]),
			.N(gen[595]),
			.NE(gen[596]),

			.O(gen[654]),
			.E(gen[656]),

			.SO(gen[714]),
			.S(gen[715]),
			.SE(gen[716]),

			.SELF(gen[655]),
			.cell_state(gen[655])
		); 

/******************* CELL 656 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell656 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[595]),
			.N(gen[596]),
			.NE(gen[597]),

			.O(gen[655]),
			.E(gen[657]),

			.SO(gen[715]),
			.S(gen[716]),
			.SE(gen[717]),

			.SELF(gen[656]),
			.cell_state(gen[656])
		); 

/******************* CELL 657 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell657 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[596]),
			.N(gen[597]),
			.NE(gen[598]),

			.O(gen[656]),
			.E(gen[658]),

			.SO(gen[716]),
			.S(gen[717]),
			.SE(gen[718]),

			.SELF(gen[657]),
			.cell_state(gen[657])
		); 

/******************* CELL 658 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell658 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[597]),
			.N(gen[598]),
			.NE(gen[599]),

			.O(gen[657]),
			.E(gen[659]),

			.SO(gen[717]),
			.S(gen[718]),
			.SE(gen[719]),

			.SELF(gen[658]),
			.cell_state(gen[658])
		); 

/******************* CELL 659 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell659 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[598]),
			.N(gen[599]),
			.NE(gen[598]),

			.O(gen[658]),
			.E(gen[658]),

			.SO(gen[718]),
			.S(gen[719]),
			.SE(gen[718]),

			.SELF(gen[659]),
			.cell_state(gen[659])
		); 

/******************* CELL 660 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell660 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[601]),
			.N(gen[600]),
			.NE(gen[601]),

			.O(gen[661]),
			.E(gen[661]),

			.SO(gen[721]),
			.S(gen[720]),
			.SE(gen[721]),

			.SELF(gen[660]),
			.cell_state(gen[660])
		); 

/******************* CELL 661 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell661 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[600]),
			.N(gen[601]),
			.NE(gen[602]),

			.O(gen[660]),
			.E(gen[662]),

			.SO(gen[720]),
			.S(gen[721]),
			.SE(gen[722]),

			.SELF(gen[661]),
			.cell_state(gen[661])
		); 

/******************* CELL 662 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell662 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[601]),
			.N(gen[602]),
			.NE(gen[603]),

			.O(gen[661]),
			.E(gen[663]),

			.SO(gen[721]),
			.S(gen[722]),
			.SE(gen[723]),

			.SELF(gen[662]),
			.cell_state(gen[662])
		); 

/******************* CELL 663 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell663 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[602]),
			.N(gen[603]),
			.NE(gen[604]),

			.O(gen[662]),
			.E(gen[664]),

			.SO(gen[722]),
			.S(gen[723]),
			.SE(gen[724]),

			.SELF(gen[663]),
			.cell_state(gen[663])
		); 

/******************* CELL 664 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell664 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[603]),
			.N(gen[604]),
			.NE(gen[605]),

			.O(gen[663]),
			.E(gen[665]),

			.SO(gen[723]),
			.S(gen[724]),
			.SE(gen[725]),

			.SELF(gen[664]),
			.cell_state(gen[664])
		); 

/******************* CELL 665 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell665 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[604]),
			.N(gen[605]),
			.NE(gen[606]),

			.O(gen[664]),
			.E(gen[666]),

			.SO(gen[724]),
			.S(gen[725]),
			.SE(gen[726]),

			.SELF(gen[665]),
			.cell_state(gen[665])
		); 

/******************* CELL 666 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell666 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[605]),
			.N(gen[606]),
			.NE(gen[607]),

			.O(gen[665]),
			.E(gen[667]),

			.SO(gen[725]),
			.S(gen[726]),
			.SE(gen[727]),

			.SELF(gen[666]),
			.cell_state(gen[666])
		); 

/******************* CELL 667 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell667 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[606]),
			.N(gen[607]),
			.NE(gen[608]),

			.O(gen[666]),
			.E(gen[668]),

			.SO(gen[726]),
			.S(gen[727]),
			.SE(gen[728]),

			.SELF(gen[667]),
			.cell_state(gen[667])
		); 

/******************* CELL 668 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell668 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[607]),
			.N(gen[608]),
			.NE(gen[609]),

			.O(gen[667]),
			.E(gen[669]),

			.SO(gen[727]),
			.S(gen[728]),
			.SE(gen[729]),

			.SELF(gen[668]),
			.cell_state(gen[668])
		); 

/******************* CELL 669 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell669 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[608]),
			.N(gen[609]),
			.NE(gen[610]),

			.O(gen[668]),
			.E(gen[670]),

			.SO(gen[728]),
			.S(gen[729]),
			.SE(gen[730]),

			.SELF(gen[669]),
			.cell_state(gen[669])
		); 

/******************* CELL 670 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell670 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[609]),
			.N(gen[610]),
			.NE(gen[611]),

			.O(gen[669]),
			.E(gen[671]),

			.SO(gen[729]),
			.S(gen[730]),
			.SE(gen[731]),

			.SELF(gen[670]),
			.cell_state(gen[670])
		); 

/******************* CELL 671 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell671 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[610]),
			.N(gen[611]),
			.NE(gen[612]),

			.O(gen[670]),
			.E(gen[672]),

			.SO(gen[730]),
			.S(gen[731]),
			.SE(gen[732]),

			.SELF(gen[671]),
			.cell_state(gen[671])
		); 

/******************* CELL 672 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell672 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[611]),
			.N(gen[612]),
			.NE(gen[613]),

			.O(gen[671]),
			.E(gen[673]),

			.SO(gen[731]),
			.S(gen[732]),
			.SE(gen[733]),

			.SELF(gen[672]),
			.cell_state(gen[672])
		); 

/******************* CELL 673 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell673 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[612]),
			.N(gen[613]),
			.NE(gen[614]),

			.O(gen[672]),
			.E(gen[674]),

			.SO(gen[732]),
			.S(gen[733]),
			.SE(gen[734]),

			.SELF(gen[673]),
			.cell_state(gen[673])
		); 

/******************* CELL 674 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell674 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[613]),
			.N(gen[614]),
			.NE(gen[615]),

			.O(gen[673]),
			.E(gen[675]),

			.SO(gen[733]),
			.S(gen[734]),
			.SE(gen[735]),

			.SELF(gen[674]),
			.cell_state(gen[674])
		); 

/******************* CELL 675 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell675 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[614]),
			.N(gen[615]),
			.NE(gen[616]),

			.O(gen[674]),
			.E(gen[676]),

			.SO(gen[734]),
			.S(gen[735]),
			.SE(gen[736]),

			.SELF(gen[675]),
			.cell_state(gen[675])
		); 

/******************* CELL 676 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell676 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[615]),
			.N(gen[616]),
			.NE(gen[617]),

			.O(gen[675]),
			.E(gen[677]),

			.SO(gen[735]),
			.S(gen[736]),
			.SE(gen[737]),

			.SELF(gen[676]),
			.cell_state(gen[676])
		); 

/******************* CELL 677 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell677 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[616]),
			.N(gen[617]),
			.NE(gen[618]),

			.O(gen[676]),
			.E(gen[678]),

			.SO(gen[736]),
			.S(gen[737]),
			.SE(gen[738]),

			.SELF(gen[677]),
			.cell_state(gen[677])
		); 

/******************* CELL 678 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell678 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[617]),
			.N(gen[618]),
			.NE(gen[619]),

			.O(gen[677]),
			.E(gen[679]),

			.SO(gen[737]),
			.S(gen[738]),
			.SE(gen[739]),

			.SELF(gen[678]),
			.cell_state(gen[678])
		); 

/******************* CELL 679 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell679 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[618]),
			.N(gen[619]),
			.NE(gen[620]),

			.O(gen[678]),
			.E(gen[680]),

			.SO(gen[738]),
			.S(gen[739]),
			.SE(gen[740]),

			.SELF(gen[679]),
			.cell_state(gen[679])
		); 

/******************* CELL 680 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell680 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[619]),
			.N(gen[620]),
			.NE(gen[621]),

			.O(gen[679]),
			.E(gen[681]),

			.SO(gen[739]),
			.S(gen[740]),
			.SE(gen[741]),

			.SELF(gen[680]),
			.cell_state(gen[680])
		); 

/******************* CELL 681 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell681 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[620]),
			.N(gen[621]),
			.NE(gen[622]),

			.O(gen[680]),
			.E(gen[682]),

			.SO(gen[740]),
			.S(gen[741]),
			.SE(gen[742]),

			.SELF(gen[681]),
			.cell_state(gen[681])
		); 

/******************* CELL 682 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell682 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[621]),
			.N(gen[622]),
			.NE(gen[623]),

			.O(gen[681]),
			.E(gen[683]),

			.SO(gen[741]),
			.S(gen[742]),
			.SE(gen[743]),

			.SELF(gen[682]),
			.cell_state(gen[682])
		); 

/******************* CELL 683 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell683 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[622]),
			.N(gen[623]),
			.NE(gen[624]),

			.O(gen[682]),
			.E(gen[684]),

			.SO(gen[742]),
			.S(gen[743]),
			.SE(gen[744]),

			.SELF(gen[683]),
			.cell_state(gen[683])
		); 

/******************* CELL 684 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell684 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[623]),
			.N(gen[624]),
			.NE(gen[625]),

			.O(gen[683]),
			.E(gen[685]),

			.SO(gen[743]),
			.S(gen[744]),
			.SE(gen[745]),

			.SELF(gen[684]),
			.cell_state(gen[684])
		); 

/******************* CELL 685 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell685 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[624]),
			.N(gen[625]),
			.NE(gen[626]),

			.O(gen[684]),
			.E(gen[686]),

			.SO(gen[744]),
			.S(gen[745]),
			.SE(gen[746]),

			.SELF(gen[685]),
			.cell_state(gen[685])
		); 

/******************* CELL 686 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell686 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[625]),
			.N(gen[626]),
			.NE(gen[627]),

			.O(gen[685]),
			.E(gen[687]),

			.SO(gen[745]),
			.S(gen[746]),
			.SE(gen[747]),

			.SELF(gen[686]),
			.cell_state(gen[686])
		); 

/******************* CELL 687 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell687 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[626]),
			.N(gen[627]),
			.NE(gen[628]),

			.O(gen[686]),
			.E(gen[688]),

			.SO(gen[746]),
			.S(gen[747]),
			.SE(gen[748]),

			.SELF(gen[687]),
			.cell_state(gen[687])
		); 

/******************* CELL 688 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell688 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[627]),
			.N(gen[628]),
			.NE(gen[629]),

			.O(gen[687]),
			.E(gen[689]),

			.SO(gen[747]),
			.S(gen[748]),
			.SE(gen[749]),

			.SELF(gen[688]),
			.cell_state(gen[688])
		); 

/******************* CELL 689 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell689 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[628]),
			.N(gen[629]),
			.NE(gen[630]),

			.O(gen[688]),
			.E(gen[690]),

			.SO(gen[748]),
			.S(gen[749]),
			.SE(gen[750]),

			.SELF(gen[689]),
			.cell_state(gen[689])
		); 

/******************* CELL 690 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell690 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[629]),
			.N(gen[630]),
			.NE(gen[631]),

			.O(gen[689]),
			.E(gen[691]),

			.SO(gen[749]),
			.S(gen[750]),
			.SE(gen[751]),

			.SELF(gen[690]),
			.cell_state(gen[690])
		); 

/******************* CELL 691 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell691 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[630]),
			.N(gen[631]),
			.NE(gen[632]),

			.O(gen[690]),
			.E(gen[692]),

			.SO(gen[750]),
			.S(gen[751]),
			.SE(gen[752]),

			.SELF(gen[691]),
			.cell_state(gen[691])
		); 

/******************* CELL 692 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell692 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[631]),
			.N(gen[632]),
			.NE(gen[633]),

			.O(gen[691]),
			.E(gen[693]),

			.SO(gen[751]),
			.S(gen[752]),
			.SE(gen[753]),

			.SELF(gen[692]),
			.cell_state(gen[692])
		); 

/******************* CELL 693 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell693 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[632]),
			.N(gen[633]),
			.NE(gen[634]),

			.O(gen[692]),
			.E(gen[694]),

			.SO(gen[752]),
			.S(gen[753]),
			.SE(gen[754]),

			.SELF(gen[693]),
			.cell_state(gen[693])
		); 

/******************* CELL 694 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell694 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[633]),
			.N(gen[634]),
			.NE(gen[635]),

			.O(gen[693]),
			.E(gen[695]),

			.SO(gen[753]),
			.S(gen[754]),
			.SE(gen[755]),

			.SELF(gen[694]),
			.cell_state(gen[694])
		); 

/******************* CELL 695 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell695 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[634]),
			.N(gen[635]),
			.NE(gen[636]),

			.O(gen[694]),
			.E(gen[696]),

			.SO(gen[754]),
			.S(gen[755]),
			.SE(gen[756]),

			.SELF(gen[695]),
			.cell_state(gen[695])
		); 

/******************* CELL 696 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell696 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[635]),
			.N(gen[636]),
			.NE(gen[637]),

			.O(gen[695]),
			.E(gen[697]),

			.SO(gen[755]),
			.S(gen[756]),
			.SE(gen[757]),

			.SELF(gen[696]),
			.cell_state(gen[696])
		); 

/******************* CELL 697 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell697 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[636]),
			.N(gen[637]),
			.NE(gen[638]),

			.O(gen[696]),
			.E(gen[698]),

			.SO(gen[756]),
			.S(gen[757]),
			.SE(gen[758]),

			.SELF(gen[697]),
			.cell_state(gen[697])
		); 

/******************* CELL 698 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell698 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[637]),
			.N(gen[638]),
			.NE(gen[639]),

			.O(gen[697]),
			.E(gen[699]),

			.SO(gen[757]),
			.S(gen[758]),
			.SE(gen[759]),

			.SELF(gen[698]),
			.cell_state(gen[698])
		); 

/******************* CELL 699 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell699 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[638]),
			.N(gen[639]),
			.NE(gen[640]),

			.O(gen[698]),
			.E(gen[700]),

			.SO(gen[758]),
			.S(gen[759]),
			.SE(gen[760]),

			.SELF(gen[699]),
			.cell_state(gen[699])
		); 

/******************* CELL 700 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell700 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[639]),
			.N(gen[640]),
			.NE(gen[641]),

			.O(gen[699]),
			.E(gen[701]),

			.SO(gen[759]),
			.S(gen[760]),
			.SE(gen[761]),

			.SELF(gen[700]),
			.cell_state(gen[700])
		); 

/******************* CELL 701 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell701 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[640]),
			.N(gen[641]),
			.NE(gen[642]),

			.O(gen[700]),
			.E(gen[702]),

			.SO(gen[760]),
			.S(gen[761]),
			.SE(gen[762]),

			.SELF(gen[701]),
			.cell_state(gen[701])
		); 

/******************* CELL 702 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell702 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[641]),
			.N(gen[642]),
			.NE(gen[643]),

			.O(gen[701]),
			.E(gen[703]),

			.SO(gen[761]),
			.S(gen[762]),
			.SE(gen[763]),

			.SELF(gen[702]),
			.cell_state(gen[702])
		); 

/******************* CELL 703 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell703 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[642]),
			.N(gen[643]),
			.NE(gen[644]),

			.O(gen[702]),
			.E(gen[704]),

			.SO(gen[762]),
			.S(gen[763]),
			.SE(gen[764]),

			.SELF(gen[703]),
			.cell_state(gen[703])
		); 

/******************* CELL 704 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell704 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[643]),
			.N(gen[644]),
			.NE(gen[645]),

			.O(gen[703]),
			.E(gen[705]),

			.SO(gen[763]),
			.S(gen[764]),
			.SE(gen[765]),

			.SELF(gen[704]),
			.cell_state(gen[704])
		); 

/******************* CELL 705 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell705 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[644]),
			.N(gen[645]),
			.NE(gen[646]),

			.O(gen[704]),
			.E(gen[706]),

			.SO(gen[764]),
			.S(gen[765]),
			.SE(gen[766]),

			.SELF(gen[705]),
			.cell_state(gen[705])
		); 

/******************* CELL 706 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell706 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[645]),
			.N(gen[646]),
			.NE(gen[647]),

			.O(gen[705]),
			.E(gen[707]),

			.SO(gen[765]),
			.S(gen[766]),
			.SE(gen[767]),

			.SELF(gen[706]),
			.cell_state(gen[706])
		); 

/******************* CELL 707 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell707 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[646]),
			.N(gen[647]),
			.NE(gen[648]),

			.O(gen[706]),
			.E(gen[708]),

			.SO(gen[766]),
			.S(gen[767]),
			.SE(gen[768]),

			.SELF(gen[707]),
			.cell_state(gen[707])
		); 

/******************* CELL 708 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell708 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[647]),
			.N(gen[648]),
			.NE(gen[649]),

			.O(gen[707]),
			.E(gen[709]),

			.SO(gen[767]),
			.S(gen[768]),
			.SE(gen[769]),

			.SELF(gen[708]),
			.cell_state(gen[708])
		); 

/******************* CELL 709 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell709 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[648]),
			.N(gen[649]),
			.NE(gen[650]),

			.O(gen[708]),
			.E(gen[710]),

			.SO(gen[768]),
			.S(gen[769]),
			.SE(gen[770]),

			.SELF(gen[709]),
			.cell_state(gen[709])
		); 

/******************* CELL 710 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell710 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[649]),
			.N(gen[650]),
			.NE(gen[651]),

			.O(gen[709]),
			.E(gen[711]),

			.SO(gen[769]),
			.S(gen[770]),
			.SE(gen[771]),

			.SELF(gen[710]),
			.cell_state(gen[710])
		); 

/******************* CELL 711 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell711 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[650]),
			.N(gen[651]),
			.NE(gen[652]),

			.O(gen[710]),
			.E(gen[712]),

			.SO(gen[770]),
			.S(gen[771]),
			.SE(gen[772]),

			.SELF(gen[711]),
			.cell_state(gen[711])
		); 

/******************* CELL 712 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell712 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[651]),
			.N(gen[652]),
			.NE(gen[653]),

			.O(gen[711]),
			.E(gen[713]),

			.SO(gen[771]),
			.S(gen[772]),
			.SE(gen[773]),

			.SELF(gen[712]),
			.cell_state(gen[712])
		); 

/******************* CELL 713 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell713 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[652]),
			.N(gen[653]),
			.NE(gen[654]),

			.O(gen[712]),
			.E(gen[714]),

			.SO(gen[772]),
			.S(gen[773]),
			.SE(gen[774]),

			.SELF(gen[713]),
			.cell_state(gen[713])
		); 

/******************* CELL 714 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell714 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[653]),
			.N(gen[654]),
			.NE(gen[655]),

			.O(gen[713]),
			.E(gen[715]),

			.SO(gen[773]),
			.S(gen[774]),
			.SE(gen[775]),

			.SELF(gen[714]),
			.cell_state(gen[714])
		); 

/******************* CELL 715 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell715 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[654]),
			.N(gen[655]),
			.NE(gen[656]),

			.O(gen[714]),
			.E(gen[716]),

			.SO(gen[774]),
			.S(gen[775]),
			.SE(gen[776]),

			.SELF(gen[715]),
			.cell_state(gen[715])
		); 

/******************* CELL 716 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell716 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[655]),
			.N(gen[656]),
			.NE(gen[657]),

			.O(gen[715]),
			.E(gen[717]),

			.SO(gen[775]),
			.S(gen[776]),
			.SE(gen[777]),

			.SELF(gen[716]),
			.cell_state(gen[716])
		); 

/******************* CELL 717 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell717 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[656]),
			.N(gen[657]),
			.NE(gen[658]),

			.O(gen[716]),
			.E(gen[718]),

			.SO(gen[776]),
			.S(gen[777]),
			.SE(gen[778]),

			.SELF(gen[717]),
			.cell_state(gen[717])
		); 

/******************* CELL 718 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell718 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[657]),
			.N(gen[658]),
			.NE(gen[659]),

			.O(gen[717]),
			.E(gen[719]),

			.SO(gen[777]),
			.S(gen[778]),
			.SE(gen[779]),

			.SELF(gen[718]),
			.cell_state(gen[718])
		); 

/******************* CELL 719 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell719 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[658]),
			.N(gen[659]),
			.NE(gen[658]),

			.O(gen[718]),
			.E(gen[718]),

			.SO(gen[778]),
			.S(gen[779]),
			.SE(gen[778]),

			.SELF(gen[719]),
			.cell_state(gen[719])
		); 

/******************* CELL 720 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell720 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[661]),
			.N(gen[660]),
			.NE(gen[661]),

			.O(gen[721]),
			.E(gen[721]),

			.SO(gen[781]),
			.S(gen[780]),
			.SE(gen[781]),

			.SELF(gen[720]),
			.cell_state(gen[720])
		); 

/******************* CELL 721 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell721 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[660]),
			.N(gen[661]),
			.NE(gen[662]),

			.O(gen[720]),
			.E(gen[722]),

			.SO(gen[780]),
			.S(gen[781]),
			.SE(gen[782]),

			.SELF(gen[721]),
			.cell_state(gen[721])
		); 

/******************* CELL 722 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell722 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[661]),
			.N(gen[662]),
			.NE(gen[663]),

			.O(gen[721]),
			.E(gen[723]),

			.SO(gen[781]),
			.S(gen[782]),
			.SE(gen[783]),

			.SELF(gen[722]),
			.cell_state(gen[722])
		); 

/******************* CELL 723 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell723 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[662]),
			.N(gen[663]),
			.NE(gen[664]),

			.O(gen[722]),
			.E(gen[724]),

			.SO(gen[782]),
			.S(gen[783]),
			.SE(gen[784]),

			.SELF(gen[723]),
			.cell_state(gen[723])
		); 

/******************* CELL 724 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell724 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[663]),
			.N(gen[664]),
			.NE(gen[665]),

			.O(gen[723]),
			.E(gen[725]),

			.SO(gen[783]),
			.S(gen[784]),
			.SE(gen[785]),

			.SELF(gen[724]),
			.cell_state(gen[724])
		); 

/******************* CELL 725 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell725 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[664]),
			.N(gen[665]),
			.NE(gen[666]),

			.O(gen[724]),
			.E(gen[726]),

			.SO(gen[784]),
			.S(gen[785]),
			.SE(gen[786]),

			.SELF(gen[725]),
			.cell_state(gen[725])
		); 

/******************* CELL 726 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell726 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[665]),
			.N(gen[666]),
			.NE(gen[667]),

			.O(gen[725]),
			.E(gen[727]),

			.SO(gen[785]),
			.S(gen[786]),
			.SE(gen[787]),

			.SELF(gen[726]),
			.cell_state(gen[726])
		); 

/******************* CELL 727 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell727 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[666]),
			.N(gen[667]),
			.NE(gen[668]),

			.O(gen[726]),
			.E(gen[728]),

			.SO(gen[786]),
			.S(gen[787]),
			.SE(gen[788]),

			.SELF(gen[727]),
			.cell_state(gen[727])
		); 

/******************* CELL 728 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell728 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[667]),
			.N(gen[668]),
			.NE(gen[669]),

			.O(gen[727]),
			.E(gen[729]),

			.SO(gen[787]),
			.S(gen[788]),
			.SE(gen[789]),

			.SELF(gen[728]),
			.cell_state(gen[728])
		); 

/******************* CELL 729 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell729 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[668]),
			.N(gen[669]),
			.NE(gen[670]),

			.O(gen[728]),
			.E(gen[730]),

			.SO(gen[788]),
			.S(gen[789]),
			.SE(gen[790]),

			.SELF(gen[729]),
			.cell_state(gen[729])
		); 

/******************* CELL 730 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell730 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[669]),
			.N(gen[670]),
			.NE(gen[671]),

			.O(gen[729]),
			.E(gen[731]),

			.SO(gen[789]),
			.S(gen[790]),
			.SE(gen[791]),

			.SELF(gen[730]),
			.cell_state(gen[730])
		); 

/******************* CELL 731 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell731 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[670]),
			.N(gen[671]),
			.NE(gen[672]),

			.O(gen[730]),
			.E(gen[732]),

			.SO(gen[790]),
			.S(gen[791]),
			.SE(gen[792]),

			.SELF(gen[731]),
			.cell_state(gen[731])
		); 

/******************* CELL 732 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell732 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[671]),
			.N(gen[672]),
			.NE(gen[673]),

			.O(gen[731]),
			.E(gen[733]),

			.SO(gen[791]),
			.S(gen[792]),
			.SE(gen[793]),

			.SELF(gen[732]),
			.cell_state(gen[732])
		); 

/******************* CELL 733 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell733 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[672]),
			.N(gen[673]),
			.NE(gen[674]),

			.O(gen[732]),
			.E(gen[734]),

			.SO(gen[792]),
			.S(gen[793]),
			.SE(gen[794]),

			.SELF(gen[733]),
			.cell_state(gen[733])
		); 

/******************* CELL 734 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell734 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[673]),
			.N(gen[674]),
			.NE(gen[675]),

			.O(gen[733]),
			.E(gen[735]),

			.SO(gen[793]),
			.S(gen[794]),
			.SE(gen[795]),

			.SELF(gen[734]),
			.cell_state(gen[734])
		); 

/******************* CELL 735 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell735 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[674]),
			.N(gen[675]),
			.NE(gen[676]),

			.O(gen[734]),
			.E(gen[736]),

			.SO(gen[794]),
			.S(gen[795]),
			.SE(gen[796]),

			.SELF(gen[735]),
			.cell_state(gen[735])
		); 

/******************* CELL 736 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell736 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[675]),
			.N(gen[676]),
			.NE(gen[677]),

			.O(gen[735]),
			.E(gen[737]),

			.SO(gen[795]),
			.S(gen[796]),
			.SE(gen[797]),

			.SELF(gen[736]),
			.cell_state(gen[736])
		); 

/******************* CELL 737 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell737 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[676]),
			.N(gen[677]),
			.NE(gen[678]),

			.O(gen[736]),
			.E(gen[738]),

			.SO(gen[796]),
			.S(gen[797]),
			.SE(gen[798]),

			.SELF(gen[737]),
			.cell_state(gen[737])
		); 

/******************* CELL 738 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell738 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[677]),
			.N(gen[678]),
			.NE(gen[679]),

			.O(gen[737]),
			.E(gen[739]),

			.SO(gen[797]),
			.S(gen[798]),
			.SE(gen[799]),

			.SELF(gen[738]),
			.cell_state(gen[738])
		); 

/******************* CELL 739 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell739 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[678]),
			.N(gen[679]),
			.NE(gen[680]),

			.O(gen[738]),
			.E(gen[740]),

			.SO(gen[798]),
			.S(gen[799]),
			.SE(gen[800]),

			.SELF(gen[739]),
			.cell_state(gen[739])
		); 

/******************* CELL 740 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell740 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[679]),
			.N(gen[680]),
			.NE(gen[681]),

			.O(gen[739]),
			.E(gen[741]),

			.SO(gen[799]),
			.S(gen[800]),
			.SE(gen[801]),

			.SELF(gen[740]),
			.cell_state(gen[740])
		); 

/******************* CELL 741 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell741 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[680]),
			.N(gen[681]),
			.NE(gen[682]),

			.O(gen[740]),
			.E(gen[742]),

			.SO(gen[800]),
			.S(gen[801]),
			.SE(gen[802]),

			.SELF(gen[741]),
			.cell_state(gen[741])
		); 

/******************* CELL 742 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell742 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[681]),
			.N(gen[682]),
			.NE(gen[683]),

			.O(gen[741]),
			.E(gen[743]),

			.SO(gen[801]),
			.S(gen[802]),
			.SE(gen[803]),

			.SELF(gen[742]),
			.cell_state(gen[742])
		); 

/******************* CELL 743 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell743 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[682]),
			.N(gen[683]),
			.NE(gen[684]),

			.O(gen[742]),
			.E(gen[744]),

			.SO(gen[802]),
			.S(gen[803]),
			.SE(gen[804]),

			.SELF(gen[743]),
			.cell_state(gen[743])
		); 

/******************* CELL 744 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell744 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[683]),
			.N(gen[684]),
			.NE(gen[685]),

			.O(gen[743]),
			.E(gen[745]),

			.SO(gen[803]),
			.S(gen[804]),
			.SE(gen[805]),

			.SELF(gen[744]),
			.cell_state(gen[744])
		); 

/******************* CELL 745 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell745 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[684]),
			.N(gen[685]),
			.NE(gen[686]),

			.O(gen[744]),
			.E(gen[746]),

			.SO(gen[804]),
			.S(gen[805]),
			.SE(gen[806]),

			.SELF(gen[745]),
			.cell_state(gen[745])
		); 

/******************* CELL 746 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell746 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[685]),
			.N(gen[686]),
			.NE(gen[687]),

			.O(gen[745]),
			.E(gen[747]),

			.SO(gen[805]),
			.S(gen[806]),
			.SE(gen[807]),

			.SELF(gen[746]),
			.cell_state(gen[746])
		); 

/******************* CELL 747 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell747 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[686]),
			.N(gen[687]),
			.NE(gen[688]),

			.O(gen[746]),
			.E(gen[748]),

			.SO(gen[806]),
			.S(gen[807]),
			.SE(gen[808]),

			.SELF(gen[747]),
			.cell_state(gen[747])
		); 

/******************* CELL 748 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell748 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[687]),
			.N(gen[688]),
			.NE(gen[689]),

			.O(gen[747]),
			.E(gen[749]),

			.SO(gen[807]),
			.S(gen[808]),
			.SE(gen[809]),

			.SELF(gen[748]),
			.cell_state(gen[748])
		); 

/******************* CELL 749 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell749 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[688]),
			.N(gen[689]),
			.NE(gen[690]),

			.O(gen[748]),
			.E(gen[750]),

			.SO(gen[808]),
			.S(gen[809]),
			.SE(gen[810]),

			.SELF(gen[749]),
			.cell_state(gen[749])
		); 

/******************* CELL 750 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell750 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[689]),
			.N(gen[690]),
			.NE(gen[691]),

			.O(gen[749]),
			.E(gen[751]),

			.SO(gen[809]),
			.S(gen[810]),
			.SE(gen[811]),

			.SELF(gen[750]),
			.cell_state(gen[750])
		); 

/******************* CELL 751 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell751 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[690]),
			.N(gen[691]),
			.NE(gen[692]),

			.O(gen[750]),
			.E(gen[752]),

			.SO(gen[810]),
			.S(gen[811]),
			.SE(gen[812]),

			.SELF(gen[751]),
			.cell_state(gen[751])
		); 

/******************* CELL 752 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell752 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[691]),
			.N(gen[692]),
			.NE(gen[693]),

			.O(gen[751]),
			.E(gen[753]),

			.SO(gen[811]),
			.S(gen[812]),
			.SE(gen[813]),

			.SELF(gen[752]),
			.cell_state(gen[752])
		); 

/******************* CELL 753 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell753 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[692]),
			.N(gen[693]),
			.NE(gen[694]),

			.O(gen[752]),
			.E(gen[754]),

			.SO(gen[812]),
			.S(gen[813]),
			.SE(gen[814]),

			.SELF(gen[753]),
			.cell_state(gen[753])
		); 

/******************* CELL 754 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell754 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[693]),
			.N(gen[694]),
			.NE(gen[695]),

			.O(gen[753]),
			.E(gen[755]),

			.SO(gen[813]),
			.S(gen[814]),
			.SE(gen[815]),

			.SELF(gen[754]),
			.cell_state(gen[754])
		); 

/******************* CELL 755 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell755 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[694]),
			.N(gen[695]),
			.NE(gen[696]),

			.O(gen[754]),
			.E(gen[756]),

			.SO(gen[814]),
			.S(gen[815]),
			.SE(gen[816]),

			.SELF(gen[755]),
			.cell_state(gen[755])
		); 

/******************* CELL 756 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell756 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[695]),
			.N(gen[696]),
			.NE(gen[697]),

			.O(gen[755]),
			.E(gen[757]),

			.SO(gen[815]),
			.S(gen[816]),
			.SE(gen[817]),

			.SELF(gen[756]),
			.cell_state(gen[756])
		); 

/******************* CELL 757 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell757 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[696]),
			.N(gen[697]),
			.NE(gen[698]),

			.O(gen[756]),
			.E(gen[758]),

			.SO(gen[816]),
			.S(gen[817]),
			.SE(gen[818]),

			.SELF(gen[757]),
			.cell_state(gen[757])
		); 

/******************* CELL 758 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell758 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[697]),
			.N(gen[698]),
			.NE(gen[699]),

			.O(gen[757]),
			.E(gen[759]),

			.SO(gen[817]),
			.S(gen[818]),
			.SE(gen[819]),

			.SELF(gen[758]),
			.cell_state(gen[758])
		); 

/******************* CELL 759 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell759 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[698]),
			.N(gen[699]),
			.NE(gen[700]),

			.O(gen[758]),
			.E(gen[760]),

			.SO(gen[818]),
			.S(gen[819]),
			.SE(gen[820]),

			.SELF(gen[759]),
			.cell_state(gen[759])
		); 

/******************* CELL 760 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell760 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[699]),
			.N(gen[700]),
			.NE(gen[701]),

			.O(gen[759]),
			.E(gen[761]),

			.SO(gen[819]),
			.S(gen[820]),
			.SE(gen[821]),

			.SELF(gen[760]),
			.cell_state(gen[760])
		); 

/******************* CELL 761 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell761 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[700]),
			.N(gen[701]),
			.NE(gen[702]),

			.O(gen[760]),
			.E(gen[762]),

			.SO(gen[820]),
			.S(gen[821]),
			.SE(gen[822]),

			.SELF(gen[761]),
			.cell_state(gen[761])
		); 

/******************* CELL 762 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell762 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[701]),
			.N(gen[702]),
			.NE(gen[703]),

			.O(gen[761]),
			.E(gen[763]),

			.SO(gen[821]),
			.S(gen[822]),
			.SE(gen[823]),

			.SELF(gen[762]),
			.cell_state(gen[762])
		); 

/******************* CELL 763 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell763 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[702]),
			.N(gen[703]),
			.NE(gen[704]),

			.O(gen[762]),
			.E(gen[764]),

			.SO(gen[822]),
			.S(gen[823]),
			.SE(gen[824]),

			.SELF(gen[763]),
			.cell_state(gen[763])
		); 

/******************* CELL 764 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell764 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[703]),
			.N(gen[704]),
			.NE(gen[705]),

			.O(gen[763]),
			.E(gen[765]),

			.SO(gen[823]),
			.S(gen[824]),
			.SE(gen[825]),

			.SELF(gen[764]),
			.cell_state(gen[764])
		); 

/******************* CELL 765 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell765 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[704]),
			.N(gen[705]),
			.NE(gen[706]),

			.O(gen[764]),
			.E(gen[766]),

			.SO(gen[824]),
			.S(gen[825]),
			.SE(gen[826]),

			.SELF(gen[765]),
			.cell_state(gen[765])
		); 

/******************* CELL 766 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell766 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[705]),
			.N(gen[706]),
			.NE(gen[707]),

			.O(gen[765]),
			.E(gen[767]),

			.SO(gen[825]),
			.S(gen[826]),
			.SE(gen[827]),

			.SELF(gen[766]),
			.cell_state(gen[766])
		); 

/******************* CELL 767 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell767 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[706]),
			.N(gen[707]),
			.NE(gen[708]),

			.O(gen[766]),
			.E(gen[768]),

			.SO(gen[826]),
			.S(gen[827]),
			.SE(gen[828]),

			.SELF(gen[767]),
			.cell_state(gen[767])
		); 

/******************* CELL 768 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell768 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[707]),
			.N(gen[708]),
			.NE(gen[709]),

			.O(gen[767]),
			.E(gen[769]),

			.SO(gen[827]),
			.S(gen[828]),
			.SE(gen[829]),

			.SELF(gen[768]),
			.cell_state(gen[768])
		); 

/******************* CELL 769 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell769 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[708]),
			.N(gen[709]),
			.NE(gen[710]),

			.O(gen[768]),
			.E(gen[770]),

			.SO(gen[828]),
			.S(gen[829]),
			.SE(gen[830]),

			.SELF(gen[769]),
			.cell_state(gen[769])
		); 

/******************* CELL 770 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell770 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[709]),
			.N(gen[710]),
			.NE(gen[711]),

			.O(gen[769]),
			.E(gen[771]),

			.SO(gen[829]),
			.S(gen[830]),
			.SE(gen[831]),

			.SELF(gen[770]),
			.cell_state(gen[770])
		); 

/******************* CELL 771 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell771 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[710]),
			.N(gen[711]),
			.NE(gen[712]),

			.O(gen[770]),
			.E(gen[772]),

			.SO(gen[830]),
			.S(gen[831]),
			.SE(gen[832]),

			.SELF(gen[771]),
			.cell_state(gen[771])
		); 

/******************* CELL 772 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell772 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[711]),
			.N(gen[712]),
			.NE(gen[713]),

			.O(gen[771]),
			.E(gen[773]),

			.SO(gen[831]),
			.S(gen[832]),
			.SE(gen[833]),

			.SELF(gen[772]),
			.cell_state(gen[772])
		); 

/******************* CELL 773 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell773 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[712]),
			.N(gen[713]),
			.NE(gen[714]),

			.O(gen[772]),
			.E(gen[774]),

			.SO(gen[832]),
			.S(gen[833]),
			.SE(gen[834]),

			.SELF(gen[773]),
			.cell_state(gen[773])
		); 

/******************* CELL 774 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell774 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[713]),
			.N(gen[714]),
			.NE(gen[715]),

			.O(gen[773]),
			.E(gen[775]),

			.SO(gen[833]),
			.S(gen[834]),
			.SE(gen[835]),

			.SELF(gen[774]),
			.cell_state(gen[774])
		); 

/******************* CELL 775 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell775 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[714]),
			.N(gen[715]),
			.NE(gen[716]),

			.O(gen[774]),
			.E(gen[776]),

			.SO(gen[834]),
			.S(gen[835]),
			.SE(gen[836]),

			.SELF(gen[775]),
			.cell_state(gen[775])
		); 

/******************* CELL 776 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell776 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[715]),
			.N(gen[716]),
			.NE(gen[717]),

			.O(gen[775]),
			.E(gen[777]),

			.SO(gen[835]),
			.S(gen[836]),
			.SE(gen[837]),

			.SELF(gen[776]),
			.cell_state(gen[776])
		); 

/******************* CELL 777 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell777 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[716]),
			.N(gen[717]),
			.NE(gen[718]),

			.O(gen[776]),
			.E(gen[778]),

			.SO(gen[836]),
			.S(gen[837]),
			.SE(gen[838]),

			.SELF(gen[777]),
			.cell_state(gen[777])
		); 

/******************* CELL 778 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell778 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[717]),
			.N(gen[718]),
			.NE(gen[719]),

			.O(gen[777]),
			.E(gen[779]),

			.SO(gen[837]),
			.S(gen[838]),
			.SE(gen[839]),

			.SELF(gen[778]),
			.cell_state(gen[778])
		); 

/******************* CELL 779 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell779 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[718]),
			.N(gen[719]),
			.NE(gen[718]),

			.O(gen[778]),
			.E(gen[778]),

			.SO(gen[838]),
			.S(gen[839]),
			.SE(gen[838]),

			.SELF(gen[779]),
			.cell_state(gen[779])
		); 

/******************* CELL 780 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell780 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[721]),
			.N(gen[720]),
			.NE(gen[721]),

			.O(gen[781]),
			.E(gen[781]),

			.SO(gen[841]),
			.S(gen[840]),
			.SE(gen[841]),

			.SELF(gen[780]),
			.cell_state(gen[780])
		); 

/******************* CELL 781 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell781 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[720]),
			.N(gen[721]),
			.NE(gen[722]),

			.O(gen[780]),
			.E(gen[782]),

			.SO(gen[840]),
			.S(gen[841]),
			.SE(gen[842]),

			.SELF(gen[781]),
			.cell_state(gen[781])
		); 

/******************* CELL 782 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell782 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[721]),
			.N(gen[722]),
			.NE(gen[723]),

			.O(gen[781]),
			.E(gen[783]),

			.SO(gen[841]),
			.S(gen[842]),
			.SE(gen[843]),

			.SELF(gen[782]),
			.cell_state(gen[782])
		); 

/******************* CELL 783 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell783 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[722]),
			.N(gen[723]),
			.NE(gen[724]),

			.O(gen[782]),
			.E(gen[784]),

			.SO(gen[842]),
			.S(gen[843]),
			.SE(gen[844]),

			.SELF(gen[783]),
			.cell_state(gen[783])
		); 

/******************* CELL 784 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell784 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[723]),
			.N(gen[724]),
			.NE(gen[725]),

			.O(gen[783]),
			.E(gen[785]),

			.SO(gen[843]),
			.S(gen[844]),
			.SE(gen[845]),

			.SELF(gen[784]),
			.cell_state(gen[784])
		); 

/******************* CELL 785 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell785 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[724]),
			.N(gen[725]),
			.NE(gen[726]),

			.O(gen[784]),
			.E(gen[786]),

			.SO(gen[844]),
			.S(gen[845]),
			.SE(gen[846]),

			.SELF(gen[785]),
			.cell_state(gen[785])
		); 

/******************* CELL 786 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell786 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[725]),
			.N(gen[726]),
			.NE(gen[727]),

			.O(gen[785]),
			.E(gen[787]),

			.SO(gen[845]),
			.S(gen[846]),
			.SE(gen[847]),

			.SELF(gen[786]),
			.cell_state(gen[786])
		); 

/******************* CELL 787 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell787 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[726]),
			.N(gen[727]),
			.NE(gen[728]),

			.O(gen[786]),
			.E(gen[788]),

			.SO(gen[846]),
			.S(gen[847]),
			.SE(gen[848]),

			.SELF(gen[787]),
			.cell_state(gen[787])
		); 

/******************* CELL 788 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell788 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[727]),
			.N(gen[728]),
			.NE(gen[729]),

			.O(gen[787]),
			.E(gen[789]),

			.SO(gen[847]),
			.S(gen[848]),
			.SE(gen[849]),

			.SELF(gen[788]),
			.cell_state(gen[788])
		); 

/******************* CELL 789 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell789 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[728]),
			.N(gen[729]),
			.NE(gen[730]),

			.O(gen[788]),
			.E(gen[790]),

			.SO(gen[848]),
			.S(gen[849]),
			.SE(gen[850]),

			.SELF(gen[789]),
			.cell_state(gen[789])
		); 

/******************* CELL 790 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell790 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[729]),
			.N(gen[730]),
			.NE(gen[731]),

			.O(gen[789]),
			.E(gen[791]),

			.SO(gen[849]),
			.S(gen[850]),
			.SE(gen[851]),

			.SELF(gen[790]),
			.cell_state(gen[790])
		); 

/******************* CELL 791 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell791 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[730]),
			.N(gen[731]),
			.NE(gen[732]),

			.O(gen[790]),
			.E(gen[792]),

			.SO(gen[850]),
			.S(gen[851]),
			.SE(gen[852]),

			.SELF(gen[791]),
			.cell_state(gen[791])
		); 

/******************* CELL 792 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell792 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[731]),
			.N(gen[732]),
			.NE(gen[733]),

			.O(gen[791]),
			.E(gen[793]),

			.SO(gen[851]),
			.S(gen[852]),
			.SE(gen[853]),

			.SELF(gen[792]),
			.cell_state(gen[792])
		); 

/******************* CELL 793 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell793 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[732]),
			.N(gen[733]),
			.NE(gen[734]),

			.O(gen[792]),
			.E(gen[794]),

			.SO(gen[852]),
			.S(gen[853]),
			.SE(gen[854]),

			.SELF(gen[793]),
			.cell_state(gen[793])
		); 

/******************* CELL 794 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell794 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[733]),
			.N(gen[734]),
			.NE(gen[735]),

			.O(gen[793]),
			.E(gen[795]),

			.SO(gen[853]),
			.S(gen[854]),
			.SE(gen[855]),

			.SELF(gen[794]),
			.cell_state(gen[794])
		); 

/******************* CELL 795 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell795 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[734]),
			.N(gen[735]),
			.NE(gen[736]),

			.O(gen[794]),
			.E(gen[796]),

			.SO(gen[854]),
			.S(gen[855]),
			.SE(gen[856]),

			.SELF(gen[795]),
			.cell_state(gen[795])
		); 

/******************* CELL 796 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell796 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[735]),
			.N(gen[736]),
			.NE(gen[737]),

			.O(gen[795]),
			.E(gen[797]),

			.SO(gen[855]),
			.S(gen[856]),
			.SE(gen[857]),

			.SELF(gen[796]),
			.cell_state(gen[796])
		); 

/******************* CELL 797 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell797 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[736]),
			.N(gen[737]),
			.NE(gen[738]),

			.O(gen[796]),
			.E(gen[798]),

			.SO(gen[856]),
			.S(gen[857]),
			.SE(gen[858]),

			.SELF(gen[797]),
			.cell_state(gen[797])
		); 

/******************* CELL 798 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell798 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[737]),
			.N(gen[738]),
			.NE(gen[739]),

			.O(gen[797]),
			.E(gen[799]),

			.SO(gen[857]),
			.S(gen[858]),
			.SE(gen[859]),

			.SELF(gen[798]),
			.cell_state(gen[798])
		); 

/******************* CELL 799 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell799 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[738]),
			.N(gen[739]),
			.NE(gen[740]),

			.O(gen[798]),
			.E(gen[800]),

			.SO(gen[858]),
			.S(gen[859]),
			.SE(gen[860]),

			.SELF(gen[799]),
			.cell_state(gen[799])
		); 

/******************* CELL 800 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell800 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[739]),
			.N(gen[740]),
			.NE(gen[741]),

			.O(gen[799]),
			.E(gen[801]),

			.SO(gen[859]),
			.S(gen[860]),
			.SE(gen[861]),

			.SELF(gen[800]),
			.cell_state(gen[800])
		); 

/******************* CELL 801 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell801 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[740]),
			.N(gen[741]),
			.NE(gen[742]),

			.O(gen[800]),
			.E(gen[802]),

			.SO(gen[860]),
			.S(gen[861]),
			.SE(gen[862]),

			.SELF(gen[801]),
			.cell_state(gen[801])
		); 

/******************* CELL 802 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell802 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[741]),
			.N(gen[742]),
			.NE(gen[743]),

			.O(gen[801]),
			.E(gen[803]),

			.SO(gen[861]),
			.S(gen[862]),
			.SE(gen[863]),

			.SELF(gen[802]),
			.cell_state(gen[802])
		); 

/******************* CELL 803 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell803 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[742]),
			.N(gen[743]),
			.NE(gen[744]),

			.O(gen[802]),
			.E(gen[804]),

			.SO(gen[862]),
			.S(gen[863]),
			.SE(gen[864]),

			.SELF(gen[803]),
			.cell_state(gen[803])
		); 

/******************* CELL 804 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell804 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[743]),
			.N(gen[744]),
			.NE(gen[745]),

			.O(gen[803]),
			.E(gen[805]),

			.SO(gen[863]),
			.S(gen[864]),
			.SE(gen[865]),

			.SELF(gen[804]),
			.cell_state(gen[804])
		); 

/******************* CELL 805 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell805 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[744]),
			.N(gen[745]),
			.NE(gen[746]),

			.O(gen[804]),
			.E(gen[806]),

			.SO(gen[864]),
			.S(gen[865]),
			.SE(gen[866]),

			.SELF(gen[805]),
			.cell_state(gen[805])
		); 

/******************* CELL 806 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell806 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[745]),
			.N(gen[746]),
			.NE(gen[747]),

			.O(gen[805]),
			.E(gen[807]),

			.SO(gen[865]),
			.S(gen[866]),
			.SE(gen[867]),

			.SELF(gen[806]),
			.cell_state(gen[806])
		); 

/******************* CELL 807 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell807 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[746]),
			.N(gen[747]),
			.NE(gen[748]),

			.O(gen[806]),
			.E(gen[808]),

			.SO(gen[866]),
			.S(gen[867]),
			.SE(gen[868]),

			.SELF(gen[807]),
			.cell_state(gen[807])
		); 

/******************* CELL 808 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell808 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[747]),
			.N(gen[748]),
			.NE(gen[749]),

			.O(gen[807]),
			.E(gen[809]),

			.SO(gen[867]),
			.S(gen[868]),
			.SE(gen[869]),

			.SELF(gen[808]),
			.cell_state(gen[808])
		); 

/******************* CELL 809 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell809 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[748]),
			.N(gen[749]),
			.NE(gen[750]),

			.O(gen[808]),
			.E(gen[810]),

			.SO(gen[868]),
			.S(gen[869]),
			.SE(gen[870]),

			.SELF(gen[809]),
			.cell_state(gen[809])
		); 

/******************* CELL 810 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell810 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[749]),
			.N(gen[750]),
			.NE(gen[751]),

			.O(gen[809]),
			.E(gen[811]),

			.SO(gen[869]),
			.S(gen[870]),
			.SE(gen[871]),

			.SELF(gen[810]),
			.cell_state(gen[810])
		); 

/******************* CELL 811 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell811 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[750]),
			.N(gen[751]),
			.NE(gen[752]),

			.O(gen[810]),
			.E(gen[812]),

			.SO(gen[870]),
			.S(gen[871]),
			.SE(gen[872]),

			.SELF(gen[811]),
			.cell_state(gen[811])
		); 

/******************* CELL 812 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell812 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[751]),
			.N(gen[752]),
			.NE(gen[753]),

			.O(gen[811]),
			.E(gen[813]),

			.SO(gen[871]),
			.S(gen[872]),
			.SE(gen[873]),

			.SELF(gen[812]),
			.cell_state(gen[812])
		); 

/******************* CELL 813 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell813 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[752]),
			.N(gen[753]),
			.NE(gen[754]),

			.O(gen[812]),
			.E(gen[814]),

			.SO(gen[872]),
			.S(gen[873]),
			.SE(gen[874]),

			.SELF(gen[813]),
			.cell_state(gen[813])
		); 

/******************* CELL 814 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell814 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[753]),
			.N(gen[754]),
			.NE(gen[755]),

			.O(gen[813]),
			.E(gen[815]),

			.SO(gen[873]),
			.S(gen[874]),
			.SE(gen[875]),

			.SELF(gen[814]),
			.cell_state(gen[814])
		); 

/******************* CELL 815 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell815 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[754]),
			.N(gen[755]),
			.NE(gen[756]),

			.O(gen[814]),
			.E(gen[816]),

			.SO(gen[874]),
			.S(gen[875]),
			.SE(gen[876]),

			.SELF(gen[815]),
			.cell_state(gen[815])
		); 

/******************* CELL 816 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell816 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[755]),
			.N(gen[756]),
			.NE(gen[757]),

			.O(gen[815]),
			.E(gen[817]),

			.SO(gen[875]),
			.S(gen[876]),
			.SE(gen[877]),

			.SELF(gen[816]),
			.cell_state(gen[816])
		); 

/******************* CELL 817 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell817 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[756]),
			.N(gen[757]),
			.NE(gen[758]),

			.O(gen[816]),
			.E(gen[818]),

			.SO(gen[876]),
			.S(gen[877]),
			.SE(gen[878]),

			.SELF(gen[817]),
			.cell_state(gen[817])
		); 

/******************* CELL 818 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell818 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[757]),
			.N(gen[758]),
			.NE(gen[759]),

			.O(gen[817]),
			.E(gen[819]),

			.SO(gen[877]),
			.S(gen[878]),
			.SE(gen[879]),

			.SELF(gen[818]),
			.cell_state(gen[818])
		); 

/******************* CELL 819 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell819 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[758]),
			.N(gen[759]),
			.NE(gen[760]),

			.O(gen[818]),
			.E(gen[820]),

			.SO(gen[878]),
			.S(gen[879]),
			.SE(gen[880]),

			.SELF(gen[819]),
			.cell_state(gen[819])
		); 

/******************* CELL 820 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell820 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[759]),
			.N(gen[760]),
			.NE(gen[761]),

			.O(gen[819]),
			.E(gen[821]),

			.SO(gen[879]),
			.S(gen[880]),
			.SE(gen[881]),

			.SELF(gen[820]),
			.cell_state(gen[820])
		); 

/******************* CELL 821 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell821 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[760]),
			.N(gen[761]),
			.NE(gen[762]),

			.O(gen[820]),
			.E(gen[822]),

			.SO(gen[880]),
			.S(gen[881]),
			.SE(gen[882]),

			.SELF(gen[821]),
			.cell_state(gen[821])
		); 

/******************* CELL 822 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell822 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[761]),
			.N(gen[762]),
			.NE(gen[763]),

			.O(gen[821]),
			.E(gen[823]),

			.SO(gen[881]),
			.S(gen[882]),
			.SE(gen[883]),

			.SELF(gen[822]),
			.cell_state(gen[822])
		); 

/******************* CELL 823 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell823 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[762]),
			.N(gen[763]),
			.NE(gen[764]),

			.O(gen[822]),
			.E(gen[824]),

			.SO(gen[882]),
			.S(gen[883]),
			.SE(gen[884]),

			.SELF(gen[823]),
			.cell_state(gen[823])
		); 

/******************* CELL 824 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell824 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[763]),
			.N(gen[764]),
			.NE(gen[765]),

			.O(gen[823]),
			.E(gen[825]),

			.SO(gen[883]),
			.S(gen[884]),
			.SE(gen[885]),

			.SELF(gen[824]),
			.cell_state(gen[824])
		); 

/******************* CELL 825 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell825 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[764]),
			.N(gen[765]),
			.NE(gen[766]),

			.O(gen[824]),
			.E(gen[826]),

			.SO(gen[884]),
			.S(gen[885]),
			.SE(gen[886]),

			.SELF(gen[825]),
			.cell_state(gen[825])
		); 

/******************* CELL 826 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell826 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[765]),
			.N(gen[766]),
			.NE(gen[767]),

			.O(gen[825]),
			.E(gen[827]),

			.SO(gen[885]),
			.S(gen[886]),
			.SE(gen[887]),

			.SELF(gen[826]),
			.cell_state(gen[826])
		); 

/******************* CELL 827 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell827 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[766]),
			.N(gen[767]),
			.NE(gen[768]),

			.O(gen[826]),
			.E(gen[828]),

			.SO(gen[886]),
			.S(gen[887]),
			.SE(gen[888]),

			.SELF(gen[827]),
			.cell_state(gen[827])
		); 

/******************* CELL 828 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell828 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[767]),
			.N(gen[768]),
			.NE(gen[769]),

			.O(gen[827]),
			.E(gen[829]),

			.SO(gen[887]),
			.S(gen[888]),
			.SE(gen[889]),

			.SELF(gen[828]),
			.cell_state(gen[828])
		); 

/******************* CELL 829 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell829 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[768]),
			.N(gen[769]),
			.NE(gen[770]),

			.O(gen[828]),
			.E(gen[830]),

			.SO(gen[888]),
			.S(gen[889]),
			.SE(gen[890]),

			.SELF(gen[829]),
			.cell_state(gen[829])
		); 

/******************* CELL 830 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell830 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[769]),
			.N(gen[770]),
			.NE(gen[771]),

			.O(gen[829]),
			.E(gen[831]),

			.SO(gen[889]),
			.S(gen[890]),
			.SE(gen[891]),

			.SELF(gen[830]),
			.cell_state(gen[830])
		); 

/******************* CELL 831 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell831 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[770]),
			.N(gen[771]),
			.NE(gen[772]),

			.O(gen[830]),
			.E(gen[832]),

			.SO(gen[890]),
			.S(gen[891]),
			.SE(gen[892]),

			.SELF(gen[831]),
			.cell_state(gen[831])
		); 

/******************* CELL 832 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell832 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[771]),
			.N(gen[772]),
			.NE(gen[773]),

			.O(gen[831]),
			.E(gen[833]),

			.SO(gen[891]),
			.S(gen[892]),
			.SE(gen[893]),

			.SELF(gen[832]),
			.cell_state(gen[832])
		); 

/******************* CELL 833 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell833 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[772]),
			.N(gen[773]),
			.NE(gen[774]),

			.O(gen[832]),
			.E(gen[834]),

			.SO(gen[892]),
			.S(gen[893]),
			.SE(gen[894]),

			.SELF(gen[833]),
			.cell_state(gen[833])
		); 

/******************* CELL 834 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell834 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[773]),
			.N(gen[774]),
			.NE(gen[775]),

			.O(gen[833]),
			.E(gen[835]),

			.SO(gen[893]),
			.S(gen[894]),
			.SE(gen[895]),

			.SELF(gen[834]),
			.cell_state(gen[834])
		); 

/******************* CELL 835 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell835 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[774]),
			.N(gen[775]),
			.NE(gen[776]),

			.O(gen[834]),
			.E(gen[836]),

			.SO(gen[894]),
			.S(gen[895]),
			.SE(gen[896]),

			.SELF(gen[835]),
			.cell_state(gen[835])
		); 

/******************* CELL 836 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell836 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[775]),
			.N(gen[776]),
			.NE(gen[777]),

			.O(gen[835]),
			.E(gen[837]),

			.SO(gen[895]),
			.S(gen[896]),
			.SE(gen[897]),

			.SELF(gen[836]),
			.cell_state(gen[836])
		); 

/******************* CELL 837 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell837 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[776]),
			.N(gen[777]),
			.NE(gen[778]),

			.O(gen[836]),
			.E(gen[838]),

			.SO(gen[896]),
			.S(gen[897]),
			.SE(gen[898]),

			.SELF(gen[837]),
			.cell_state(gen[837])
		); 

/******************* CELL 838 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell838 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[777]),
			.N(gen[778]),
			.NE(gen[779]),

			.O(gen[837]),
			.E(gen[839]),

			.SO(gen[897]),
			.S(gen[898]),
			.SE(gen[899]),

			.SELF(gen[838]),
			.cell_state(gen[838])
		); 

/******************* CELL 839 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell839 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[778]),
			.N(gen[779]),
			.NE(gen[778]),

			.O(gen[838]),
			.E(gen[838]),

			.SO(gen[898]),
			.S(gen[899]),
			.SE(gen[898]),

			.SELF(gen[839]),
			.cell_state(gen[839])
		); 

/******************* CELL 840 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell840 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[781]),
			.N(gen[780]),
			.NE(gen[781]),

			.O(gen[841]),
			.E(gen[841]),

			.SO(gen[901]),
			.S(gen[900]),
			.SE(gen[901]),

			.SELF(gen[840]),
			.cell_state(gen[840])
		); 

/******************* CELL 841 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell841 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[780]),
			.N(gen[781]),
			.NE(gen[782]),

			.O(gen[840]),
			.E(gen[842]),

			.SO(gen[900]),
			.S(gen[901]),
			.SE(gen[902]),

			.SELF(gen[841]),
			.cell_state(gen[841])
		); 

/******************* CELL 842 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell842 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[781]),
			.N(gen[782]),
			.NE(gen[783]),

			.O(gen[841]),
			.E(gen[843]),

			.SO(gen[901]),
			.S(gen[902]),
			.SE(gen[903]),

			.SELF(gen[842]),
			.cell_state(gen[842])
		); 

/******************* CELL 843 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell843 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[782]),
			.N(gen[783]),
			.NE(gen[784]),

			.O(gen[842]),
			.E(gen[844]),

			.SO(gen[902]),
			.S(gen[903]),
			.SE(gen[904]),

			.SELF(gen[843]),
			.cell_state(gen[843])
		); 

/******************* CELL 844 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell844 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[783]),
			.N(gen[784]),
			.NE(gen[785]),

			.O(gen[843]),
			.E(gen[845]),

			.SO(gen[903]),
			.S(gen[904]),
			.SE(gen[905]),

			.SELF(gen[844]),
			.cell_state(gen[844])
		); 

/******************* CELL 845 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell845 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[784]),
			.N(gen[785]),
			.NE(gen[786]),

			.O(gen[844]),
			.E(gen[846]),

			.SO(gen[904]),
			.S(gen[905]),
			.SE(gen[906]),

			.SELF(gen[845]),
			.cell_state(gen[845])
		); 

/******************* CELL 846 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell846 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[785]),
			.N(gen[786]),
			.NE(gen[787]),

			.O(gen[845]),
			.E(gen[847]),

			.SO(gen[905]),
			.S(gen[906]),
			.SE(gen[907]),

			.SELF(gen[846]),
			.cell_state(gen[846])
		); 

/******************* CELL 847 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell847 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[786]),
			.N(gen[787]),
			.NE(gen[788]),

			.O(gen[846]),
			.E(gen[848]),

			.SO(gen[906]),
			.S(gen[907]),
			.SE(gen[908]),

			.SELF(gen[847]),
			.cell_state(gen[847])
		); 

/******************* CELL 848 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell848 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[787]),
			.N(gen[788]),
			.NE(gen[789]),

			.O(gen[847]),
			.E(gen[849]),

			.SO(gen[907]),
			.S(gen[908]),
			.SE(gen[909]),

			.SELF(gen[848]),
			.cell_state(gen[848])
		); 

/******************* CELL 849 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell849 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[788]),
			.N(gen[789]),
			.NE(gen[790]),

			.O(gen[848]),
			.E(gen[850]),

			.SO(gen[908]),
			.S(gen[909]),
			.SE(gen[910]),

			.SELF(gen[849]),
			.cell_state(gen[849])
		); 

/******************* CELL 850 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell850 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[789]),
			.N(gen[790]),
			.NE(gen[791]),

			.O(gen[849]),
			.E(gen[851]),

			.SO(gen[909]),
			.S(gen[910]),
			.SE(gen[911]),

			.SELF(gen[850]),
			.cell_state(gen[850])
		); 

/******************* CELL 851 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell851 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[790]),
			.N(gen[791]),
			.NE(gen[792]),

			.O(gen[850]),
			.E(gen[852]),

			.SO(gen[910]),
			.S(gen[911]),
			.SE(gen[912]),

			.SELF(gen[851]),
			.cell_state(gen[851])
		); 

/******************* CELL 852 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell852 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[791]),
			.N(gen[792]),
			.NE(gen[793]),

			.O(gen[851]),
			.E(gen[853]),

			.SO(gen[911]),
			.S(gen[912]),
			.SE(gen[913]),

			.SELF(gen[852]),
			.cell_state(gen[852])
		); 

/******************* CELL 853 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell853 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[792]),
			.N(gen[793]),
			.NE(gen[794]),

			.O(gen[852]),
			.E(gen[854]),

			.SO(gen[912]),
			.S(gen[913]),
			.SE(gen[914]),

			.SELF(gen[853]),
			.cell_state(gen[853])
		); 

/******************* CELL 854 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell854 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[793]),
			.N(gen[794]),
			.NE(gen[795]),

			.O(gen[853]),
			.E(gen[855]),

			.SO(gen[913]),
			.S(gen[914]),
			.SE(gen[915]),

			.SELF(gen[854]),
			.cell_state(gen[854])
		); 

/******************* CELL 855 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell855 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[794]),
			.N(gen[795]),
			.NE(gen[796]),

			.O(gen[854]),
			.E(gen[856]),

			.SO(gen[914]),
			.S(gen[915]),
			.SE(gen[916]),

			.SELF(gen[855]),
			.cell_state(gen[855])
		); 

/******************* CELL 856 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell856 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[795]),
			.N(gen[796]),
			.NE(gen[797]),

			.O(gen[855]),
			.E(gen[857]),

			.SO(gen[915]),
			.S(gen[916]),
			.SE(gen[917]),

			.SELF(gen[856]),
			.cell_state(gen[856])
		); 

/******************* CELL 857 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell857 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[796]),
			.N(gen[797]),
			.NE(gen[798]),

			.O(gen[856]),
			.E(gen[858]),

			.SO(gen[916]),
			.S(gen[917]),
			.SE(gen[918]),

			.SELF(gen[857]),
			.cell_state(gen[857])
		); 

/******************* CELL 858 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell858 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[797]),
			.N(gen[798]),
			.NE(gen[799]),

			.O(gen[857]),
			.E(gen[859]),

			.SO(gen[917]),
			.S(gen[918]),
			.SE(gen[919]),

			.SELF(gen[858]),
			.cell_state(gen[858])
		); 

/******************* CELL 859 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell859 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[798]),
			.N(gen[799]),
			.NE(gen[800]),

			.O(gen[858]),
			.E(gen[860]),

			.SO(gen[918]),
			.S(gen[919]),
			.SE(gen[920]),

			.SELF(gen[859]),
			.cell_state(gen[859])
		); 

/******************* CELL 860 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell860 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[799]),
			.N(gen[800]),
			.NE(gen[801]),

			.O(gen[859]),
			.E(gen[861]),

			.SO(gen[919]),
			.S(gen[920]),
			.SE(gen[921]),

			.SELF(gen[860]),
			.cell_state(gen[860])
		); 

/******************* CELL 861 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell861 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[800]),
			.N(gen[801]),
			.NE(gen[802]),

			.O(gen[860]),
			.E(gen[862]),

			.SO(gen[920]),
			.S(gen[921]),
			.SE(gen[922]),

			.SELF(gen[861]),
			.cell_state(gen[861])
		); 

/******************* CELL 862 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell862 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[801]),
			.N(gen[802]),
			.NE(gen[803]),

			.O(gen[861]),
			.E(gen[863]),

			.SO(gen[921]),
			.S(gen[922]),
			.SE(gen[923]),

			.SELF(gen[862]),
			.cell_state(gen[862])
		); 

/******************* CELL 863 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell863 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[802]),
			.N(gen[803]),
			.NE(gen[804]),

			.O(gen[862]),
			.E(gen[864]),

			.SO(gen[922]),
			.S(gen[923]),
			.SE(gen[924]),

			.SELF(gen[863]),
			.cell_state(gen[863])
		); 

/******************* CELL 864 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell864 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[803]),
			.N(gen[804]),
			.NE(gen[805]),

			.O(gen[863]),
			.E(gen[865]),

			.SO(gen[923]),
			.S(gen[924]),
			.SE(gen[925]),

			.SELF(gen[864]),
			.cell_state(gen[864])
		); 

/******************* CELL 865 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell865 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[804]),
			.N(gen[805]),
			.NE(gen[806]),

			.O(gen[864]),
			.E(gen[866]),

			.SO(gen[924]),
			.S(gen[925]),
			.SE(gen[926]),

			.SELF(gen[865]),
			.cell_state(gen[865])
		); 

/******************* CELL 866 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell866 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[805]),
			.N(gen[806]),
			.NE(gen[807]),

			.O(gen[865]),
			.E(gen[867]),

			.SO(gen[925]),
			.S(gen[926]),
			.SE(gen[927]),

			.SELF(gen[866]),
			.cell_state(gen[866])
		); 

/******************* CELL 867 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell867 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[806]),
			.N(gen[807]),
			.NE(gen[808]),

			.O(gen[866]),
			.E(gen[868]),

			.SO(gen[926]),
			.S(gen[927]),
			.SE(gen[928]),

			.SELF(gen[867]),
			.cell_state(gen[867])
		); 

/******************* CELL 868 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell868 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[807]),
			.N(gen[808]),
			.NE(gen[809]),

			.O(gen[867]),
			.E(gen[869]),

			.SO(gen[927]),
			.S(gen[928]),
			.SE(gen[929]),

			.SELF(gen[868]),
			.cell_state(gen[868])
		); 

/******************* CELL 869 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell869 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[808]),
			.N(gen[809]),
			.NE(gen[810]),

			.O(gen[868]),
			.E(gen[870]),

			.SO(gen[928]),
			.S(gen[929]),
			.SE(gen[930]),

			.SELF(gen[869]),
			.cell_state(gen[869])
		); 

/******************* CELL 870 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell870 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[809]),
			.N(gen[810]),
			.NE(gen[811]),

			.O(gen[869]),
			.E(gen[871]),

			.SO(gen[929]),
			.S(gen[930]),
			.SE(gen[931]),

			.SELF(gen[870]),
			.cell_state(gen[870])
		); 

/******************* CELL 871 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell871 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[810]),
			.N(gen[811]),
			.NE(gen[812]),

			.O(gen[870]),
			.E(gen[872]),

			.SO(gen[930]),
			.S(gen[931]),
			.SE(gen[932]),

			.SELF(gen[871]),
			.cell_state(gen[871])
		); 

/******************* CELL 872 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell872 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[811]),
			.N(gen[812]),
			.NE(gen[813]),

			.O(gen[871]),
			.E(gen[873]),

			.SO(gen[931]),
			.S(gen[932]),
			.SE(gen[933]),

			.SELF(gen[872]),
			.cell_state(gen[872])
		); 

/******************* CELL 873 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell873 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[812]),
			.N(gen[813]),
			.NE(gen[814]),

			.O(gen[872]),
			.E(gen[874]),

			.SO(gen[932]),
			.S(gen[933]),
			.SE(gen[934]),

			.SELF(gen[873]),
			.cell_state(gen[873])
		); 

/******************* CELL 874 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell874 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[813]),
			.N(gen[814]),
			.NE(gen[815]),

			.O(gen[873]),
			.E(gen[875]),

			.SO(gen[933]),
			.S(gen[934]),
			.SE(gen[935]),

			.SELF(gen[874]),
			.cell_state(gen[874])
		); 

/******************* CELL 875 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell875 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[814]),
			.N(gen[815]),
			.NE(gen[816]),

			.O(gen[874]),
			.E(gen[876]),

			.SO(gen[934]),
			.S(gen[935]),
			.SE(gen[936]),

			.SELF(gen[875]),
			.cell_state(gen[875])
		); 

/******************* CELL 876 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell876 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[815]),
			.N(gen[816]),
			.NE(gen[817]),

			.O(gen[875]),
			.E(gen[877]),

			.SO(gen[935]),
			.S(gen[936]),
			.SE(gen[937]),

			.SELF(gen[876]),
			.cell_state(gen[876])
		); 

/******************* CELL 877 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell877 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[816]),
			.N(gen[817]),
			.NE(gen[818]),

			.O(gen[876]),
			.E(gen[878]),

			.SO(gen[936]),
			.S(gen[937]),
			.SE(gen[938]),

			.SELF(gen[877]),
			.cell_state(gen[877])
		); 

/******************* CELL 878 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell878 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[817]),
			.N(gen[818]),
			.NE(gen[819]),

			.O(gen[877]),
			.E(gen[879]),

			.SO(gen[937]),
			.S(gen[938]),
			.SE(gen[939]),

			.SELF(gen[878]),
			.cell_state(gen[878])
		); 

/******************* CELL 879 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell879 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[818]),
			.N(gen[819]),
			.NE(gen[820]),

			.O(gen[878]),
			.E(gen[880]),

			.SO(gen[938]),
			.S(gen[939]),
			.SE(gen[940]),

			.SELF(gen[879]),
			.cell_state(gen[879])
		); 

/******************* CELL 880 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell880 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[819]),
			.N(gen[820]),
			.NE(gen[821]),

			.O(gen[879]),
			.E(gen[881]),

			.SO(gen[939]),
			.S(gen[940]),
			.SE(gen[941]),

			.SELF(gen[880]),
			.cell_state(gen[880])
		); 

/******************* CELL 881 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell881 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[820]),
			.N(gen[821]),
			.NE(gen[822]),

			.O(gen[880]),
			.E(gen[882]),

			.SO(gen[940]),
			.S(gen[941]),
			.SE(gen[942]),

			.SELF(gen[881]),
			.cell_state(gen[881])
		); 

/******************* CELL 882 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell882 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[821]),
			.N(gen[822]),
			.NE(gen[823]),

			.O(gen[881]),
			.E(gen[883]),

			.SO(gen[941]),
			.S(gen[942]),
			.SE(gen[943]),

			.SELF(gen[882]),
			.cell_state(gen[882])
		); 

/******************* CELL 883 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell883 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[822]),
			.N(gen[823]),
			.NE(gen[824]),

			.O(gen[882]),
			.E(gen[884]),

			.SO(gen[942]),
			.S(gen[943]),
			.SE(gen[944]),

			.SELF(gen[883]),
			.cell_state(gen[883])
		); 

/******************* CELL 884 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell884 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[823]),
			.N(gen[824]),
			.NE(gen[825]),

			.O(gen[883]),
			.E(gen[885]),

			.SO(gen[943]),
			.S(gen[944]),
			.SE(gen[945]),

			.SELF(gen[884]),
			.cell_state(gen[884])
		); 

/******************* CELL 885 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell885 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[824]),
			.N(gen[825]),
			.NE(gen[826]),

			.O(gen[884]),
			.E(gen[886]),

			.SO(gen[944]),
			.S(gen[945]),
			.SE(gen[946]),

			.SELF(gen[885]),
			.cell_state(gen[885])
		); 

/******************* CELL 886 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell886 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[825]),
			.N(gen[826]),
			.NE(gen[827]),

			.O(gen[885]),
			.E(gen[887]),

			.SO(gen[945]),
			.S(gen[946]),
			.SE(gen[947]),

			.SELF(gen[886]),
			.cell_state(gen[886])
		); 

/******************* CELL 887 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell887 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[826]),
			.N(gen[827]),
			.NE(gen[828]),

			.O(gen[886]),
			.E(gen[888]),

			.SO(gen[946]),
			.S(gen[947]),
			.SE(gen[948]),

			.SELF(gen[887]),
			.cell_state(gen[887])
		); 

/******************* CELL 888 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell888 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[827]),
			.N(gen[828]),
			.NE(gen[829]),

			.O(gen[887]),
			.E(gen[889]),

			.SO(gen[947]),
			.S(gen[948]),
			.SE(gen[949]),

			.SELF(gen[888]),
			.cell_state(gen[888])
		); 

/******************* CELL 889 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell889 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[828]),
			.N(gen[829]),
			.NE(gen[830]),

			.O(gen[888]),
			.E(gen[890]),

			.SO(gen[948]),
			.S(gen[949]),
			.SE(gen[950]),

			.SELF(gen[889]),
			.cell_state(gen[889])
		); 

/******************* CELL 890 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell890 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[829]),
			.N(gen[830]),
			.NE(gen[831]),

			.O(gen[889]),
			.E(gen[891]),

			.SO(gen[949]),
			.S(gen[950]),
			.SE(gen[951]),

			.SELF(gen[890]),
			.cell_state(gen[890])
		); 

/******************* CELL 891 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell891 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[830]),
			.N(gen[831]),
			.NE(gen[832]),

			.O(gen[890]),
			.E(gen[892]),

			.SO(gen[950]),
			.S(gen[951]),
			.SE(gen[952]),

			.SELF(gen[891]),
			.cell_state(gen[891])
		); 

/******************* CELL 892 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell892 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[831]),
			.N(gen[832]),
			.NE(gen[833]),

			.O(gen[891]),
			.E(gen[893]),

			.SO(gen[951]),
			.S(gen[952]),
			.SE(gen[953]),

			.SELF(gen[892]),
			.cell_state(gen[892])
		); 

/******************* CELL 893 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell893 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[832]),
			.N(gen[833]),
			.NE(gen[834]),

			.O(gen[892]),
			.E(gen[894]),

			.SO(gen[952]),
			.S(gen[953]),
			.SE(gen[954]),

			.SELF(gen[893]),
			.cell_state(gen[893])
		); 

/******************* CELL 894 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell894 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[833]),
			.N(gen[834]),
			.NE(gen[835]),

			.O(gen[893]),
			.E(gen[895]),

			.SO(gen[953]),
			.S(gen[954]),
			.SE(gen[955]),

			.SELF(gen[894]),
			.cell_state(gen[894])
		); 

/******************* CELL 895 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell895 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[834]),
			.N(gen[835]),
			.NE(gen[836]),

			.O(gen[894]),
			.E(gen[896]),

			.SO(gen[954]),
			.S(gen[955]),
			.SE(gen[956]),

			.SELF(gen[895]),
			.cell_state(gen[895])
		); 

/******************* CELL 896 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell896 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[835]),
			.N(gen[836]),
			.NE(gen[837]),

			.O(gen[895]),
			.E(gen[897]),

			.SO(gen[955]),
			.S(gen[956]),
			.SE(gen[957]),

			.SELF(gen[896]),
			.cell_state(gen[896])
		); 

/******************* CELL 897 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell897 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[836]),
			.N(gen[837]),
			.NE(gen[838]),

			.O(gen[896]),
			.E(gen[898]),

			.SO(gen[956]),
			.S(gen[957]),
			.SE(gen[958]),

			.SELF(gen[897]),
			.cell_state(gen[897])
		); 

/******************* CELL 898 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell898 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[837]),
			.N(gen[838]),
			.NE(gen[839]),

			.O(gen[897]),
			.E(gen[899]),

			.SO(gen[957]),
			.S(gen[958]),
			.SE(gen[959]),

			.SELF(gen[898]),
			.cell_state(gen[898])
		); 

/******************* CELL 899 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell899 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[838]),
			.N(gen[839]),
			.NE(gen[838]),

			.O(gen[898]),
			.E(gen[898]),

			.SO(gen[958]),
			.S(gen[959]),
			.SE(gen[958]),

			.SELF(gen[899]),
			.cell_state(gen[899])
		); 

/******************* CELL 900 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell900 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[841]),
			.N(gen[840]),
			.NE(gen[841]),

			.O(gen[901]),
			.E(gen[901]),

			.SO(gen[961]),
			.S(gen[960]),
			.SE(gen[961]),

			.SELF(gen[900]),
			.cell_state(gen[900])
		); 

/******************* CELL 901 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell901 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[840]),
			.N(gen[841]),
			.NE(gen[842]),

			.O(gen[900]),
			.E(gen[902]),

			.SO(gen[960]),
			.S(gen[961]),
			.SE(gen[962]),

			.SELF(gen[901]),
			.cell_state(gen[901])
		); 

/******************* CELL 902 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell902 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[841]),
			.N(gen[842]),
			.NE(gen[843]),

			.O(gen[901]),
			.E(gen[903]),

			.SO(gen[961]),
			.S(gen[962]),
			.SE(gen[963]),

			.SELF(gen[902]),
			.cell_state(gen[902])
		); 

/******************* CELL 903 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell903 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[842]),
			.N(gen[843]),
			.NE(gen[844]),

			.O(gen[902]),
			.E(gen[904]),

			.SO(gen[962]),
			.S(gen[963]),
			.SE(gen[964]),

			.SELF(gen[903]),
			.cell_state(gen[903])
		); 

/******************* CELL 904 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell904 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[843]),
			.N(gen[844]),
			.NE(gen[845]),

			.O(gen[903]),
			.E(gen[905]),

			.SO(gen[963]),
			.S(gen[964]),
			.SE(gen[965]),

			.SELF(gen[904]),
			.cell_state(gen[904])
		); 

/******************* CELL 905 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell905 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[844]),
			.N(gen[845]),
			.NE(gen[846]),

			.O(gen[904]),
			.E(gen[906]),

			.SO(gen[964]),
			.S(gen[965]),
			.SE(gen[966]),

			.SELF(gen[905]),
			.cell_state(gen[905])
		); 

/******************* CELL 906 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell906 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[845]),
			.N(gen[846]),
			.NE(gen[847]),

			.O(gen[905]),
			.E(gen[907]),

			.SO(gen[965]),
			.S(gen[966]),
			.SE(gen[967]),

			.SELF(gen[906]),
			.cell_state(gen[906])
		); 

/******************* CELL 907 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell907 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[846]),
			.N(gen[847]),
			.NE(gen[848]),

			.O(gen[906]),
			.E(gen[908]),

			.SO(gen[966]),
			.S(gen[967]),
			.SE(gen[968]),

			.SELF(gen[907]),
			.cell_state(gen[907])
		); 

/******************* CELL 908 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell908 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[847]),
			.N(gen[848]),
			.NE(gen[849]),

			.O(gen[907]),
			.E(gen[909]),

			.SO(gen[967]),
			.S(gen[968]),
			.SE(gen[969]),

			.SELF(gen[908]),
			.cell_state(gen[908])
		); 

/******************* CELL 909 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell909 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[848]),
			.N(gen[849]),
			.NE(gen[850]),

			.O(gen[908]),
			.E(gen[910]),

			.SO(gen[968]),
			.S(gen[969]),
			.SE(gen[970]),

			.SELF(gen[909]),
			.cell_state(gen[909])
		); 

/******************* CELL 910 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell910 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[849]),
			.N(gen[850]),
			.NE(gen[851]),

			.O(gen[909]),
			.E(gen[911]),

			.SO(gen[969]),
			.S(gen[970]),
			.SE(gen[971]),

			.SELF(gen[910]),
			.cell_state(gen[910])
		); 

/******************* CELL 911 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell911 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[850]),
			.N(gen[851]),
			.NE(gen[852]),

			.O(gen[910]),
			.E(gen[912]),

			.SO(gen[970]),
			.S(gen[971]),
			.SE(gen[972]),

			.SELF(gen[911]),
			.cell_state(gen[911])
		); 

/******************* CELL 912 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell912 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[851]),
			.N(gen[852]),
			.NE(gen[853]),

			.O(gen[911]),
			.E(gen[913]),

			.SO(gen[971]),
			.S(gen[972]),
			.SE(gen[973]),

			.SELF(gen[912]),
			.cell_state(gen[912])
		); 

/******************* CELL 913 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell913 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[852]),
			.N(gen[853]),
			.NE(gen[854]),

			.O(gen[912]),
			.E(gen[914]),

			.SO(gen[972]),
			.S(gen[973]),
			.SE(gen[974]),

			.SELF(gen[913]),
			.cell_state(gen[913])
		); 

/******************* CELL 914 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell914 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[853]),
			.N(gen[854]),
			.NE(gen[855]),

			.O(gen[913]),
			.E(gen[915]),

			.SO(gen[973]),
			.S(gen[974]),
			.SE(gen[975]),

			.SELF(gen[914]),
			.cell_state(gen[914])
		); 

/******************* CELL 915 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell915 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[854]),
			.N(gen[855]),
			.NE(gen[856]),

			.O(gen[914]),
			.E(gen[916]),

			.SO(gen[974]),
			.S(gen[975]),
			.SE(gen[976]),

			.SELF(gen[915]),
			.cell_state(gen[915])
		); 

/******************* CELL 916 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell916 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[855]),
			.N(gen[856]),
			.NE(gen[857]),

			.O(gen[915]),
			.E(gen[917]),

			.SO(gen[975]),
			.S(gen[976]),
			.SE(gen[977]),

			.SELF(gen[916]),
			.cell_state(gen[916])
		); 

/******************* CELL 917 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell917 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[856]),
			.N(gen[857]),
			.NE(gen[858]),

			.O(gen[916]),
			.E(gen[918]),

			.SO(gen[976]),
			.S(gen[977]),
			.SE(gen[978]),

			.SELF(gen[917]),
			.cell_state(gen[917])
		); 

/******************* CELL 918 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell918 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[857]),
			.N(gen[858]),
			.NE(gen[859]),

			.O(gen[917]),
			.E(gen[919]),

			.SO(gen[977]),
			.S(gen[978]),
			.SE(gen[979]),

			.SELF(gen[918]),
			.cell_state(gen[918])
		); 

/******************* CELL 919 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell919 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[858]),
			.N(gen[859]),
			.NE(gen[860]),

			.O(gen[918]),
			.E(gen[920]),

			.SO(gen[978]),
			.S(gen[979]),
			.SE(gen[980]),

			.SELF(gen[919]),
			.cell_state(gen[919])
		); 

/******************* CELL 920 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell920 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[859]),
			.N(gen[860]),
			.NE(gen[861]),

			.O(gen[919]),
			.E(gen[921]),

			.SO(gen[979]),
			.S(gen[980]),
			.SE(gen[981]),

			.SELF(gen[920]),
			.cell_state(gen[920])
		); 

/******************* CELL 921 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell921 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[860]),
			.N(gen[861]),
			.NE(gen[862]),

			.O(gen[920]),
			.E(gen[922]),

			.SO(gen[980]),
			.S(gen[981]),
			.SE(gen[982]),

			.SELF(gen[921]),
			.cell_state(gen[921])
		); 

/******************* CELL 922 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell922 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[861]),
			.N(gen[862]),
			.NE(gen[863]),

			.O(gen[921]),
			.E(gen[923]),

			.SO(gen[981]),
			.S(gen[982]),
			.SE(gen[983]),

			.SELF(gen[922]),
			.cell_state(gen[922])
		); 

/******************* CELL 923 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell923 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[862]),
			.N(gen[863]),
			.NE(gen[864]),

			.O(gen[922]),
			.E(gen[924]),

			.SO(gen[982]),
			.S(gen[983]),
			.SE(gen[984]),

			.SELF(gen[923]),
			.cell_state(gen[923])
		); 

/******************* CELL 924 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell924 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[863]),
			.N(gen[864]),
			.NE(gen[865]),

			.O(gen[923]),
			.E(gen[925]),

			.SO(gen[983]),
			.S(gen[984]),
			.SE(gen[985]),

			.SELF(gen[924]),
			.cell_state(gen[924])
		); 

/******************* CELL 925 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell925 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[864]),
			.N(gen[865]),
			.NE(gen[866]),

			.O(gen[924]),
			.E(gen[926]),

			.SO(gen[984]),
			.S(gen[985]),
			.SE(gen[986]),

			.SELF(gen[925]),
			.cell_state(gen[925])
		); 

/******************* CELL 926 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell926 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[865]),
			.N(gen[866]),
			.NE(gen[867]),

			.O(gen[925]),
			.E(gen[927]),

			.SO(gen[985]),
			.S(gen[986]),
			.SE(gen[987]),

			.SELF(gen[926]),
			.cell_state(gen[926])
		); 

/******************* CELL 927 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell927 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[866]),
			.N(gen[867]),
			.NE(gen[868]),

			.O(gen[926]),
			.E(gen[928]),

			.SO(gen[986]),
			.S(gen[987]),
			.SE(gen[988]),

			.SELF(gen[927]),
			.cell_state(gen[927])
		); 

/******************* CELL 928 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell928 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[867]),
			.N(gen[868]),
			.NE(gen[869]),

			.O(gen[927]),
			.E(gen[929]),

			.SO(gen[987]),
			.S(gen[988]),
			.SE(gen[989]),

			.SELF(gen[928]),
			.cell_state(gen[928])
		); 

/******************* CELL 929 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell929 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[868]),
			.N(gen[869]),
			.NE(gen[870]),

			.O(gen[928]),
			.E(gen[930]),

			.SO(gen[988]),
			.S(gen[989]),
			.SE(gen[990]),

			.SELF(gen[929]),
			.cell_state(gen[929])
		); 

/******************* CELL 930 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell930 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[869]),
			.N(gen[870]),
			.NE(gen[871]),

			.O(gen[929]),
			.E(gen[931]),

			.SO(gen[989]),
			.S(gen[990]),
			.SE(gen[991]),

			.SELF(gen[930]),
			.cell_state(gen[930])
		); 

/******************* CELL 931 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell931 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[870]),
			.N(gen[871]),
			.NE(gen[872]),

			.O(gen[930]),
			.E(gen[932]),

			.SO(gen[990]),
			.S(gen[991]),
			.SE(gen[992]),

			.SELF(gen[931]),
			.cell_state(gen[931])
		); 

/******************* CELL 932 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell932 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[871]),
			.N(gen[872]),
			.NE(gen[873]),

			.O(gen[931]),
			.E(gen[933]),

			.SO(gen[991]),
			.S(gen[992]),
			.SE(gen[993]),

			.SELF(gen[932]),
			.cell_state(gen[932])
		); 

/******************* CELL 933 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell933 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[872]),
			.N(gen[873]),
			.NE(gen[874]),

			.O(gen[932]),
			.E(gen[934]),

			.SO(gen[992]),
			.S(gen[993]),
			.SE(gen[994]),

			.SELF(gen[933]),
			.cell_state(gen[933])
		); 

/******************* CELL 934 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell934 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[873]),
			.N(gen[874]),
			.NE(gen[875]),

			.O(gen[933]),
			.E(gen[935]),

			.SO(gen[993]),
			.S(gen[994]),
			.SE(gen[995]),

			.SELF(gen[934]),
			.cell_state(gen[934])
		); 

/******************* CELL 935 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell935 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[874]),
			.N(gen[875]),
			.NE(gen[876]),

			.O(gen[934]),
			.E(gen[936]),

			.SO(gen[994]),
			.S(gen[995]),
			.SE(gen[996]),

			.SELF(gen[935]),
			.cell_state(gen[935])
		); 

/******************* CELL 936 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell936 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[875]),
			.N(gen[876]),
			.NE(gen[877]),

			.O(gen[935]),
			.E(gen[937]),

			.SO(gen[995]),
			.S(gen[996]),
			.SE(gen[997]),

			.SELF(gen[936]),
			.cell_state(gen[936])
		); 

/******************* CELL 937 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell937 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[876]),
			.N(gen[877]),
			.NE(gen[878]),

			.O(gen[936]),
			.E(gen[938]),

			.SO(gen[996]),
			.S(gen[997]),
			.SE(gen[998]),

			.SELF(gen[937]),
			.cell_state(gen[937])
		); 

/******************* CELL 938 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell938 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[877]),
			.N(gen[878]),
			.NE(gen[879]),

			.O(gen[937]),
			.E(gen[939]),

			.SO(gen[997]),
			.S(gen[998]),
			.SE(gen[999]),

			.SELF(gen[938]),
			.cell_state(gen[938])
		); 

/******************* CELL 939 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell939 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[878]),
			.N(gen[879]),
			.NE(gen[880]),

			.O(gen[938]),
			.E(gen[940]),

			.SO(gen[998]),
			.S(gen[999]),
			.SE(gen[1000]),

			.SELF(gen[939]),
			.cell_state(gen[939])
		); 

/******************* CELL 940 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell940 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[879]),
			.N(gen[880]),
			.NE(gen[881]),

			.O(gen[939]),
			.E(gen[941]),

			.SO(gen[999]),
			.S(gen[1000]),
			.SE(gen[1001]),

			.SELF(gen[940]),
			.cell_state(gen[940])
		); 

/******************* CELL 941 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell941 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[880]),
			.N(gen[881]),
			.NE(gen[882]),

			.O(gen[940]),
			.E(gen[942]),

			.SO(gen[1000]),
			.S(gen[1001]),
			.SE(gen[1002]),

			.SELF(gen[941]),
			.cell_state(gen[941])
		); 

/******************* CELL 942 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell942 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[881]),
			.N(gen[882]),
			.NE(gen[883]),

			.O(gen[941]),
			.E(gen[943]),

			.SO(gen[1001]),
			.S(gen[1002]),
			.SE(gen[1003]),

			.SELF(gen[942]),
			.cell_state(gen[942])
		); 

/******************* CELL 943 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell943 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[882]),
			.N(gen[883]),
			.NE(gen[884]),

			.O(gen[942]),
			.E(gen[944]),

			.SO(gen[1002]),
			.S(gen[1003]),
			.SE(gen[1004]),

			.SELF(gen[943]),
			.cell_state(gen[943])
		); 

/******************* CELL 944 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell944 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[883]),
			.N(gen[884]),
			.NE(gen[885]),

			.O(gen[943]),
			.E(gen[945]),

			.SO(gen[1003]),
			.S(gen[1004]),
			.SE(gen[1005]),

			.SELF(gen[944]),
			.cell_state(gen[944])
		); 

/******************* CELL 945 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell945 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[884]),
			.N(gen[885]),
			.NE(gen[886]),

			.O(gen[944]),
			.E(gen[946]),

			.SO(gen[1004]),
			.S(gen[1005]),
			.SE(gen[1006]),

			.SELF(gen[945]),
			.cell_state(gen[945])
		); 

/******************* CELL 946 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell946 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[885]),
			.N(gen[886]),
			.NE(gen[887]),

			.O(gen[945]),
			.E(gen[947]),

			.SO(gen[1005]),
			.S(gen[1006]),
			.SE(gen[1007]),

			.SELF(gen[946]),
			.cell_state(gen[946])
		); 

/******************* CELL 947 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell947 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[886]),
			.N(gen[887]),
			.NE(gen[888]),

			.O(gen[946]),
			.E(gen[948]),

			.SO(gen[1006]),
			.S(gen[1007]),
			.SE(gen[1008]),

			.SELF(gen[947]),
			.cell_state(gen[947])
		); 

/******************* CELL 948 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell948 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[887]),
			.N(gen[888]),
			.NE(gen[889]),

			.O(gen[947]),
			.E(gen[949]),

			.SO(gen[1007]),
			.S(gen[1008]),
			.SE(gen[1009]),

			.SELF(gen[948]),
			.cell_state(gen[948])
		); 

/******************* CELL 949 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell949 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[888]),
			.N(gen[889]),
			.NE(gen[890]),

			.O(gen[948]),
			.E(gen[950]),

			.SO(gen[1008]),
			.S(gen[1009]),
			.SE(gen[1010]),

			.SELF(gen[949]),
			.cell_state(gen[949])
		); 

/******************* CELL 950 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell950 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[889]),
			.N(gen[890]),
			.NE(gen[891]),

			.O(gen[949]),
			.E(gen[951]),

			.SO(gen[1009]),
			.S(gen[1010]),
			.SE(gen[1011]),

			.SELF(gen[950]),
			.cell_state(gen[950])
		); 

/******************* CELL 951 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell951 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[890]),
			.N(gen[891]),
			.NE(gen[892]),

			.O(gen[950]),
			.E(gen[952]),

			.SO(gen[1010]),
			.S(gen[1011]),
			.SE(gen[1012]),

			.SELF(gen[951]),
			.cell_state(gen[951])
		); 

/******************* CELL 952 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell952 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[891]),
			.N(gen[892]),
			.NE(gen[893]),

			.O(gen[951]),
			.E(gen[953]),

			.SO(gen[1011]),
			.S(gen[1012]),
			.SE(gen[1013]),

			.SELF(gen[952]),
			.cell_state(gen[952])
		); 

/******************* CELL 953 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell953 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[892]),
			.N(gen[893]),
			.NE(gen[894]),

			.O(gen[952]),
			.E(gen[954]),

			.SO(gen[1012]),
			.S(gen[1013]),
			.SE(gen[1014]),

			.SELF(gen[953]),
			.cell_state(gen[953])
		); 

/******************* CELL 954 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell954 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[893]),
			.N(gen[894]),
			.NE(gen[895]),

			.O(gen[953]),
			.E(gen[955]),

			.SO(gen[1013]),
			.S(gen[1014]),
			.SE(gen[1015]),

			.SELF(gen[954]),
			.cell_state(gen[954])
		); 

/******************* CELL 955 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell955 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[894]),
			.N(gen[895]),
			.NE(gen[896]),

			.O(gen[954]),
			.E(gen[956]),

			.SO(gen[1014]),
			.S(gen[1015]),
			.SE(gen[1016]),

			.SELF(gen[955]),
			.cell_state(gen[955])
		); 

/******************* CELL 956 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell956 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[895]),
			.N(gen[896]),
			.NE(gen[897]),

			.O(gen[955]),
			.E(gen[957]),

			.SO(gen[1015]),
			.S(gen[1016]),
			.SE(gen[1017]),

			.SELF(gen[956]),
			.cell_state(gen[956])
		); 

/******************* CELL 957 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell957 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[896]),
			.N(gen[897]),
			.NE(gen[898]),

			.O(gen[956]),
			.E(gen[958]),

			.SO(gen[1016]),
			.S(gen[1017]),
			.SE(gen[1018]),

			.SELF(gen[957]),
			.cell_state(gen[957])
		); 

/******************* CELL 958 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell958 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[897]),
			.N(gen[898]),
			.NE(gen[899]),

			.O(gen[957]),
			.E(gen[959]),

			.SO(gen[1017]),
			.S(gen[1018]),
			.SE(gen[1019]),

			.SELF(gen[958]),
			.cell_state(gen[958])
		); 

/******************* CELL 959 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell959 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[898]),
			.N(gen[899]),
			.NE(gen[898]),

			.O(gen[958]),
			.E(gen[958]),

			.SO(gen[1018]),
			.S(gen[1019]),
			.SE(gen[1018]),

			.SELF(gen[959]),
			.cell_state(gen[959])
		); 

/******************* CELL 960 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell960 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[901]),
			.N(gen[900]),
			.NE(gen[901]),

			.O(gen[961]),
			.E(gen[961]),

			.SO(gen[1021]),
			.S(gen[1020]),
			.SE(gen[1021]),

			.SELF(gen[960]),
			.cell_state(gen[960])
		); 

/******************* CELL 961 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell961 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[900]),
			.N(gen[901]),
			.NE(gen[902]),

			.O(gen[960]),
			.E(gen[962]),

			.SO(gen[1020]),
			.S(gen[1021]),
			.SE(gen[1022]),

			.SELF(gen[961]),
			.cell_state(gen[961])
		); 

/******************* CELL 962 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell962 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[901]),
			.N(gen[902]),
			.NE(gen[903]),

			.O(gen[961]),
			.E(gen[963]),

			.SO(gen[1021]),
			.S(gen[1022]),
			.SE(gen[1023]),

			.SELF(gen[962]),
			.cell_state(gen[962])
		); 

/******************* CELL 963 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell963 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[902]),
			.N(gen[903]),
			.NE(gen[904]),

			.O(gen[962]),
			.E(gen[964]),

			.SO(gen[1022]),
			.S(gen[1023]),
			.SE(gen[1024]),

			.SELF(gen[963]),
			.cell_state(gen[963])
		); 

/******************* CELL 964 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell964 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[903]),
			.N(gen[904]),
			.NE(gen[905]),

			.O(gen[963]),
			.E(gen[965]),

			.SO(gen[1023]),
			.S(gen[1024]),
			.SE(gen[1025]),

			.SELF(gen[964]),
			.cell_state(gen[964])
		); 

/******************* CELL 965 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell965 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[904]),
			.N(gen[905]),
			.NE(gen[906]),

			.O(gen[964]),
			.E(gen[966]),

			.SO(gen[1024]),
			.S(gen[1025]),
			.SE(gen[1026]),

			.SELF(gen[965]),
			.cell_state(gen[965])
		); 

/******************* CELL 966 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell966 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[905]),
			.N(gen[906]),
			.NE(gen[907]),

			.O(gen[965]),
			.E(gen[967]),

			.SO(gen[1025]),
			.S(gen[1026]),
			.SE(gen[1027]),

			.SELF(gen[966]),
			.cell_state(gen[966])
		); 

/******************* CELL 967 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell967 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[906]),
			.N(gen[907]),
			.NE(gen[908]),

			.O(gen[966]),
			.E(gen[968]),

			.SO(gen[1026]),
			.S(gen[1027]),
			.SE(gen[1028]),

			.SELF(gen[967]),
			.cell_state(gen[967])
		); 

/******************* CELL 968 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell968 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[907]),
			.N(gen[908]),
			.NE(gen[909]),

			.O(gen[967]),
			.E(gen[969]),

			.SO(gen[1027]),
			.S(gen[1028]),
			.SE(gen[1029]),

			.SELF(gen[968]),
			.cell_state(gen[968])
		); 

/******************* CELL 969 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell969 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[908]),
			.N(gen[909]),
			.NE(gen[910]),

			.O(gen[968]),
			.E(gen[970]),

			.SO(gen[1028]),
			.S(gen[1029]),
			.SE(gen[1030]),

			.SELF(gen[969]),
			.cell_state(gen[969])
		); 

/******************* CELL 970 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell970 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[909]),
			.N(gen[910]),
			.NE(gen[911]),

			.O(gen[969]),
			.E(gen[971]),

			.SO(gen[1029]),
			.S(gen[1030]),
			.SE(gen[1031]),

			.SELF(gen[970]),
			.cell_state(gen[970])
		); 

/******************* CELL 971 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell971 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[910]),
			.N(gen[911]),
			.NE(gen[912]),

			.O(gen[970]),
			.E(gen[972]),

			.SO(gen[1030]),
			.S(gen[1031]),
			.SE(gen[1032]),

			.SELF(gen[971]),
			.cell_state(gen[971])
		); 

/******************* CELL 972 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell972 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[911]),
			.N(gen[912]),
			.NE(gen[913]),

			.O(gen[971]),
			.E(gen[973]),

			.SO(gen[1031]),
			.S(gen[1032]),
			.SE(gen[1033]),

			.SELF(gen[972]),
			.cell_state(gen[972])
		); 

/******************* CELL 973 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell973 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[912]),
			.N(gen[913]),
			.NE(gen[914]),

			.O(gen[972]),
			.E(gen[974]),

			.SO(gen[1032]),
			.S(gen[1033]),
			.SE(gen[1034]),

			.SELF(gen[973]),
			.cell_state(gen[973])
		); 

/******************* CELL 974 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell974 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[913]),
			.N(gen[914]),
			.NE(gen[915]),

			.O(gen[973]),
			.E(gen[975]),

			.SO(gen[1033]),
			.S(gen[1034]),
			.SE(gen[1035]),

			.SELF(gen[974]),
			.cell_state(gen[974])
		); 

/******************* CELL 975 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell975 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[914]),
			.N(gen[915]),
			.NE(gen[916]),

			.O(gen[974]),
			.E(gen[976]),

			.SO(gen[1034]),
			.S(gen[1035]),
			.SE(gen[1036]),

			.SELF(gen[975]),
			.cell_state(gen[975])
		); 

/******************* CELL 976 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell976 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[915]),
			.N(gen[916]),
			.NE(gen[917]),

			.O(gen[975]),
			.E(gen[977]),

			.SO(gen[1035]),
			.S(gen[1036]),
			.SE(gen[1037]),

			.SELF(gen[976]),
			.cell_state(gen[976])
		); 

/******************* CELL 977 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell977 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[916]),
			.N(gen[917]),
			.NE(gen[918]),

			.O(gen[976]),
			.E(gen[978]),

			.SO(gen[1036]),
			.S(gen[1037]),
			.SE(gen[1038]),

			.SELF(gen[977]),
			.cell_state(gen[977])
		); 

/******************* CELL 978 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell978 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[917]),
			.N(gen[918]),
			.NE(gen[919]),

			.O(gen[977]),
			.E(gen[979]),

			.SO(gen[1037]),
			.S(gen[1038]),
			.SE(gen[1039]),

			.SELF(gen[978]),
			.cell_state(gen[978])
		); 

/******************* CELL 979 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell979 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[918]),
			.N(gen[919]),
			.NE(gen[920]),

			.O(gen[978]),
			.E(gen[980]),

			.SO(gen[1038]),
			.S(gen[1039]),
			.SE(gen[1040]),

			.SELF(gen[979]),
			.cell_state(gen[979])
		); 

/******************* CELL 980 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell980 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[919]),
			.N(gen[920]),
			.NE(gen[921]),

			.O(gen[979]),
			.E(gen[981]),

			.SO(gen[1039]),
			.S(gen[1040]),
			.SE(gen[1041]),

			.SELF(gen[980]),
			.cell_state(gen[980])
		); 

/******************* CELL 981 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell981 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[920]),
			.N(gen[921]),
			.NE(gen[922]),

			.O(gen[980]),
			.E(gen[982]),

			.SO(gen[1040]),
			.S(gen[1041]),
			.SE(gen[1042]),

			.SELF(gen[981]),
			.cell_state(gen[981])
		); 

/******************* CELL 982 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell982 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[921]),
			.N(gen[922]),
			.NE(gen[923]),

			.O(gen[981]),
			.E(gen[983]),

			.SO(gen[1041]),
			.S(gen[1042]),
			.SE(gen[1043]),

			.SELF(gen[982]),
			.cell_state(gen[982])
		); 

/******************* CELL 983 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell983 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[922]),
			.N(gen[923]),
			.NE(gen[924]),

			.O(gen[982]),
			.E(gen[984]),

			.SO(gen[1042]),
			.S(gen[1043]),
			.SE(gen[1044]),

			.SELF(gen[983]),
			.cell_state(gen[983])
		); 

/******************* CELL 984 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell984 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[923]),
			.N(gen[924]),
			.NE(gen[925]),

			.O(gen[983]),
			.E(gen[985]),

			.SO(gen[1043]),
			.S(gen[1044]),
			.SE(gen[1045]),

			.SELF(gen[984]),
			.cell_state(gen[984])
		); 

/******************* CELL 985 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell985 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[924]),
			.N(gen[925]),
			.NE(gen[926]),

			.O(gen[984]),
			.E(gen[986]),

			.SO(gen[1044]),
			.S(gen[1045]),
			.SE(gen[1046]),

			.SELF(gen[985]),
			.cell_state(gen[985])
		); 

/******************* CELL 986 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell986 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[925]),
			.N(gen[926]),
			.NE(gen[927]),

			.O(gen[985]),
			.E(gen[987]),

			.SO(gen[1045]),
			.S(gen[1046]),
			.SE(gen[1047]),

			.SELF(gen[986]),
			.cell_state(gen[986])
		); 

/******************* CELL 987 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell987 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[926]),
			.N(gen[927]),
			.NE(gen[928]),

			.O(gen[986]),
			.E(gen[988]),

			.SO(gen[1046]),
			.S(gen[1047]),
			.SE(gen[1048]),

			.SELF(gen[987]),
			.cell_state(gen[987])
		); 

/******************* CELL 988 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell988 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[927]),
			.N(gen[928]),
			.NE(gen[929]),

			.O(gen[987]),
			.E(gen[989]),

			.SO(gen[1047]),
			.S(gen[1048]),
			.SE(gen[1049]),

			.SELF(gen[988]),
			.cell_state(gen[988])
		); 

/******************* CELL 989 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell989 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[928]),
			.N(gen[929]),
			.NE(gen[930]),

			.O(gen[988]),
			.E(gen[990]),

			.SO(gen[1048]),
			.S(gen[1049]),
			.SE(gen[1050]),

			.SELF(gen[989]),
			.cell_state(gen[989])
		); 

/******************* CELL 990 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell990 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[929]),
			.N(gen[930]),
			.NE(gen[931]),

			.O(gen[989]),
			.E(gen[991]),

			.SO(gen[1049]),
			.S(gen[1050]),
			.SE(gen[1051]),

			.SELF(gen[990]),
			.cell_state(gen[990])
		); 

/******************* CELL 991 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell991 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[930]),
			.N(gen[931]),
			.NE(gen[932]),

			.O(gen[990]),
			.E(gen[992]),

			.SO(gen[1050]),
			.S(gen[1051]),
			.SE(gen[1052]),

			.SELF(gen[991]),
			.cell_state(gen[991])
		); 

/******************* CELL 992 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell992 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[931]),
			.N(gen[932]),
			.NE(gen[933]),

			.O(gen[991]),
			.E(gen[993]),

			.SO(gen[1051]),
			.S(gen[1052]),
			.SE(gen[1053]),

			.SELF(gen[992]),
			.cell_state(gen[992])
		); 

/******************* CELL 993 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell993 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[932]),
			.N(gen[933]),
			.NE(gen[934]),

			.O(gen[992]),
			.E(gen[994]),

			.SO(gen[1052]),
			.S(gen[1053]),
			.SE(gen[1054]),

			.SELF(gen[993]),
			.cell_state(gen[993])
		); 

/******************* CELL 994 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell994 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[933]),
			.N(gen[934]),
			.NE(gen[935]),

			.O(gen[993]),
			.E(gen[995]),

			.SO(gen[1053]),
			.S(gen[1054]),
			.SE(gen[1055]),

			.SELF(gen[994]),
			.cell_state(gen[994])
		); 

/******************* CELL 995 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell995 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[934]),
			.N(gen[935]),
			.NE(gen[936]),

			.O(gen[994]),
			.E(gen[996]),

			.SO(gen[1054]),
			.S(gen[1055]),
			.SE(gen[1056]),

			.SELF(gen[995]),
			.cell_state(gen[995])
		); 

/******************* CELL 996 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell996 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[935]),
			.N(gen[936]),
			.NE(gen[937]),

			.O(gen[995]),
			.E(gen[997]),

			.SO(gen[1055]),
			.S(gen[1056]),
			.SE(gen[1057]),

			.SELF(gen[996]),
			.cell_state(gen[996])
		); 

/******************* CELL 997 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell997 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[936]),
			.N(gen[937]),
			.NE(gen[938]),

			.O(gen[996]),
			.E(gen[998]),

			.SO(gen[1056]),
			.S(gen[1057]),
			.SE(gen[1058]),

			.SELF(gen[997]),
			.cell_state(gen[997])
		); 

/******************* CELL 998 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell998 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[937]),
			.N(gen[938]),
			.NE(gen[939]),

			.O(gen[997]),
			.E(gen[999]),

			.SO(gen[1057]),
			.S(gen[1058]),
			.SE(gen[1059]),

			.SELF(gen[998]),
			.cell_state(gen[998])
		); 

/******************* CELL 999 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell999 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[938]),
			.N(gen[939]),
			.NE(gen[940]),

			.O(gen[998]),
			.E(gen[1000]),

			.SO(gen[1058]),
			.S(gen[1059]),
			.SE(gen[1060]),

			.SELF(gen[999]),
			.cell_state(gen[999])
		); 

/******************* CELL 1000 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1000 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[939]),
			.N(gen[940]),
			.NE(gen[941]),

			.O(gen[999]),
			.E(gen[1001]),

			.SO(gen[1059]),
			.S(gen[1060]),
			.SE(gen[1061]),

			.SELF(gen[1000]),
			.cell_state(gen[1000])
		); 

/******************* CELL 1001 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1001 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[940]),
			.N(gen[941]),
			.NE(gen[942]),

			.O(gen[1000]),
			.E(gen[1002]),

			.SO(gen[1060]),
			.S(gen[1061]),
			.SE(gen[1062]),

			.SELF(gen[1001]),
			.cell_state(gen[1001])
		); 

/******************* CELL 1002 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1002 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[941]),
			.N(gen[942]),
			.NE(gen[943]),

			.O(gen[1001]),
			.E(gen[1003]),

			.SO(gen[1061]),
			.S(gen[1062]),
			.SE(gen[1063]),

			.SELF(gen[1002]),
			.cell_state(gen[1002])
		); 

/******************* CELL 1003 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1003 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[942]),
			.N(gen[943]),
			.NE(gen[944]),

			.O(gen[1002]),
			.E(gen[1004]),

			.SO(gen[1062]),
			.S(gen[1063]),
			.SE(gen[1064]),

			.SELF(gen[1003]),
			.cell_state(gen[1003])
		); 

/******************* CELL 1004 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1004 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[943]),
			.N(gen[944]),
			.NE(gen[945]),

			.O(gen[1003]),
			.E(gen[1005]),

			.SO(gen[1063]),
			.S(gen[1064]),
			.SE(gen[1065]),

			.SELF(gen[1004]),
			.cell_state(gen[1004])
		); 

/******************* CELL 1005 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1005 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[944]),
			.N(gen[945]),
			.NE(gen[946]),

			.O(gen[1004]),
			.E(gen[1006]),

			.SO(gen[1064]),
			.S(gen[1065]),
			.SE(gen[1066]),

			.SELF(gen[1005]),
			.cell_state(gen[1005])
		); 

/******************* CELL 1006 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1006 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[945]),
			.N(gen[946]),
			.NE(gen[947]),

			.O(gen[1005]),
			.E(gen[1007]),

			.SO(gen[1065]),
			.S(gen[1066]),
			.SE(gen[1067]),

			.SELF(gen[1006]),
			.cell_state(gen[1006])
		); 

/******************* CELL 1007 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1007 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[946]),
			.N(gen[947]),
			.NE(gen[948]),

			.O(gen[1006]),
			.E(gen[1008]),

			.SO(gen[1066]),
			.S(gen[1067]),
			.SE(gen[1068]),

			.SELF(gen[1007]),
			.cell_state(gen[1007])
		); 

/******************* CELL 1008 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1008 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[947]),
			.N(gen[948]),
			.NE(gen[949]),

			.O(gen[1007]),
			.E(gen[1009]),

			.SO(gen[1067]),
			.S(gen[1068]),
			.SE(gen[1069]),

			.SELF(gen[1008]),
			.cell_state(gen[1008])
		); 

/******************* CELL 1009 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1009 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[948]),
			.N(gen[949]),
			.NE(gen[950]),

			.O(gen[1008]),
			.E(gen[1010]),

			.SO(gen[1068]),
			.S(gen[1069]),
			.SE(gen[1070]),

			.SELF(gen[1009]),
			.cell_state(gen[1009])
		); 

/******************* CELL 1010 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1010 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[949]),
			.N(gen[950]),
			.NE(gen[951]),

			.O(gen[1009]),
			.E(gen[1011]),

			.SO(gen[1069]),
			.S(gen[1070]),
			.SE(gen[1071]),

			.SELF(gen[1010]),
			.cell_state(gen[1010])
		); 

/******************* CELL 1011 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1011 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[950]),
			.N(gen[951]),
			.NE(gen[952]),

			.O(gen[1010]),
			.E(gen[1012]),

			.SO(gen[1070]),
			.S(gen[1071]),
			.SE(gen[1072]),

			.SELF(gen[1011]),
			.cell_state(gen[1011])
		); 

/******************* CELL 1012 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1012 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[951]),
			.N(gen[952]),
			.NE(gen[953]),

			.O(gen[1011]),
			.E(gen[1013]),

			.SO(gen[1071]),
			.S(gen[1072]),
			.SE(gen[1073]),

			.SELF(gen[1012]),
			.cell_state(gen[1012])
		); 

/******************* CELL 1013 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1013 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[952]),
			.N(gen[953]),
			.NE(gen[954]),

			.O(gen[1012]),
			.E(gen[1014]),

			.SO(gen[1072]),
			.S(gen[1073]),
			.SE(gen[1074]),

			.SELF(gen[1013]),
			.cell_state(gen[1013])
		); 

/******************* CELL 1014 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1014 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[953]),
			.N(gen[954]),
			.NE(gen[955]),

			.O(gen[1013]),
			.E(gen[1015]),

			.SO(gen[1073]),
			.S(gen[1074]),
			.SE(gen[1075]),

			.SELF(gen[1014]),
			.cell_state(gen[1014])
		); 

/******************* CELL 1015 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1015 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[954]),
			.N(gen[955]),
			.NE(gen[956]),

			.O(gen[1014]),
			.E(gen[1016]),

			.SO(gen[1074]),
			.S(gen[1075]),
			.SE(gen[1076]),

			.SELF(gen[1015]),
			.cell_state(gen[1015])
		); 

/******************* CELL 1016 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1016 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[955]),
			.N(gen[956]),
			.NE(gen[957]),

			.O(gen[1015]),
			.E(gen[1017]),

			.SO(gen[1075]),
			.S(gen[1076]),
			.SE(gen[1077]),

			.SELF(gen[1016]),
			.cell_state(gen[1016])
		); 

/******************* CELL 1017 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1017 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[956]),
			.N(gen[957]),
			.NE(gen[958]),

			.O(gen[1016]),
			.E(gen[1018]),

			.SO(gen[1076]),
			.S(gen[1077]),
			.SE(gen[1078]),

			.SELF(gen[1017]),
			.cell_state(gen[1017])
		); 

/******************* CELL 1018 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1018 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[957]),
			.N(gen[958]),
			.NE(gen[959]),

			.O(gen[1017]),
			.E(gen[1019]),

			.SO(gen[1077]),
			.S(gen[1078]),
			.SE(gen[1079]),

			.SELF(gen[1018]),
			.cell_state(gen[1018])
		); 

/******************* CELL 1019 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1019 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[958]),
			.N(gen[959]),
			.NE(gen[958]),

			.O(gen[1018]),
			.E(gen[1018]),

			.SO(gen[1078]),
			.S(gen[1079]),
			.SE(gen[1078]),

			.SELF(gen[1019]),
			.cell_state(gen[1019])
		); 

/******************* CELL 1020 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1020 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[961]),
			.N(gen[960]),
			.NE(gen[961]),

			.O(gen[1021]),
			.E(gen[1021]),

			.SO(gen[1081]),
			.S(gen[1080]),
			.SE(gen[1081]),

			.SELF(gen[1020]),
			.cell_state(gen[1020])
		); 

/******************* CELL 1021 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1021 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[960]),
			.N(gen[961]),
			.NE(gen[962]),

			.O(gen[1020]),
			.E(gen[1022]),

			.SO(gen[1080]),
			.S(gen[1081]),
			.SE(gen[1082]),

			.SELF(gen[1021]),
			.cell_state(gen[1021])
		); 

/******************* CELL 1022 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1022 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[961]),
			.N(gen[962]),
			.NE(gen[963]),

			.O(gen[1021]),
			.E(gen[1023]),

			.SO(gen[1081]),
			.S(gen[1082]),
			.SE(gen[1083]),

			.SELF(gen[1022]),
			.cell_state(gen[1022])
		); 

/******************* CELL 1023 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1023 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[962]),
			.N(gen[963]),
			.NE(gen[964]),

			.O(gen[1022]),
			.E(gen[1024]),

			.SO(gen[1082]),
			.S(gen[1083]),
			.SE(gen[1084]),

			.SELF(gen[1023]),
			.cell_state(gen[1023])
		); 

/******************* CELL 1024 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1024 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[963]),
			.N(gen[964]),
			.NE(gen[965]),

			.O(gen[1023]),
			.E(gen[1025]),

			.SO(gen[1083]),
			.S(gen[1084]),
			.SE(gen[1085]),

			.SELF(gen[1024]),
			.cell_state(gen[1024])
		); 

/******************* CELL 1025 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1025 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[964]),
			.N(gen[965]),
			.NE(gen[966]),

			.O(gen[1024]),
			.E(gen[1026]),

			.SO(gen[1084]),
			.S(gen[1085]),
			.SE(gen[1086]),

			.SELF(gen[1025]),
			.cell_state(gen[1025])
		); 

/******************* CELL 1026 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1026 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[965]),
			.N(gen[966]),
			.NE(gen[967]),

			.O(gen[1025]),
			.E(gen[1027]),

			.SO(gen[1085]),
			.S(gen[1086]),
			.SE(gen[1087]),

			.SELF(gen[1026]),
			.cell_state(gen[1026])
		); 

/******************* CELL 1027 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1027 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[966]),
			.N(gen[967]),
			.NE(gen[968]),

			.O(gen[1026]),
			.E(gen[1028]),

			.SO(gen[1086]),
			.S(gen[1087]),
			.SE(gen[1088]),

			.SELF(gen[1027]),
			.cell_state(gen[1027])
		); 

/******************* CELL 1028 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1028 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[967]),
			.N(gen[968]),
			.NE(gen[969]),

			.O(gen[1027]),
			.E(gen[1029]),

			.SO(gen[1087]),
			.S(gen[1088]),
			.SE(gen[1089]),

			.SELF(gen[1028]),
			.cell_state(gen[1028])
		); 

/******************* CELL 1029 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1029 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[968]),
			.N(gen[969]),
			.NE(gen[970]),

			.O(gen[1028]),
			.E(gen[1030]),

			.SO(gen[1088]),
			.S(gen[1089]),
			.SE(gen[1090]),

			.SELF(gen[1029]),
			.cell_state(gen[1029])
		); 

/******************* CELL 1030 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1030 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[969]),
			.N(gen[970]),
			.NE(gen[971]),

			.O(gen[1029]),
			.E(gen[1031]),

			.SO(gen[1089]),
			.S(gen[1090]),
			.SE(gen[1091]),

			.SELF(gen[1030]),
			.cell_state(gen[1030])
		); 

/******************* CELL 1031 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1031 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[970]),
			.N(gen[971]),
			.NE(gen[972]),

			.O(gen[1030]),
			.E(gen[1032]),

			.SO(gen[1090]),
			.S(gen[1091]),
			.SE(gen[1092]),

			.SELF(gen[1031]),
			.cell_state(gen[1031])
		); 

/******************* CELL 1032 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1032 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[971]),
			.N(gen[972]),
			.NE(gen[973]),

			.O(gen[1031]),
			.E(gen[1033]),

			.SO(gen[1091]),
			.S(gen[1092]),
			.SE(gen[1093]),

			.SELF(gen[1032]),
			.cell_state(gen[1032])
		); 

/******************* CELL 1033 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1033 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[972]),
			.N(gen[973]),
			.NE(gen[974]),

			.O(gen[1032]),
			.E(gen[1034]),

			.SO(gen[1092]),
			.S(gen[1093]),
			.SE(gen[1094]),

			.SELF(gen[1033]),
			.cell_state(gen[1033])
		); 

/******************* CELL 1034 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1034 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[973]),
			.N(gen[974]),
			.NE(gen[975]),

			.O(gen[1033]),
			.E(gen[1035]),

			.SO(gen[1093]),
			.S(gen[1094]),
			.SE(gen[1095]),

			.SELF(gen[1034]),
			.cell_state(gen[1034])
		); 

/******************* CELL 1035 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1035 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[974]),
			.N(gen[975]),
			.NE(gen[976]),

			.O(gen[1034]),
			.E(gen[1036]),

			.SO(gen[1094]),
			.S(gen[1095]),
			.SE(gen[1096]),

			.SELF(gen[1035]),
			.cell_state(gen[1035])
		); 

/******************* CELL 1036 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1036 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[975]),
			.N(gen[976]),
			.NE(gen[977]),

			.O(gen[1035]),
			.E(gen[1037]),

			.SO(gen[1095]),
			.S(gen[1096]),
			.SE(gen[1097]),

			.SELF(gen[1036]),
			.cell_state(gen[1036])
		); 

/******************* CELL 1037 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1037 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[976]),
			.N(gen[977]),
			.NE(gen[978]),

			.O(gen[1036]),
			.E(gen[1038]),

			.SO(gen[1096]),
			.S(gen[1097]),
			.SE(gen[1098]),

			.SELF(gen[1037]),
			.cell_state(gen[1037])
		); 

/******************* CELL 1038 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1038 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[977]),
			.N(gen[978]),
			.NE(gen[979]),

			.O(gen[1037]),
			.E(gen[1039]),

			.SO(gen[1097]),
			.S(gen[1098]),
			.SE(gen[1099]),

			.SELF(gen[1038]),
			.cell_state(gen[1038])
		); 

/******************* CELL 1039 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1039 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[978]),
			.N(gen[979]),
			.NE(gen[980]),

			.O(gen[1038]),
			.E(gen[1040]),

			.SO(gen[1098]),
			.S(gen[1099]),
			.SE(gen[1100]),

			.SELF(gen[1039]),
			.cell_state(gen[1039])
		); 

/******************* CELL 1040 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1040 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[979]),
			.N(gen[980]),
			.NE(gen[981]),

			.O(gen[1039]),
			.E(gen[1041]),

			.SO(gen[1099]),
			.S(gen[1100]),
			.SE(gen[1101]),

			.SELF(gen[1040]),
			.cell_state(gen[1040])
		); 

/******************* CELL 1041 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1041 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[980]),
			.N(gen[981]),
			.NE(gen[982]),

			.O(gen[1040]),
			.E(gen[1042]),

			.SO(gen[1100]),
			.S(gen[1101]),
			.SE(gen[1102]),

			.SELF(gen[1041]),
			.cell_state(gen[1041])
		); 

/******************* CELL 1042 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1042 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[981]),
			.N(gen[982]),
			.NE(gen[983]),

			.O(gen[1041]),
			.E(gen[1043]),

			.SO(gen[1101]),
			.S(gen[1102]),
			.SE(gen[1103]),

			.SELF(gen[1042]),
			.cell_state(gen[1042])
		); 

/******************* CELL 1043 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1043 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[982]),
			.N(gen[983]),
			.NE(gen[984]),

			.O(gen[1042]),
			.E(gen[1044]),

			.SO(gen[1102]),
			.S(gen[1103]),
			.SE(gen[1104]),

			.SELF(gen[1043]),
			.cell_state(gen[1043])
		); 

/******************* CELL 1044 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1044 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[983]),
			.N(gen[984]),
			.NE(gen[985]),

			.O(gen[1043]),
			.E(gen[1045]),

			.SO(gen[1103]),
			.S(gen[1104]),
			.SE(gen[1105]),

			.SELF(gen[1044]),
			.cell_state(gen[1044])
		); 

/******************* CELL 1045 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1045 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[984]),
			.N(gen[985]),
			.NE(gen[986]),

			.O(gen[1044]),
			.E(gen[1046]),

			.SO(gen[1104]),
			.S(gen[1105]),
			.SE(gen[1106]),

			.SELF(gen[1045]),
			.cell_state(gen[1045])
		); 

/******************* CELL 1046 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1046 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[985]),
			.N(gen[986]),
			.NE(gen[987]),

			.O(gen[1045]),
			.E(gen[1047]),

			.SO(gen[1105]),
			.S(gen[1106]),
			.SE(gen[1107]),

			.SELF(gen[1046]),
			.cell_state(gen[1046])
		); 

/******************* CELL 1047 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1047 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[986]),
			.N(gen[987]),
			.NE(gen[988]),

			.O(gen[1046]),
			.E(gen[1048]),

			.SO(gen[1106]),
			.S(gen[1107]),
			.SE(gen[1108]),

			.SELF(gen[1047]),
			.cell_state(gen[1047])
		); 

/******************* CELL 1048 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1048 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[987]),
			.N(gen[988]),
			.NE(gen[989]),

			.O(gen[1047]),
			.E(gen[1049]),

			.SO(gen[1107]),
			.S(gen[1108]),
			.SE(gen[1109]),

			.SELF(gen[1048]),
			.cell_state(gen[1048])
		); 

/******************* CELL 1049 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1049 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[988]),
			.N(gen[989]),
			.NE(gen[990]),

			.O(gen[1048]),
			.E(gen[1050]),

			.SO(gen[1108]),
			.S(gen[1109]),
			.SE(gen[1110]),

			.SELF(gen[1049]),
			.cell_state(gen[1049])
		); 

/******************* CELL 1050 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1050 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[989]),
			.N(gen[990]),
			.NE(gen[991]),

			.O(gen[1049]),
			.E(gen[1051]),

			.SO(gen[1109]),
			.S(gen[1110]),
			.SE(gen[1111]),

			.SELF(gen[1050]),
			.cell_state(gen[1050])
		); 

/******************* CELL 1051 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1051 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[990]),
			.N(gen[991]),
			.NE(gen[992]),

			.O(gen[1050]),
			.E(gen[1052]),

			.SO(gen[1110]),
			.S(gen[1111]),
			.SE(gen[1112]),

			.SELF(gen[1051]),
			.cell_state(gen[1051])
		); 

/******************* CELL 1052 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1052 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[991]),
			.N(gen[992]),
			.NE(gen[993]),

			.O(gen[1051]),
			.E(gen[1053]),

			.SO(gen[1111]),
			.S(gen[1112]),
			.SE(gen[1113]),

			.SELF(gen[1052]),
			.cell_state(gen[1052])
		); 

/******************* CELL 1053 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1053 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[992]),
			.N(gen[993]),
			.NE(gen[994]),

			.O(gen[1052]),
			.E(gen[1054]),

			.SO(gen[1112]),
			.S(gen[1113]),
			.SE(gen[1114]),

			.SELF(gen[1053]),
			.cell_state(gen[1053])
		); 

/******************* CELL 1054 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1054 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[993]),
			.N(gen[994]),
			.NE(gen[995]),

			.O(gen[1053]),
			.E(gen[1055]),

			.SO(gen[1113]),
			.S(gen[1114]),
			.SE(gen[1115]),

			.SELF(gen[1054]),
			.cell_state(gen[1054])
		); 

/******************* CELL 1055 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1055 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[994]),
			.N(gen[995]),
			.NE(gen[996]),

			.O(gen[1054]),
			.E(gen[1056]),

			.SO(gen[1114]),
			.S(gen[1115]),
			.SE(gen[1116]),

			.SELF(gen[1055]),
			.cell_state(gen[1055])
		); 

/******************* CELL 1056 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1056 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[995]),
			.N(gen[996]),
			.NE(gen[997]),

			.O(gen[1055]),
			.E(gen[1057]),

			.SO(gen[1115]),
			.S(gen[1116]),
			.SE(gen[1117]),

			.SELF(gen[1056]),
			.cell_state(gen[1056])
		); 

/******************* CELL 1057 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1057 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[996]),
			.N(gen[997]),
			.NE(gen[998]),

			.O(gen[1056]),
			.E(gen[1058]),

			.SO(gen[1116]),
			.S(gen[1117]),
			.SE(gen[1118]),

			.SELF(gen[1057]),
			.cell_state(gen[1057])
		); 

/******************* CELL 1058 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1058 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[997]),
			.N(gen[998]),
			.NE(gen[999]),

			.O(gen[1057]),
			.E(gen[1059]),

			.SO(gen[1117]),
			.S(gen[1118]),
			.SE(gen[1119]),

			.SELF(gen[1058]),
			.cell_state(gen[1058])
		); 

/******************* CELL 1059 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1059 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[998]),
			.N(gen[999]),
			.NE(gen[1000]),

			.O(gen[1058]),
			.E(gen[1060]),

			.SO(gen[1118]),
			.S(gen[1119]),
			.SE(gen[1120]),

			.SELF(gen[1059]),
			.cell_state(gen[1059])
		); 

/******************* CELL 1060 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1060 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[999]),
			.N(gen[1000]),
			.NE(gen[1001]),

			.O(gen[1059]),
			.E(gen[1061]),

			.SO(gen[1119]),
			.S(gen[1120]),
			.SE(gen[1121]),

			.SELF(gen[1060]),
			.cell_state(gen[1060])
		); 

/******************* CELL 1061 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1061 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1000]),
			.N(gen[1001]),
			.NE(gen[1002]),

			.O(gen[1060]),
			.E(gen[1062]),

			.SO(gen[1120]),
			.S(gen[1121]),
			.SE(gen[1122]),

			.SELF(gen[1061]),
			.cell_state(gen[1061])
		); 

/******************* CELL 1062 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1062 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1001]),
			.N(gen[1002]),
			.NE(gen[1003]),

			.O(gen[1061]),
			.E(gen[1063]),

			.SO(gen[1121]),
			.S(gen[1122]),
			.SE(gen[1123]),

			.SELF(gen[1062]),
			.cell_state(gen[1062])
		); 

/******************* CELL 1063 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1063 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1002]),
			.N(gen[1003]),
			.NE(gen[1004]),

			.O(gen[1062]),
			.E(gen[1064]),

			.SO(gen[1122]),
			.S(gen[1123]),
			.SE(gen[1124]),

			.SELF(gen[1063]),
			.cell_state(gen[1063])
		); 

/******************* CELL 1064 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1064 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1003]),
			.N(gen[1004]),
			.NE(gen[1005]),

			.O(gen[1063]),
			.E(gen[1065]),

			.SO(gen[1123]),
			.S(gen[1124]),
			.SE(gen[1125]),

			.SELF(gen[1064]),
			.cell_state(gen[1064])
		); 

/******************* CELL 1065 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1065 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1004]),
			.N(gen[1005]),
			.NE(gen[1006]),

			.O(gen[1064]),
			.E(gen[1066]),

			.SO(gen[1124]),
			.S(gen[1125]),
			.SE(gen[1126]),

			.SELF(gen[1065]),
			.cell_state(gen[1065])
		); 

/******************* CELL 1066 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1066 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1005]),
			.N(gen[1006]),
			.NE(gen[1007]),

			.O(gen[1065]),
			.E(gen[1067]),

			.SO(gen[1125]),
			.S(gen[1126]),
			.SE(gen[1127]),

			.SELF(gen[1066]),
			.cell_state(gen[1066])
		); 

/******************* CELL 1067 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1067 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1006]),
			.N(gen[1007]),
			.NE(gen[1008]),

			.O(gen[1066]),
			.E(gen[1068]),

			.SO(gen[1126]),
			.S(gen[1127]),
			.SE(gen[1128]),

			.SELF(gen[1067]),
			.cell_state(gen[1067])
		); 

/******************* CELL 1068 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1068 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1007]),
			.N(gen[1008]),
			.NE(gen[1009]),

			.O(gen[1067]),
			.E(gen[1069]),

			.SO(gen[1127]),
			.S(gen[1128]),
			.SE(gen[1129]),

			.SELF(gen[1068]),
			.cell_state(gen[1068])
		); 

/******************* CELL 1069 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1069 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1008]),
			.N(gen[1009]),
			.NE(gen[1010]),

			.O(gen[1068]),
			.E(gen[1070]),

			.SO(gen[1128]),
			.S(gen[1129]),
			.SE(gen[1130]),

			.SELF(gen[1069]),
			.cell_state(gen[1069])
		); 

/******************* CELL 1070 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1070 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1009]),
			.N(gen[1010]),
			.NE(gen[1011]),

			.O(gen[1069]),
			.E(gen[1071]),

			.SO(gen[1129]),
			.S(gen[1130]),
			.SE(gen[1131]),

			.SELF(gen[1070]),
			.cell_state(gen[1070])
		); 

/******************* CELL 1071 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1071 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1010]),
			.N(gen[1011]),
			.NE(gen[1012]),

			.O(gen[1070]),
			.E(gen[1072]),

			.SO(gen[1130]),
			.S(gen[1131]),
			.SE(gen[1132]),

			.SELF(gen[1071]),
			.cell_state(gen[1071])
		); 

/******************* CELL 1072 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1072 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1011]),
			.N(gen[1012]),
			.NE(gen[1013]),

			.O(gen[1071]),
			.E(gen[1073]),

			.SO(gen[1131]),
			.S(gen[1132]),
			.SE(gen[1133]),

			.SELF(gen[1072]),
			.cell_state(gen[1072])
		); 

/******************* CELL 1073 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1073 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1012]),
			.N(gen[1013]),
			.NE(gen[1014]),

			.O(gen[1072]),
			.E(gen[1074]),

			.SO(gen[1132]),
			.S(gen[1133]),
			.SE(gen[1134]),

			.SELF(gen[1073]),
			.cell_state(gen[1073])
		); 

/******************* CELL 1074 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1074 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1013]),
			.N(gen[1014]),
			.NE(gen[1015]),

			.O(gen[1073]),
			.E(gen[1075]),

			.SO(gen[1133]),
			.S(gen[1134]),
			.SE(gen[1135]),

			.SELF(gen[1074]),
			.cell_state(gen[1074])
		); 

/******************* CELL 1075 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1075 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1014]),
			.N(gen[1015]),
			.NE(gen[1016]),

			.O(gen[1074]),
			.E(gen[1076]),

			.SO(gen[1134]),
			.S(gen[1135]),
			.SE(gen[1136]),

			.SELF(gen[1075]),
			.cell_state(gen[1075])
		); 

/******************* CELL 1076 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1076 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1015]),
			.N(gen[1016]),
			.NE(gen[1017]),

			.O(gen[1075]),
			.E(gen[1077]),

			.SO(gen[1135]),
			.S(gen[1136]),
			.SE(gen[1137]),

			.SELF(gen[1076]),
			.cell_state(gen[1076])
		); 

/******************* CELL 1077 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1077 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1016]),
			.N(gen[1017]),
			.NE(gen[1018]),

			.O(gen[1076]),
			.E(gen[1078]),

			.SO(gen[1136]),
			.S(gen[1137]),
			.SE(gen[1138]),

			.SELF(gen[1077]),
			.cell_state(gen[1077])
		); 

/******************* CELL 1078 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1078 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1017]),
			.N(gen[1018]),
			.NE(gen[1019]),

			.O(gen[1077]),
			.E(gen[1079]),

			.SO(gen[1137]),
			.S(gen[1138]),
			.SE(gen[1139]),

			.SELF(gen[1078]),
			.cell_state(gen[1078])
		); 

/******************* CELL 1079 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1079 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1018]),
			.N(gen[1019]),
			.NE(gen[1018]),

			.O(gen[1078]),
			.E(gen[1078]),

			.SO(gen[1138]),
			.S(gen[1139]),
			.SE(gen[1138]),

			.SELF(gen[1079]),
			.cell_state(gen[1079])
		); 

/******************* CELL 1080 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1080 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1021]),
			.N(gen[1020]),
			.NE(gen[1021]),

			.O(gen[1081]),
			.E(gen[1081]),

			.SO(gen[1141]),
			.S(gen[1140]),
			.SE(gen[1141]),

			.SELF(gen[1080]),
			.cell_state(gen[1080])
		); 

/******************* CELL 1081 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1081 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1020]),
			.N(gen[1021]),
			.NE(gen[1022]),

			.O(gen[1080]),
			.E(gen[1082]),

			.SO(gen[1140]),
			.S(gen[1141]),
			.SE(gen[1142]),

			.SELF(gen[1081]),
			.cell_state(gen[1081])
		); 

/******************* CELL 1082 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1082 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1021]),
			.N(gen[1022]),
			.NE(gen[1023]),

			.O(gen[1081]),
			.E(gen[1083]),

			.SO(gen[1141]),
			.S(gen[1142]),
			.SE(gen[1143]),

			.SELF(gen[1082]),
			.cell_state(gen[1082])
		); 

/******************* CELL 1083 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1083 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1022]),
			.N(gen[1023]),
			.NE(gen[1024]),

			.O(gen[1082]),
			.E(gen[1084]),

			.SO(gen[1142]),
			.S(gen[1143]),
			.SE(gen[1144]),

			.SELF(gen[1083]),
			.cell_state(gen[1083])
		); 

/******************* CELL 1084 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1084 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1023]),
			.N(gen[1024]),
			.NE(gen[1025]),

			.O(gen[1083]),
			.E(gen[1085]),

			.SO(gen[1143]),
			.S(gen[1144]),
			.SE(gen[1145]),

			.SELF(gen[1084]),
			.cell_state(gen[1084])
		); 

/******************* CELL 1085 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1085 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1024]),
			.N(gen[1025]),
			.NE(gen[1026]),

			.O(gen[1084]),
			.E(gen[1086]),

			.SO(gen[1144]),
			.S(gen[1145]),
			.SE(gen[1146]),

			.SELF(gen[1085]),
			.cell_state(gen[1085])
		); 

/******************* CELL 1086 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1086 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1025]),
			.N(gen[1026]),
			.NE(gen[1027]),

			.O(gen[1085]),
			.E(gen[1087]),

			.SO(gen[1145]),
			.S(gen[1146]),
			.SE(gen[1147]),

			.SELF(gen[1086]),
			.cell_state(gen[1086])
		); 

/******************* CELL 1087 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1087 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1026]),
			.N(gen[1027]),
			.NE(gen[1028]),

			.O(gen[1086]),
			.E(gen[1088]),

			.SO(gen[1146]),
			.S(gen[1147]),
			.SE(gen[1148]),

			.SELF(gen[1087]),
			.cell_state(gen[1087])
		); 

/******************* CELL 1088 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1088 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1027]),
			.N(gen[1028]),
			.NE(gen[1029]),

			.O(gen[1087]),
			.E(gen[1089]),

			.SO(gen[1147]),
			.S(gen[1148]),
			.SE(gen[1149]),

			.SELF(gen[1088]),
			.cell_state(gen[1088])
		); 

/******************* CELL 1089 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1089 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1028]),
			.N(gen[1029]),
			.NE(gen[1030]),

			.O(gen[1088]),
			.E(gen[1090]),

			.SO(gen[1148]),
			.S(gen[1149]),
			.SE(gen[1150]),

			.SELF(gen[1089]),
			.cell_state(gen[1089])
		); 

/******************* CELL 1090 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1090 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1029]),
			.N(gen[1030]),
			.NE(gen[1031]),

			.O(gen[1089]),
			.E(gen[1091]),

			.SO(gen[1149]),
			.S(gen[1150]),
			.SE(gen[1151]),

			.SELF(gen[1090]),
			.cell_state(gen[1090])
		); 

/******************* CELL 1091 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1091 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1030]),
			.N(gen[1031]),
			.NE(gen[1032]),

			.O(gen[1090]),
			.E(gen[1092]),

			.SO(gen[1150]),
			.S(gen[1151]),
			.SE(gen[1152]),

			.SELF(gen[1091]),
			.cell_state(gen[1091])
		); 

/******************* CELL 1092 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1092 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1031]),
			.N(gen[1032]),
			.NE(gen[1033]),

			.O(gen[1091]),
			.E(gen[1093]),

			.SO(gen[1151]),
			.S(gen[1152]),
			.SE(gen[1153]),

			.SELF(gen[1092]),
			.cell_state(gen[1092])
		); 

/******************* CELL 1093 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1093 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1032]),
			.N(gen[1033]),
			.NE(gen[1034]),

			.O(gen[1092]),
			.E(gen[1094]),

			.SO(gen[1152]),
			.S(gen[1153]),
			.SE(gen[1154]),

			.SELF(gen[1093]),
			.cell_state(gen[1093])
		); 

/******************* CELL 1094 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1094 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1033]),
			.N(gen[1034]),
			.NE(gen[1035]),

			.O(gen[1093]),
			.E(gen[1095]),

			.SO(gen[1153]),
			.S(gen[1154]),
			.SE(gen[1155]),

			.SELF(gen[1094]),
			.cell_state(gen[1094])
		); 

/******************* CELL 1095 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1095 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1034]),
			.N(gen[1035]),
			.NE(gen[1036]),

			.O(gen[1094]),
			.E(gen[1096]),

			.SO(gen[1154]),
			.S(gen[1155]),
			.SE(gen[1156]),

			.SELF(gen[1095]),
			.cell_state(gen[1095])
		); 

/******************* CELL 1096 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1096 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1035]),
			.N(gen[1036]),
			.NE(gen[1037]),

			.O(gen[1095]),
			.E(gen[1097]),

			.SO(gen[1155]),
			.S(gen[1156]),
			.SE(gen[1157]),

			.SELF(gen[1096]),
			.cell_state(gen[1096])
		); 

/******************* CELL 1097 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1097 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1036]),
			.N(gen[1037]),
			.NE(gen[1038]),

			.O(gen[1096]),
			.E(gen[1098]),

			.SO(gen[1156]),
			.S(gen[1157]),
			.SE(gen[1158]),

			.SELF(gen[1097]),
			.cell_state(gen[1097])
		); 

/******************* CELL 1098 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1098 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1037]),
			.N(gen[1038]),
			.NE(gen[1039]),

			.O(gen[1097]),
			.E(gen[1099]),

			.SO(gen[1157]),
			.S(gen[1158]),
			.SE(gen[1159]),

			.SELF(gen[1098]),
			.cell_state(gen[1098])
		); 

/******************* CELL 1099 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1099 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1038]),
			.N(gen[1039]),
			.NE(gen[1040]),

			.O(gen[1098]),
			.E(gen[1100]),

			.SO(gen[1158]),
			.S(gen[1159]),
			.SE(gen[1160]),

			.SELF(gen[1099]),
			.cell_state(gen[1099])
		); 

/******************* CELL 1100 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1100 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1039]),
			.N(gen[1040]),
			.NE(gen[1041]),

			.O(gen[1099]),
			.E(gen[1101]),

			.SO(gen[1159]),
			.S(gen[1160]),
			.SE(gen[1161]),

			.SELF(gen[1100]),
			.cell_state(gen[1100])
		); 

/******************* CELL 1101 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1101 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1040]),
			.N(gen[1041]),
			.NE(gen[1042]),

			.O(gen[1100]),
			.E(gen[1102]),

			.SO(gen[1160]),
			.S(gen[1161]),
			.SE(gen[1162]),

			.SELF(gen[1101]),
			.cell_state(gen[1101])
		); 

/******************* CELL 1102 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1102 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1041]),
			.N(gen[1042]),
			.NE(gen[1043]),

			.O(gen[1101]),
			.E(gen[1103]),

			.SO(gen[1161]),
			.S(gen[1162]),
			.SE(gen[1163]),

			.SELF(gen[1102]),
			.cell_state(gen[1102])
		); 

/******************* CELL 1103 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1103 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1042]),
			.N(gen[1043]),
			.NE(gen[1044]),

			.O(gen[1102]),
			.E(gen[1104]),

			.SO(gen[1162]),
			.S(gen[1163]),
			.SE(gen[1164]),

			.SELF(gen[1103]),
			.cell_state(gen[1103])
		); 

/******************* CELL 1104 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1104 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1043]),
			.N(gen[1044]),
			.NE(gen[1045]),

			.O(gen[1103]),
			.E(gen[1105]),

			.SO(gen[1163]),
			.S(gen[1164]),
			.SE(gen[1165]),

			.SELF(gen[1104]),
			.cell_state(gen[1104])
		); 

/******************* CELL 1105 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1105 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1044]),
			.N(gen[1045]),
			.NE(gen[1046]),

			.O(gen[1104]),
			.E(gen[1106]),

			.SO(gen[1164]),
			.S(gen[1165]),
			.SE(gen[1166]),

			.SELF(gen[1105]),
			.cell_state(gen[1105])
		); 

/******************* CELL 1106 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1106 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1045]),
			.N(gen[1046]),
			.NE(gen[1047]),

			.O(gen[1105]),
			.E(gen[1107]),

			.SO(gen[1165]),
			.S(gen[1166]),
			.SE(gen[1167]),

			.SELF(gen[1106]),
			.cell_state(gen[1106])
		); 

/******************* CELL 1107 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1107 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1046]),
			.N(gen[1047]),
			.NE(gen[1048]),

			.O(gen[1106]),
			.E(gen[1108]),

			.SO(gen[1166]),
			.S(gen[1167]),
			.SE(gen[1168]),

			.SELF(gen[1107]),
			.cell_state(gen[1107])
		); 

/******************* CELL 1108 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1108 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1047]),
			.N(gen[1048]),
			.NE(gen[1049]),

			.O(gen[1107]),
			.E(gen[1109]),

			.SO(gen[1167]),
			.S(gen[1168]),
			.SE(gen[1169]),

			.SELF(gen[1108]),
			.cell_state(gen[1108])
		); 

/******************* CELL 1109 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1109 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1048]),
			.N(gen[1049]),
			.NE(gen[1050]),

			.O(gen[1108]),
			.E(gen[1110]),

			.SO(gen[1168]),
			.S(gen[1169]),
			.SE(gen[1170]),

			.SELF(gen[1109]),
			.cell_state(gen[1109])
		); 

/******************* CELL 1110 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1110 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1049]),
			.N(gen[1050]),
			.NE(gen[1051]),

			.O(gen[1109]),
			.E(gen[1111]),

			.SO(gen[1169]),
			.S(gen[1170]),
			.SE(gen[1171]),

			.SELF(gen[1110]),
			.cell_state(gen[1110])
		); 

/******************* CELL 1111 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1111 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1050]),
			.N(gen[1051]),
			.NE(gen[1052]),

			.O(gen[1110]),
			.E(gen[1112]),

			.SO(gen[1170]),
			.S(gen[1171]),
			.SE(gen[1172]),

			.SELF(gen[1111]),
			.cell_state(gen[1111])
		); 

/******************* CELL 1112 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1112 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1051]),
			.N(gen[1052]),
			.NE(gen[1053]),

			.O(gen[1111]),
			.E(gen[1113]),

			.SO(gen[1171]),
			.S(gen[1172]),
			.SE(gen[1173]),

			.SELF(gen[1112]),
			.cell_state(gen[1112])
		); 

/******************* CELL 1113 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1113 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1052]),
			.N(gen[1053]),
			.NE(gen[1054]),

			.O(gen[1112]),
			.E(gen[1114]),

			.SO(gen[1172]),
			.S(gen[1173]),
			.SE(gen[1174]),

			.SELF(gen[1113]),
			.cell_state(gen[1113])
		); 

/******************* CELL 1114 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1114 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1053]),
			.N(gen[1054]),
			.NE(gen[1055]),

			.O(gen[1113]),
			.E(gen[1115]),

			.SO(gen[1173]),
			.S(gen[1174]),
			.SE(gen[1175]),

			.SELF(gen[1114]),
			.cell_state(gen[1114])
		); 

/******************* CELL 1115 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1115 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1054]),
			.N(gen[1055]),
			.NE(gen[1056]),

			.O(gen[1114]),
			.E(gen[1116]),

			.SO(gen[1174]),
			.S(gen[1175]),
			.SE(gen[1176]),

			.SELF(gen[1115]),
			.cell_state(gen[1115])
		); 

/******************* CELL 1116 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1116 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1055]),
			.N(gen[1056]),
			.NE(gen[1057]),

			.O(gen[1115]),
			.E(gen[1117]),

			.SO(gen[1175]),
			.S(gen[1176]),
			.SE(gen[1177]),

			.SELF(gen[1116]),
			.cell_state(gen[1116])
		); 

/******************* CELL 1117 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1117 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1056]),
			.N(gen[1057]),
			.NE(gen[1058]),

			.O(gen[1116]),
			.E(gen[1118]),

			.SO(gen[1176]),
			.S(gen[1177]),
			.SE(gen[1178]),

			.SELF(gen[1117]),
			.cell_state(gen[1117])
		); 

/******************* CELL 1118 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1118 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1057]),
			.N(gen[1058]),
			.NE(gen[1059]),

			.O(gen[1117]),
			.E(gen[1119]),

			.SO(gen[1177]),
			.S(gen[1178]),
			.SE(gen[1179]),

			.SELF(gen[1118]),
			.cell_state(gen[1118])
		); 

/******************* CELL 1119 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1119 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1058]),
			.N(gen[1059]),
			.NE(gen[1060]),

			.O(gen[1118]),
			.E(gen[1120]),

			.SO(gen[1178]),
			.S(gen[1179]),
			.SE(gen[1180]),

			.SELF(gen[1119]),
			.cell_state(gen[1119])
		); 

/******************* CELL 1120 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1120 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1059]),
			.N(gen[1060]),
			.NE(gen[1061]),

			.O(gen[1119]),
			.E(gen[1121]),

			.SO(gen[1179]),
			.S(gen[1180]),
			.SE(gen[1181]),

			.SELF(gen[1120]),
			.cell_state(gen[1120])
		); 

/******************* CELL 1121 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1121 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1060]),
			.N(gen[1061]),
			.NE(gen[1062]),

			.O(gen[1120]),
			.E(gen[1122]),

			.SO(gen[1180]),
			.S(gen[1181]),
			.SE(gen[1182]),

			.SELF(gen[1121]),
			.cell_state(gen[1121])
		); 

/******************* CELL 1122 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1122 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1061]),
			.N(gen[1062]),
			.NE(gen[1063]),

			.O(gen[1121]),
			.E(gen[1123]),

			.SO(gen[1181]),
			.S(gen[1182]),
			.SE(gen[1183]),

			.SELF(gen[1122]),
			.cell_state(gen[1122])
		); 

/******************* CELL 1123 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1123 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1062]),
			.N(gen[1063]),
			.NE(gen[1064]),

			.O(gen[1122]),
			.E(gen[1124]),

			.SO(gen[1182]),
			.S(gen[1183]),
			.SE(gen[1184]),

			.SELF(gen[1123]),
			.cell_state(gen[1123])
		); 

/******************* CELL 1124 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1124 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1063]),
			.N(gen[1064]),
			.NE(gen[1065]),

			.O(gen[1123]),
			.E(gen[1125]),

			.SO(gen[1183]),
			.S(gen[1184]),
			.SE(gen[1185]),

			.SELF(gen[1124]),
			.cell_state(gen[1124])
		); 

/******************* CELL 1125 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1125 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1064]),
			.N(gen[1065]),
			.NE(gen[1066]),

			.O(gen[1124]),
			.E(gen[1126]),

			.SO(gen[1184]),
			.S(gen[1185]),
			.SE(gen[1186]),

			.SELF(gen[1125]),
			.cell_state(gen[1125])
		); 

/******************* CELL 1126 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1126 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1065]),
			.N(gen[1066]),
			.NE(gen[1067]),

			.O(gen[1125]),
			.E(gen[1127]),

			.SO(gen[1185]),
			.S(gen[1186]),
			.SE(gen[1187]),

			.SELF(gen[1126]),
			.cell_state(gen[1126])
		); 

/******************* CELL 1127 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1127 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1066]),
			.N(gen[1067]),
			.NE(gen[1068]),

			.O(gen[1126]),
			.E(gen[1128]),

			.SO(gen[1186]),
			.S(gen[1187]),
			.SE(gen[1188]),

			.SELF(gen[1127]),
			.cell_state(gen[1127])
		); 

/******************* CELL 1128 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1128 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1067]),
			.N(gen[1068]),
			.NE(gen[1069]),

			.O(gen[1127]),
			.E(gen[1129]),

			.SO(gen[1187]),
			.S(gen[1188]),
			.SE(gen[1189]),

			.SELF(gen[1128]),
			.cell_state(gen[1128])
		); 

/******************* CELL 1129 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1129 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1068]),
			.N(gen[1069]),
			.NE(gen[1070]),

			.O(gen[1128]),
			.E(gen[1130]),

			.SO(gen[1188]),
			.S(gen[1189]),
			.SE(gen[1190]),

			.SELF(gen[1129]),
			.cell_state(gen[1129])
		); 

/******************* CELL 1130 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1130 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1069]),
			.N(gen[1070]),
			.NE(gen[1071]),

			.O(gen[1129]),
			.E(gen[1131]),

			.SO(gen[1189]),
			.S(gen[1190]),
			.SE(gen[1191]),

			.SELF(gen[1130]),
			.cell_state(gen[1130])
		); 

/******************* CELL 1131 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1131 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1070]),
			.N(gen[1071]),
			.NE(gen[1072]),

			.O(gen[1130]),
			.E(gen[1132]),

			.SO(gen[1190]),
			.S(gen[1191]),
			.SE(gen[1192]),

			.SELF(gen[1131]),
			.cell_state(gen[1131])
		); 

/******************* CELL 1132 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1132 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1071]),
			.N(gen[1072]),
			.NE(gen[1073]),

			.O(gen[1131]),
			.E(gen[1133]),

			.SO(gen[1191]),
			.S(gen[1192]),
			.SE(gen[1193]),

			.SELF(gen[1132]),
			.cell_state(gen[1132])
		); 

/******************* CELL 1133 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1133 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1072]),
			.N(gen[1073]),
			.NE(gen[1074]),

			.O(gen[1132]),
			.E(gen[1134]),

			.SO(gen[1192]),
			.S(gen[1193]),
			.SE(gen[1194]),

			.SELF(gen[1133]),
			.cell_state(gen[1133])
		); 

/******************* CELL 1134 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1134 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1073]),
			.N(gen[1074]),
			.NE(gen[1075]),

			.O(gen[1133]),
			.E(gen[1135]),

			.SO(gen[1193]),
			.S(gen[1194]),
			.SE(gen[1195]),

			.SELF(gen[1134]),
			.cell_state(gen[1134])
		); 

/******************* CELL 1135 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1135 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1074]),
			.N(gen[1075]),
			.NE(gen[1076]),

			.O(gen[1134]),
			.E(gen[1136]),

			.SO(gen[1194]),
			.S(gen[1195]),
			.SE(gen[1196]),

			.SELF(gen[1135]),
			.cell_state(gen[1135])
		); 

/******************* CELL 1136 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1136 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1075]),
			.N(gen[1076]),
			.NE(gen[1077]),

			.O(gen[1135]),
			.E(gen[1137]),

			.SO(gen[1195]),
			.S(gen[1196]),
			.SE(gen[1197]),

			.SELF(gen[1136]),
			.cell_state(gen[1136])
		); 

/******************* CELL 1137 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1137 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1076]),
			.N(gen[1077]),
			.NE(gen[1078]),

			.O(gen[1136]),
			.E(gen[1138]),

			.SO(gen[1196]),
			.S(gen[1197]),
			.SE(gen[1198]),

			.SELF(gen[1137]),
			.cell_state(gen[1137])
		); 

/******************* CELL 1138 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1138 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1077]),
			.N(gen[1078]),
			.NE(gen[1079]),

			.O(gen[1137]),
			.E(gen[1139]),

			.SO(gen[1197]),
			.S(gen[1198]),
			.SE(gen[1199]),

			.SELF(gen[1138]),
			.cell_state(gen[1138])
		); 

/******************* CELL 1139 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1139 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1078]),
			.N(gen[1079]),
			.NE(gen[1078]),

			.O(gen[1138]),
			.E(gen[1138]),

			.SO(gen[1198]),
			.S(gen[1199]),
			.SE(gen[1198]),

			.SELF(gen[1139]),
			.cell_state(gen[1139])
		); 

/******************* CELL 1140 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1140 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1081]),
			.N(gen[1080]),
			.NE(gen[1081]),

			.O(gen[1141]),
			.E(gen[1141]),

			.SO(gen[1201]),
			.S(gen[1200]),
			.SE(gen[1201]),

			.SELF(gen[1140]),
			.cell_state(gen[1140])
		); 

/******************* CELL 1141 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1141 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1080]),
			.N(gen[1081]),
			.NE(gen[1082]),

			.O(gen[1140]),
			.E(gen[1142]),

			.SO(gen[1200]),
			.S(gen[1201]),
			.SE(gen[1202]),

			.SELF(gen[1141]),
			.cell_state(gen[1141])
		); 

/******************* CELL 1142 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1142 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1081]),
			.N(gen[1082]),
			.NE(gen[1083]),

			.O(gen[1141]),
			.E(gen[1143]),

			.SO(gen[1201]),
			.S(gen[1202]),
			.SE(gen[1203]),

			.SELF(gen[1142]),
			.cell_state(gen[1142])
		); 

/******************* CELL 1143 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1143 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1082]),
			.N(gen[1083]),
			.NE(gen[1084]),

			.O(gen[1142]),
			.E(gen[1144]),

			.SO(gen[1202]),
			.S(gen[1203]),
			.SE(gen[1204]),

			.SELF(gen[1143]),
			.cell_state(gen[1143])
		); 

/******************* CELL 1144 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1144 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1083]),
			.N(gen[1084]),
			.NE(gen[1085]),

			.O(gen[1143]),
			.E(gen[1145]),

			.SO(gen[1203]),
			.S(gen[1204]),
			.SE(gen[1205]),

			.SELF(gen[1144]),
			.cell_state(gen[1144])
		); 

/******************* CELL 1145 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1145 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1084]),
			.N(gen[1085]),
			.NE(gen[1086]),

			.O(gen[1144]),
			.E(gen[1146]),

			.SO(gen[1204]),
			.S(gen[1205]),
			.SE(gen[1206]),

			.SELF(gen[1145]),
			.cell_state(gen[1145])
		); 

/******************* CELL 1146 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1146 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1085]),
			.N(gen[1086]),
			.NE(gen[1087]),

			.O(gen[1145]),
			.E(gen[1147]),

			.SO(gen[1205]),
			.S(gen[1206]),
			.SE(gen[1207]),

			.SELF(gen[1146]),
			.cell_state(gen[1146])
		); 

/******************* CELL 1147 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1147 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1086]),
			.N(gen[1087]),
			.NE(gen[1088]),

			.O(gen[1146]),
			.E(gen[1148]),

			.SO(gen[1206]),
			.S(gen[1207]),
			.SE(gen[1208]),

			.SELF(gen[1147]),
			.cell_state(gen[1147])
		); 

/******************* CELL 1148 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1148 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1087]),
			.N(gen[1088]),
			.NE(gen[1089]),

			.O(gen[1147]),
			.E(gen[1149]),

			.SO(gen[1207]),
			.S(gen[1208]),
			.SE(gen[1209]),

			.SELF(gen[1148]),
			.cell_state(gen[1148])
		); 

/******************* CELL 1149 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1149 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1088]),
			.N(gen[1089]),
			.NE(gen[1090]),

			.O(gen[1148]),
			.E(gen[1150]),

			.SO(gen[1208]),
			.S(gen[1209]),
			.SE(gen[1210]),

			.SELF(gen[1149]),
			.cell_state(gen[1149])
		); 

/******************* CELL 1150 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1150 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1089]),
			.N(gen[1090]),
			.NE(gen[1091]),

			.O(gen[1149]),
			.E(gen[1151]),

			.SO(gen[1209]),
			.S(gen[1210]),
			.SE(gen[1211]),

			.SELF(gen[1150]),
			.cell_state(gen[1150])
		); 

/******************* CELL 1151 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1151 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1090]),
			.N(gen[1091]),
			.NE(gen[1092]),

			.O(gen[1150]),
			.E(gen[1152]),

			.SO(gen[1210]),
			.S(gen[1211]),
			.SE(gen[1212]),

			.SELF(gen[1151]),
			.cell_state(gen[1151])
		); 

/******************* CELL 1152 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1152 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1091]),
			.N(gen[1092]),
			.NE(gen[1093]),

			.O(gen[1151]),
			.E(gen[1153]),

			.SO(gen[1211]),
			.S(gen[1212]),
			.SE(gen[1213]),

			.SELF(gen[1152]),
			.cell_state(gen[1152])
		); 

/******************* CELL 1153 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1153 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1092]),
			.N(gen[1093]),
			.NE(gen[1094]),

			.O(gen[1152]),
			.E(gen[1154]),

			.SO(gen[1212]),
			.S(gen[1213]),
			.SE(gen[1214]),

			.SELF(gen[1153]),
			.cell_state(gen[1153])
		); 

/******************* CELL 1154 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1154 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1093]),
			.N(gen[1094]),
			.NE(gen[1095]),

			.O(gen[1153]),
			.E(gen[1155]),

			.SO(gen[1213]),
			.S(gen[1214]),
			.SE(gen[1215]),

			.SELF(gen[1154]),
			.cell_state(gen[1154])
		); 

/******************* CELL 1155 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1155 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1094]),
			.N(gen[1095]),
			.NE(gen[1096]),

			.O(gen[1154]),
			.E(gen[1156]),

			.SO(gen[1214]),
			.S(gen[1215]),
			.SE(gen[1216]),

			.SELF(gen[1155]),
			.cell_state(gen[1155])
		); 

/******************* CELL 1156 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1156 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1095]),
			.N(gen[1096]),
			.NE(gen[1097]),

			.O(gen[1155]),
			.E(gen[1157]),

			.SO(gen[1215]),
			.S(gen[1216]),
			.SE(gen[1217]),

			.SELF(gen[1156]),
			.cell_state(gen[1156])
		); 

/******************* CELL 1157 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1157 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1096]),
			.N(gen[1097]),
			.NE(gen[1098]),

			.O(gen[1156]),
			.E(gen[1158]),

			.SO(gen[1216]),
			.S(gen[1217]),
			.SE(gen[1218]),

			.SELF(gen[1157]),
			.cell_state(gen[1157])
		); 

/******************* CELL 1158 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1158 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1097]),
			.N(gen[1098]),
			.NE(gen[1099]),

			.O(gen[1157]),
			.E(gen[1159]),

			.SO(gen[1217]),
			.S(gen[1218]),
			.SE(gen[1219]),

			.SELF(gen[1158]),
			.cell_state(gen[1158])
		); 

/******************* CELL 1159 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1159 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1098]),
			.N(gen[1099]),
			.NE(gen[1100]),

			.O(gen[1158]),
			.E(gen[1160]),

			.SO(gen[1218]),
			.S(gen[1219]),
			.SE(gen[1220]),

			.SELF(gen[1159]),
			.cell_state(gen[1159])
		); 

/******************* CELL 1160 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1160 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1099]),
			.N(gen[1100]),
			.NE(gen[1101]),

			.O(gen[1159]),
			.E(gen[1161]),

			.SO(gen[1219]),
			.S(gen[1220]),
			.SE(gen[1221]),

			.SELF(gen[1160]),
			.cell_state(gen[1160])
		); 

/******************* CELL 1161 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1161 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1100]),
			.N(gen[1101]),
			.NE(gen[1102]),

			.O(gen[1160]),
			.E(gen[1162]),

			.SO(gen[1220]),
			.S(gen[1221]),
			.SE(gen[1222]),

			.SELF(gen[1161]),
			.cell_state(gen[1161])
		); 

/******************* CELL 1162 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1162 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1101]),
			.N(gen[1102]),
			.NE(gen[1103]),

			.O(gen[1161]),
			.E(gen[1163]),

			.SO(gen[1221]),
			.S(gen[1222]),
			.SE(gen[1223]),

			.SELF(gen[1162]),
			.cell_state(gen[1162])
		); 

/******************* CELL 1163 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1163 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1102]),
			.N(gen[1103]),
			.NE(gen[1104]),

			.O(gen[1162]),
			.E(gen[1164]),

			.SO(gen[1222]),
			.S(gen[1223]),
			.SE(gen[1224]),

			.SELF(gen[1163]),
			.cell_state(gen[1163])
		); 

/******************* CELL 1164 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1164 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1103]),
			.N(gen[1104]),
			.NE(gen[1105]),

			.O(gen[1163]),
			.E(gen[1165]),

			.SO(gen[1223]),
			.S(gen[1224]),
			.SE(gen[1225]),

			.SELF(gen[1164]),
			.cell_state(gen[1164])
		); 

/******************* CELL 1165 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1165 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1104]),
			.N(gen[1105]),
			.NE(gen[1106]),

			.O(gen[1164]),
			.E(gen[1166]),

			.SO(gen[1224]),
			.S(gen[1225]),
			.SE(gen[1226]),

			.SELF(gen[1165]),
			.cell_state(gen[1165])
		); 

/******************* CELL 1166 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1166 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1105]),
			.N(gen[1106]),
			.NE(gen[1107]),

			.O(gen[1165]),
			.E(gen[1167]),

			.SO(gen[1225]),
			.S(gen[1226]),
			.SE(gen[1227]),

			.SELF(gen[1166]),
			.cell_state(gen[1166])
		); 

/******************* CELL 1167 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1167 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1106]),
			.N(gen[1107]),
			.NE(gen[1108]),

			.O(gen[1166]),
			.E(gen[1168]),

			.SO(gen[1226]),
			.S(gen[1227]),
			.SE(gen[1228]),

			.SELF(gen[1167]),
			.cell_state(gen[1167])
		); 

/******************* CELL 1168 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1168 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1107]),
			.N(gen[1108]),
			.NE(gen[1109]),

			.O(gen[1167]),
			.E(gen[1169]),

			.SO(gen[1227]),
			.S(gen[1228]),
			.SE(gen[1229]),

			.SELF(gen[1168]),
			.cell_state(gen[1168])
		); 

/******************* CELL 1169 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1169 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1108]),
			.N(gen[1109]),
			.NE(gen[1110]),

			.O(gen[1168]),
			.E(gen[1170]),

			.SO(gen[1228]),
			.S(gen[1229]),
			.SE(gen[1230]),

			.SELF(gen[1169]),
			.cell_state(gen[1169])
		); 

/******************* CELL 1170 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1170 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1109]),
			.N(gen[1110]),
			.NE(gen[1111]),

			.O(gen[1169]),
			.E(gen[1171]),

			.SO(gen[1229]),
			.S(gen[1230]),
			.SE(gen[1231]),

			.SELF(gen[1170]),
			.cell_state(gen[1170])
		); 

/******************* CELL 1171 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1171 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1110]),
			.N(gen[1111]),
			.NE(gen[1112]),

			.O(gen[1170]),
			.E(gen[1172]),

			.SO(gen[1230]),
			.S(gen[1231]),
			.SE(gen[1232]),

			.SELF(gen[1171]),
			.cell_state(gen[1171])
		); 

/******************* CELL 1172 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1172 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1111]),
			.N(gen[1112]),
			.NE(gen[1113]),

			.O(gen[1171]),
			.E(gen[1173]),

			.SO(gen[1231]),
			.S(gen[1232]),
			.SE(gen[1233]),

			.SELF(gen[1172]),
			.cell_state(gen[1172])
		); 

/******************* CELL 1173 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1173 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1112]),
			.N(gen[1113]),
			.NE(gen[1114]),

			.O(gen[1172]),
			.E(gen[1174]),

			.SO(gen[1232]),
			.S(gen[1233]),
			.SE(gen[1234]),

			.SELF(gen[1173]),
			.cell_state(gen[1173])
		); 

/******************* CELL 1174 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1174 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1113]),
			.N(gen[1114]),
			.NE(gen[1115]),

			.O(gen[1173]),
			.E(gen[1175]),

			.SO(gen[1233]),
			.S(gen[1234]),
			.SE(gen[1235]),

			.SELF(gen[1174]),
			.cell_state(gen[1174])
		); 

/******************* CELL 1175 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1175 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1114]),
			.N(gen[1115]),
			.NE(gen[1116]),

			.O(gen[1174]),
			.E(gen[1176]),

			.SO(gen[1234]),
			.S(gen[1235]),
			.SE(gen[1236]),

			.SELF(gen[1175]),
			.cell_state(gen[1175])
		); 

/******************* CELL 1176 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1176 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1115]),
			.N(gen[1116]),
			.NE(gen[1117]),

			.O(gen[1175]),
			.E(gen[1177]),

			.SO(gen[1235]),
			.S(gen[1236]),
			.SE(gen[1237]),

			.SELF(gen[1176]),
			.cell_state(gen[1176])
		); 

/******************* CELL 1177 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1177 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1116]),
			.N(gen[1117]),
			.NE(gen[1118]),

			.O(gen[1176]),
			.E(gen[1178]),

			.SO(gen[1236]),
			.S(gen[1237]),
			.SE(gen[1238]),

			.SELF(gen[1177]),
			.cell_state(gen[1177])
		); 

/******************* CELL 1178 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1178 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1117]),
			.N(gen[1118]),
			.NE(gen[1119]),

			.O(gen[1177]),
			.E(gen[1179]),

			.SO(gen[1237]),
			.S(gen[1238]),
			.SE(gen[1239]),

			.SELF(gen[1178]),
			.cell_state(gen[1178])
		); 

/******************* CELL 1179 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1179 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1118]),
			.N(gen[1119]),
			.NE(gen[1120]),

			.O(gen[1178]),
			.E(gen[1180]),

			.SO(gen[1238]),
			.S(gen[1239]),
			.SE(gen[1240]),

			.SELF(gen[1179]),
			.cell_state(gen[1179])
		); 

/******************* CELL 1180 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1180 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1119]),
			.N(gen[1120]),
			.NE(gen[1121]),

			.O(gen[1179]),
			.E(gen[1181]),

			.SO(gen[1239]),
			.S(gen[1240]),
			.SE(gen[1241]),

			.SELF(gen[1180]),
			.cell_state(gen[1180])
		); 

/******************* CELL 1181 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1181 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1120]),
			.N(gen[1121]),
			.NE(gen[1122]),

			.O(gen[1180]),
			.E(gen[1182]),

			.SO(gen[1240]),
			.S(gen[1241]),
			.SE(gen[1242]),

			.SELF(gen[1181]),
			.cell_state(gen[1181])
		); 

/******************* CELL 1182 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1182 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1121]),
			.N(gen[1122]),
			.NE(gen[1123]),

			.O(gen[1181]),
			.E(gen[1183]),

			.SO(gen[1241]),
			.S(gen[1242]),
			.SE(gen[1243]),

			.SELF(gen[1182]),
			.cell_state(gen[1182])
		); 

/******************* CELL 1183 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1183 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1122]),
			.N(gen[1123]),
			.NE(gen[1124]),

			.O(gen[1182]),
			.E(gen[1184]),

			.SO(gen[1242]),
			.S(gen[1243]),
			.SE(gen[1244]),

			.SELF(gen[1183]),
			.cell_state(gen[1183])
		); 

/******************* CELL 1184 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1184 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1123]),
			.N(gen[1124]),
			.NE(gen[1125]),

			.O(gen[1183]),
			.E(gen[1185]),

			.SO(gen[1243]),
			.S(gen[1244]),
			.SE(gen[1245]),

			.SELF(gen[1184]),
			.cell_state(gen[1184])
		); 

/******************* CELL 1185 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1185 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1124]),
			.N(gen[1125]),
			.NE(gen[1126]),

			.O(gen[1184]),
			.E(gen[1186]),

			.SO(gen[1244]),
			.S(gen[1245]),
			.SE(gen[1246]),

			.SELF(gen[1185]),
			.cell_state(gen[1185])
		); 

/******************* CELL 1186 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1186 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1125]),
			.N(gen[1126]),
			.NE(gen[1127]),

			.O(gen[1185]),
			.E(gen[1187]),

			.SO(gen[1245]),
			.S(gen[1246]),
			.SE(gen[1247]),

			.SELF(gen[1186]),
			.cell_state(gen[1186])
		); 

/******************* CELL 1187 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1187 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1126]),
			.N(gen[1127]),
			.NE(gen[1128]),

			.O(gen[1186]),
			.E(gen[1188]),

			.SO(gen[1246]),
			.S(gen[1247]),
			.SE(gen[1248]),

			.SELF(gen[1187]),
			.cell_state(gen[1187])
		); 

/******************* CELL 1188 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1188 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1127]),
			.N(gen[1128]),
			.NE(gen[1129]),

			.O(gen[1187]),
			.E(gen[1189]),

			.SO(gen[1247]),
			.S(gen[1248]),
			.SE(gen[1249]),

			.SELF(gen[1188]),
			.cell_state(gen[1188])
		); 

/******************* CELL 1189 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1189 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1128]),
			.N(gen[1129]),
			.NE(gen[1130]),

			.O(gen[1188]),
			.E(gen[1190]),

			.SO(gen[1248]),
			.S(gen[1249]),
			.SE(gen[1250]),

			.SELF(gen[1189]),
			.cell_state(gen[1189])
		); 

/******************* CELL 1190 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1190 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1129]),
			.N(gen[1130]),
			.NE(gen[1131]),

			.O(gen[1189]),
			.E(gen[1191]),

			.SO(gen[1249]),
			.S(gen[1250]),
			.SE(gen[1251]),

			.SELF(gen[1190]),
			.cell_state(gen[1190])
		); 

/******************* CELL 1191 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1191 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1130]),
			.N(gen[1131]),
			.NE(gen[1132]),

			.O(gen[1190]),
			.E(gen[1192]),

			.SO(gen[1250]),
			.S(gen[1251]),
			.SE(gen[1252]),

			.SELF(gen[1191]),
			.cell_state(gen[1191])
		); 

/******************* CELL 1192 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1192 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1131]),
			.N(gen[1132]),
			.NE(gen[1133]),

			.O(gen[1191]),
			.E(gen[1193]),

			.SO(gen[1251]),
			.S(gen[1252]),
			.SE(gen[1253]),

			.SELF(gen[1192]),
			.cell_state(gen[1192])
		); 

/******************* CELL 1193 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1193 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1132]),
			.N(gen[1133]),
			.NE(gen[1134]),

			.O(gen[1192]),
			.E(gen[1194]),

			.SO(gen[1252]),
			.S(gen[1253]),
			.SE(gen[1254]),

			.SELF(gen[1193]),
			.cell_state(gen[1193])
		); 

/******************* CELL 1194 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1194 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1133]),
			.N(gen[1134]),
			.NE(gen[1135]),

			.O(gen[1193]),
			.E(gen[1195]),

			.SO(gen[1253]),
			.S(gen[1254]),
			.SE(gen[1255]),

			.SELF(gen[1194]),
			.cell_state(gen[1194])
		); 

/******************* CELL 1195 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1195 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1134]),
			.N(gen[1135]),
			.NE(gen[1136]),

			.O(gen[1194]),
			.E(gen[1196]),

			.SO(gen[1254]),
			.S(gen[1255]),
			.SE(gen[1256]),

			.SELF(gen[1195]),
			.cell_state(gen[1195])
		); 

/******************* CELL 1196 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1196 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1135]),
			.N(gen[1136]),
			.NE(gen[1137]),

			.O(gen[1195]),
			.E(gen[1197]),

			.SO(gen[1255]),
			.S(gen[1256]),
			.SE(gen[1257]),

			.SELF(gen[1196]),
			.cell_state(gen[1196])
		); 

/******************* CELL 1197 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1197 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1136]),
			.N(gen[1137]),
			.NE(gen[1138]),

			.O(gen[1196]),
			.E(gen[1198]),

			.SO(gen[1256]),
			.S(gen[1257]),
			.SE(gen[1258]),

			.SELF(gen[1197]),
			.cell_state(gen[1197])
		); 

/******************* CELL 1198 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1198 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1137]),
			.N(gen[1138]),
			.NE(gen[1139]),

			.O(gen[1197]),
			.E(gen[1199]),

			.SO(gen[1257]),
			.S(gen[1258]),
			.SE(gen[1259]),

			.SELF(gen[1198]),
			.cell_state(gen[1198])
		); 

/******************* CELL 1199 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1199 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1138]),
			.N(gen[1139]),
			.NE(gen[1138]),

			.O(gen[1198]),
			.E(gen[1198]),

			.SO(gen[1258]),
			.S(gen[1259]),
			.SE(gen[1258]),

			.SELF(gen[1199]),
			.cell_state(gen[1199])
		); 

/******************* CELL 1200 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1200 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1141]),
			.N(gen[1140]),
			.NE(gen[1141]),

			.O(gen[1201]),
			.E(gen[1201]),

			.SO(gen[1261]),
			.S(gen[1260]),
			.SE(gen[1261]),

			.SELF(gen[1200]),
			.cell_state(gen[1200])
		); 

/******************* CELL 1201 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1201 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1140]),
			.N(gen[1141]),
			.NE(gen[1142]),

			.O(gen[1200]),
			.E(gen[1202]),

			.SO(gen[1260]),
			.S(gen[1261]),
			.SE(gen[1262]),

			.SELF(gen[1201]),
			.cell_state(gen[1201])
		); 

/******************* CELL 1202 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1202 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1141]),
			.N(gen[1142]),
			.NE(gen[1143]),

			.O(gen[1201]),
			.E(gen[1203]),

			.SO(gen[1261]),
			.S(gen[1262]),
			.SE(gen[1263]),

			.SELF(gen[1202]),
			.cell_state(gen[1202])
		); 

/******************* CELL 1203 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1203 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1142]),
			.N(gen[1143]),
			.NE(gen[1144]),

			.O(gen[1202]),
			.E(gen[1204]),

			.SO(gen[1262]),
			.S(gen[1263]),
			.SE(gen[1264]),

			.SELF(gen[1203]),
			.cell_state(gen[1203])
		); 

/******************* CELL 1204 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1204 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1143]),
			.N(gen[1144]),
			.NE(gen[1145]),

			.O(gen[1203]),
			.E(gen[1205]),

			.SO(gen[1263]),
			.S(gen[1264]),
			.SE(gen[1265]),

			.SELF(gen[1204]),
			.cell_state(gen[1204])
		); 

/******************* CELL 1205 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1205 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1144]),
			.N(gen[1145]),
			.NE(gen[1146]),

			.O(gen[1204]),
			.E(gen[1206]),

			.SO(gen[1264]),
			.S(gen[1265]),
			.SE(gen[1266]),

			.SELF(gen[1205]),
			.cell_state(gen[1205])
		); 

/******************* CELL 1206 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1206 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1145]),
			.N(gen[1146]),
			.NE(gen[1147]),

			.O(gen[1205]),
			.E(gen[1207]),

			.SO(gen[1265]),
			.S(gen[1266]),
			.SE(gen[1267]),

			.SELF(gen[1206]),
			.cell_state(gen[1206])
		); 

/******************* CELL 1207 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1207 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1146]),
			.N(gen[1147]),
			.NE(gen[1148]),

			.O(gen[1206]),
			.E(gen[1208]),

			.SO(gen[1266]),
			.S(gen[1267]),
			.SE(gen[1268]),

			.SELF(gen[1207]),
			.cell_state(gen[1207])
		); 

/******************* CELL 1208 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1208 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1147]),
			.N(gen[1148]),
			.NE(gen[1149]),

			.O(gen[1207]),
			.E(gen[1209]),

			.SO(gen[1267]),
			.S(gen[1268]),
			.SE(gen[1269]),

			.SELF(gen[1208]),
			.cell_state(gen[1208])
		); 

/******************* CELL 1209 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1209 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1148]),
			.N(gen[1149]),
			.NE(gen[1150]),

			.O(gen[1208]),
			.E(gen[1210]),

			.SO(gen[1268]),
			.S(gen[1269]),
			.SE(gen[1270]),

			.SELF(gen[1209]),
			.cell_state(gen[1209])
		); 

/******************* CELL 1210 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1210 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1149]),
			.N(gen[1150]),
			.NE(gen[1151]),

			.O(gen[1209]),
			.E(gen[1211]),

			.SO(gen[1269]),
			.S(gen[1270]),
			.SE(gen[1271]),

			.SELF(gen[1210]),
			.cell_state(gen[1210])
		); 

/******************* CELL 1211 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1211 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1150]),
			.N(gen[1151]),
			.NE(gen[1152]),

			.O(gen[1210]),
			.E(gen[1212]),

			.SO(gen[1270]),
			.S(gen[1271]),
			.SE(gen[1272]),

			.SELF(gen[1211]),
			.cell_state(gen[1211])
		); 

/******************* CELL 1212 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1212 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1151]),
			.N(gen[1152]),
			.NE(gen[1153]),

			.O(gen[1211]),
			.E(gen[1213]),

			.SO(gen[1271]),
			.S(gen[1272]),
			.SE(gen[1273]),

			.SELF(gen[1212]),
			.cell_state(gen[1212])
		); 

/******************* CELL 1213 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1213 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1152]),
			.N(gen[1153]),
			.NE(gen[1154]),

			.O(gen[1212]),
			.E(gen[1214]),

			.SO(gen[1272]),
			.S(gen[1273]),
			.SE(gen[1274]),

			.SELF(gen[1213]),
			.cell_state(gen[1213])
		); 

/******************* CELL 1214 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1214 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1153]),
			.N(gen[1154]),
			.NE(gen[1155]),

			.O(gen[1213]),
			.E(gen[1215]),

			.SO(gen[1273]),
			.S(gen[1274]),
			.SE(gen[1275]),

			.SELF(gen[1214]),
			.cell_state(gen[1214])
		); 

/******************* CELL 1215 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1215 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1154]),
			.N(gen[1155]),
			.NE(gen[1156]),

			.O(gen[1214]),
			.E(gen[1216]),

			.SO(gen[1274]),
			.S(gen[1275]),
			.SE(gen[1276]),

			.SELF(gen[1215]),
			.cell_state(gen[1215])
		); 

/******************* CELL 1216 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1216 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1155]),
			.N(gen[1156]),
			.NE(gen[1157]),

			.O(gen[1215]),
			.E(gen[1217]),

			.SO(gen[1275]),
			.S(gen[1276]),
			.SE(gen[1277]),

			.SELF(gen[1216]),
			.cell_state(gen[1216])
		); 

/******************* CELL 1217 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1217 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1156]),
			.N(gen[1157]),
			.NE(gen[1158]),

			.O(gen[1216]),
			.E(gen[1218]),

			.SO(gen[1276]),
			.S(gen[1277]),
			.SE(gen[1278]),

			.SELF(gen[1217]),
			.cell_state(gen[1217])
		); 

/******************* CELL 1218 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1218 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1157]),
			.N(gen[1158]),
			.NE(gen[1159]),

			.O(gen[1217]),
			.E(gen[1219]),

			.SO(gen[1277]),
			.S(gen[1278]),
			.SE(gen[1279]),

			.SELF(gen[1218]),
			.cell_state(gen[1218])
		); 

/******************* CELL 1219 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1219 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1158]),
			.N(gen[1159]),
			.NE(gen[1160]),

			.O(gen[1218]),
			.E(gen[1220]),

			.SO(gen[1278]),
			.S(gen[1279]),
			.SE(gen[1280]),

			.SELF(gen[1219]),
			.cell_state(gen[1219])
		); 

/******************* CELL 1220 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1220 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1159]),
			.N(gen[1160]),
			.NE(gen[1161]),

			.O(gen[1219]),
			.E(gen[1221]),

			.SO(gen[1279]),
			.S(gen[1280]),
			.SE(gen[1281]),

			.SELF(gen[1220]),
			.cell_state(gen[1220])
		); 

/******************* CELL 1221 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1221 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1160]),
			.N(gen[1161]),
			.NE(gen[1162]),

			.O(gen[1220]),
			.E(gen[1222]),

			.SO(gen[1280]),
			.S(gen[1281]),
			.SE(gen[1282]),

			.SELF(gen[1221]),
			.cell_state(gen[1221])
		); 

/******************* CELL 1222 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1222 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1161]),
			.N(gen[1162]),
			.NE(gen[1163]),

			.O(gen[1221]),
			.E(gen[1223]),

			.SO(gen[1281]),
			.S(gen[1282]),
			.SE(gen[1283]),

			.SELF(gen[1222]),
			.cell_state(gen[1222])
		); 

/******************* CELL 1223 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1223 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1162]),
			.N(gen[1163]),
			.NE(gen[1164]),

			.O(gen[1222]),
			.E(gen[1224]),

			.SO(gen[1282]),
			.S(gen[1283]),
			.SE(gen[1284]),

			.SELF(gen[1223]),
			.cell_state(gen[1223])
		); 

/******************* CELL 1224 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1224 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1163]),
			.N(gen[1164]),
			.NE(gen[1165]),

			.O(gen[1223]),
			.E(gen[1225]),

			.SO(gen[1283]),
			.S(gen[1284]),
			.SE(gen[1285]),

			.SELF(gen[1224]),
			.cell_state(gen[1224])
		); 

/******************* CELL 1225 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1225 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1164]),
			.N(gen[1165]),
			.NE(gen[1166]),

			.O(gen[1224]),
			.E(gen[1226]),

			.SO(gen[1284]),
			.S(gen[1285]),
			.SE(gen[1286]),

			.SELF(gen[1225]),
			.cell_state(gen[1225])
		); 

/******************* CELL 1226 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1226 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1165]),
			.N(gen[1166]),
			.NE(gen[1167]),

			.O(gen[1225]),
			.E(gen[1227]),

			.SO(gen[1285]),
			.S(gen[1286]),
			.SE(gen[1287]),

			.SELF(gen[1226]),
			.cell_state(gen[1226])
		); 

/******************* CELL 1227 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1227 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1166]),
			.N(gen[1167]),
			.NE(gen[1168]),

			.O(gen[1226]),
			.E(gen[1228]),

			.SO(gen[1286]),
			.S(gen[1287]),
			.SE(gen[1288]),

			.SELF(gen[1227]),
			.cell_state(gen[1227])
		); 

/******************* CELL 1228 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1228 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1167]),
			.N(gen[1168]),
			.NE(gen[1169]),

			.O(gen[1227]),
			.E(gen[1229]),

			.SO(gen[1287]),
			.S(gen[1288]),
			.SE(gen[1289]),

			.SELF(gen[1228]),
			.cell_state(gen[1228])
		); 

/******************* CELL 1229 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1229 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1168]),
			.N(gen[1169]),
			.NE(gen[1170]),

			.O(gen[1228]),
			.E(gen[1230]),

			.SO(gen[1288]),
			.S(gen[1289]),
			.SE(gen[1290]),

			.SELF(gen[1229]),
			.cell_state(gen[1229])
		); 

/******************* CELL 1230 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1230 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1169]),
			.N(gen[1170]),
			.NE(gen[1171]),

			.O(gen[1229]),
			.E(gen[1231]),

			.SO(gen[1289]),
			.S(gen[1290]),
			.SE(gen[1291]),

			.SELF(gen[1230]),
			.cell_state(gen[1230])
		); 

/******************* CELL 1231 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1231 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1170]),
			.N(gen[1171]),
			.NE(gen[1172]),

			.O(gen[1230]),
			.E(gen[1232]),

			.SO(gen[1290]),
			.S(gen[1291]),
			.SE(gen[1292]),

			.SELF(gen[1231]),
			.cell_state(gen[1231])
		); 

/******************* CELL 1232 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1232 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1171]),
			.N(gen[1172]),
			.NE(gen[1173]),

			.O(gen[1231]),
			.E(gen[1233]),

			.SO(gen[1291]),
			.S(gen[1292]),
			.SE(gen[1293]),

			.SELF(gen[1232]),
			.cell_state(gen[1232])
		); 

/******************* CELL 1233 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1233 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1172]),
			.N(gen[1173]),
			.NE(gen[1174]),

			.O(gen[1232]),
			.E(gen[1234]),

			.SO(gen[1292]),
			.S(gen[1293]),
			.SE(gen[1294]),

			.SELF(gen[1233]),
			.cell_state(gen[1233])
		); 

/******************* CELL 1234 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1234 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1173]),
			.N(gen[1174]),
			.NE(gen[1175]),

			.O(gen[1233]),
			.E(gen[1235]),

			.SO(gen[1293]),
			.S(gen[1294]),
			.SE(gen[1295]),

			.SELF(gen[1234]),
			.cell_state(gen[1234])
		); 

/******************* CELL 1235 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1235 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1174]),
			.N(gen[1175]),
			.NE(gen[1176]),

			.O(gen[1234]),
			.E(gen[1236]),

			.SO(gen[1294]),
			.S(gen[1295]),
			.SE(gen[1296]),

			.SELF(gen[1235]),
			.cell_state(gen[1235])
		); 

/******************* CELL 1236 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1236 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1175]),
			.N(gen[1176]),
			.NE(gen[1177]),

			.O(gen[1235]),
			.E(gen[1237]),

			.SO(gen[1295]),
			.S(gen[1296]),
			.SE(gen[1297]),

			.SELF(gen[1236]),
			.cell_state(gen[1236])
		); 

/******************* CELL 1237 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1237 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1176]),
			.N(gen[1177]),
			.NE(gen[1178]),

			.O(gen[1236]),
			.E(gen[1238]),

			.SO(gen[1296]),
			.S(gen[1297]),
			.SE(gen[1298]),

			.SELF(gen[1237]),
			.cell_state(gen[1237])
		); 

/******************* CELL 1238 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1238 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1177]),
			.N(gen[1178]),
			.NE(gen[1179]),

			.O(gen[1237]),
			.E(gen[1239]),

			.SO(gen[1297]),
			.S(gen[1298]),
			.SE(gen[1299]),

			.SELF(gen[1238]),
			.cell_state(gen[1238])
		); 

/******************* CELL 1239 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1239 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1178]),
			.N(gen[1179]),
			.NE(gen[1180]),

			.O(gen[1238]),
			.E(gen[1240]),

			.SO(gen[1298]),
			.S(gen[1299]),
			.SE(gen[1300]),

			.SELF(gen[1239]),
			.cell_state(gen[1239])
		); 

/******************* CELL 1240 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1240 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1179]),
			.N(gen[1180]),
			.NE(gen[1181]),

			.O(gen[1239]),
			.E(gen[1241]),

			.SO(gen[1299]),
			.S(gen[1300]),
			.SE(gen[1301]),

			.SELF(gen[1240]),
			.cell_state(gen[1240])
		); 

/******************* CELL 1241 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1241 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1180]),
			.N(gen[1181]),
			.NE(gen[1182]),

			.O(gen[1240]),
			.E(gen[1242]),

			.SO(gen[1300]),
			.S(gen[1301]),
			.SE(gen[1302]),

			.SELF(gen[1241]),
			.cell_state(gen[1241])
		); 

/******************* CELL 1242 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1242 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1181]),
			.N(gen[1182]),
			.NE(gen[1183]),

			.O(gen[1241]),
			.E(gen[1243]),

			.SO(gen[1301]),
			.S(gen[1302]),
			.SE(gen[1303]),

			.SELF(gen[1242]),
			.cell_state(gen[1242])
		); 

/******************* CELL 1243 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1243 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1182]),
			.N(gen[1183]),
			.NE(gen[1184]),

			.O(gen[1242]),
			.E(gen[1244]),

			.SO(gen[1302]),
			.S(gen[1303]),
			.SE(gen[1304]),

			.SELF(gen[1243]),
			.cell_state(gen[1243])
		); 

/******************* CELL 1244 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1244 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1183]),
			.N(gen[1184]),
			.NE(gen[1185]),

			.O(gen[1243]),
			.E(gen[1245]),

			.SO(gen[1303]),
			.S(gen[1304]),
			.SE(gen[1305]),

			.SELF(gen[1244]),
			.cell_state(gen[1244])
		); 

/******************* CELL 1245 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1245 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1184]),
			.N(gen[1185]),
			.NE(gen[1186]),

			.O(gen[1244]),
			.E(gen[1246]),

			.SO(gen[1304]),
			.S(gen[1305]),
			.SE(gen[1306]),

			.SELF(gen[1245]),
			.cell_state(gen[1245])
		); 

/******************* CELL 1246 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1246 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1185]),
			.N(gen[1186]),
			.NE(gen[1187]),

			.O(gen[1245]),
			.E(gen[1247]),

			.SO(gen[1305]),
			.S(gen[1306]),
			.SE(gen[1307]),

			.SELF(gen[1246]),
			.cell_state(gen[1246])
		); 

/******************* CELL 1247 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1247 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1186]),
			.N(gen[1187]),
			.NE(gen[1188]),

			.O(gen[1246]),
			.E(gen[1248]),

			.SO(gen[1306]),
			.S(gen[1307]),
			.SE(gen[1308]),

			.SELF(gen[1247]),
			.cell_state(gen[1247])
		); 

/******************* CELL 1248 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1248 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1187]),
			.N(gen[1188]),
			.NE(gen[1189]),

			.O(gen[1247]),
			.E(gen[1249]),

			.SO(gen[1307]),
			.S(gen[1308]),
			.SE(gen[1309]),

			.SELF(gen[1248]),
			.cell_state(gen[1248])
		); 

/******************* CELL 1249 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1249 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1188]),
			.N(gen[1189]),
			.NE(gen[1190]),

			.O(gen[1248]),
			.E(gen[1250]),

			.SO(gen[1308]),
			.S(gen[1309]),
			.SE(gen[1310]),

			.SELF(gen[1249]),
			.cell_state(gen[1249])
		); 

/******************* CELL 1250 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1250 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1189]),
			.N(gen[1190]),
			.NE(gen[1191]),

			.O(gen[1249]),
			.E(gen[1251]),

			.SO(gen[1309]),
			.S(gen[1310]),
			.SE(gen[1311]),

			.SELF(gen[1250]),
			.cell_state(gen[1250])
		); 

/******************* CELL 1251 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1251 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1190]),
			.N(gen[1191]),
			.NE(gen[1192]),

			.O(gen[1250]),
			.E(gen[1252]),

			.SO(gen[1310]),
			.S(gen[1311]),
			.SE(gen[1312]),

			.SELF(gen[1251]),
			.cell_state(gen[1251])
		); 

/******************* CELL 1252 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1252 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1191]),
			.N(gen[1192]),
			.NE(gen[1193]),

			.O(gen[1251]),
			.E(gen[1253]),

			.SO(gen[1311]),
			.S(gen[1312]),
			.SE(gen[1313]),

			.SELF(gen[1252]),
			.cell_state(gen[1252])
		); 

/******************* CELL 1253 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1253 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1192]),
			.N(gen[1193]),
			.NE(gen[1194]),

			.O(gen[1252]),
			.E(gen[1254]),

			.SO(gen[1312]),
			.S(gen[1313]),
			.SE(gen[1314]),

			.SELF(gen[1253]),
			.cell_state(gen[1253])
		); 

/******************* CELL 1254 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1254 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1193]),
			.N(gen[1194]),
			.NE(gen[1195]),

			.O(gen[1253]),
			.E(gen[1255]),

			.SO(gen[1313]),
			.S(gen[1314]),
			.SE(gen[1315]),

			.SELF(gen[1254]),
			.cell_state(gen[1254])
		); 

/******************* CELL 1255 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1255 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1194]),
			.N(gen[1195]),
			.NE(gen[1196]),

			.O(gen[1254]),
			.E(gen[1256]),

			.SO(gen[1314]),
			.S(gen[1315]),
			.SE(gen[1316]),

			.SELF(gen[1255]),
			.cell_state(gen[1255])
		); 

/******************* CELL 1256 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1256 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1195]),
			.N(gen[1196]),
			.NE(gen[1197]),

			.O(gen[1255]),
			.E(gen[1257]),

			.SO(gen[1315]),
			.S(gen[1316]),
			.SE(gen[1317]),

			.SELF(gen[1256]),
			.cell_state(gen[1256])
		); 

/******************* CELL 1257 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1257 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1196]),
			.N(gen[1197]),
			.NE(gen[1198]),

			.O(gen[1256]),
			.E(gen[1258]),

			.SO(gen[1316]),
			.S(gen[1317]),
			.SE(gen[1318]),

			.SELF(gen[1257]),
			.cell_state(gen[1257])
		); 

/******************* CELL 1258 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1258 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1197]),
			.N(gen[1198]),
			.NE(gen[1199]),

			.O(gen[1257]),
			.E(gen[1259]),

			.SO(gen[1317]),
			.S(gen[1318]),
			.SE(gen[1319]),

			.SELF(gen[1258]),
			.cell_state(gen[1258])
		); 

/******************* CELL 1259 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1259 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1198]),
			.N(gen[1199]),
			.NE(gen[1198]),

			.O(gen[1258]),
			.E(gen[1258]),

			.SO(gen[1318]),
			.S(gen[1319]),
			.SE(gen[1318]),

			.SELF(gen[1259]),
			.cell_state(gen[1259])
		); 

/******************* CELL 1260 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1260 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1201]),
			.N(gen[1200]),
			.NE(gen[1201]),

			.O(gen[1261]),
			.E(gen[1261]),

			.SO(gen[1321]),
			.S(gen[1320]),
			.SE(gen[1321]),

			.SELF(gen[1260]),
			.cell_state(gen[1260])
		); 

/******************* CELL 1261 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1261 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1200]),
			.N(gen[1201]),
			.NE(gen[1202]),

			.O(gen[1260]),
			.E(gen[1262]),

			.SO(gen[1320]),
			.S(gen[1321]),
			.SE(gen[1322]),

			.SELF(gen[1261]),
			.cell_state(gen[1261])
		); 

/******************* CELL 1262 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1262 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1201]),
			.N(gen[1202]),
			.NE(gen[1203]),

			.O(gen[1261]),
			.E(gen[1263]),

			.SO(gen[1321]),
			.S(gen[1322]),
			.SE(gen[1323]),

			.SELF(gen[1262]),
			.cell_state(gen[1262])
		); 

/******************* CELL 1263 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1263 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1202]),
			.N(gen[1203]),
			.NE(gen[1204]),

			.O(gen[1262]),
			.E(gen[1264]),

			.SO(gen[1322]),
			.S(gen[1323]),
			.SE(gen[1324]),

			.SELF(gen[1263]),
			.cell_state(gen[1263])
		); 

/******************* CELL 1264 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1264 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1203]),
			.N(gen[1204]),
			.NE(gen[1205]),

			.O(gen[1263]),
			.E(gen[1265]),

			.SO(gen[1323]),
			.S(gen[1324]),
			.SE(gen[1325]),

			.SELF(gen[1264]),
			.cell_state(gen[1264])
		); 

/******************* CELL 1265 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1265 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1204]),
			.N(gen[1205]),
			.NE(gen[1206]),

			.O(gen[1264]),
			.E(gen[1266]),

			.SO(gen[1324]),
			.S(gen[1325]),
			.SE(gen[1326]),

			.SELF(gen[1265]),
			.cell_state(gen[1265])
		); 

/******************* CELL 1266 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1266 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1205]),
			.N(gen[1206]),
			.NE(gen[1207]),

			.O(gen[1265]),
			.E(gen[1267]),

			.SO(gen[1325]),
			.S(gen[1326]),
			.SE(gen[1327]),

			.SELF(gen[1266]),
			.cell_state(gen[1266])
		); 

/******************* CELL 1267 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1267 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1206]),
			.N(gen[1207]),
			.NE(gen[1208]),

			.O(gen[1266]),
			.E(gen[1268]),

			.SO(gen[1326]),
			.S(gen[1327]),
			.SE(gen[1328]),

			.SELF(gen[1267]),
			.cell_state(gen[1267])
		); 

/******************* CELL 1268 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1268 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1207]),
			.N(gen[1208]),
			.NE(gen[1209]),

			.O(gen[1267]),
			.E(gen[1269]),

			.SO(gen[1327]),
			.S(gen[1328]),
			.SE(gen[1329]),

			.SELF(gen[1268]),
			.cell_state(gen[1268])
		); 

/******************* CELL 1269 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1269 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1208]),
			.N(gen[1209]),
			.NE(gen[1210]),

			.O(gen[1268]),
			.E(gen[1270]),

			.SO(gen[1328]),
			.S(gen[1329]),
			.SE(gen[1330]),

			.SELF(gen[1269]),
			.cell_state(gen[1269])
		); 

/******************* CELL 1270 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1270 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1209]),
			.N(gen[1210]),
			.NE(gen[1211]),

			.O(gen[1269]),
			.E(gen[1271]),

			.SO(gen[1329]),
			.S(gen[1330]),
			.SE(gen[1331]),

			.SELF(gen[1270]),
			.cell_state(gen[1270])
		); 

/******************* CELL 1271 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1271 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1210]),
			.N(gen[1211]),
			.NE(gen[1212]),

			.O(gen[1270]),
			.E(gen[1272]),

			.SO(gen[1330]),
			.S(gen[1331]),
			.SE(gen[1332]),

			.SELF(gen[1271]),
			.cell_state(gen[1271])
		); 

/******************* CELL 1272 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1272 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1211]),
			.N(gen[1212]),
			.NE(gen[1213]),

			.O(gen[1271]),
			.E(gen[1273]),

			.SO(gen[1331]),
			.S(gen[1332]),
			.SE(gen[1333]),

			.SELF(gen[1272]),
			.cell_state(gen[1272])
		); 

/******************* CELL 1273 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1273 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1212]),
			.N(gen[1213]),
			.NE(gen[1214]),

			.O(gen[1272]),
			.E(gen[1274]),

			.SO(gen[1332]),
			.S(gen[1333]),
			.SE(gen[1334]),

			.SELF(gen[1273]),
			.cell_state(gen[1273])
		); 

/******************* CELL 1274 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1274 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1213]),
			.N(gen[1214]),
			.NE(gen[1215]),

			.O(gen[1273]),
			.E(gen[1275]),

			.SO(gen[1333]),
			.S(gen[1334]),
			.SE(gen[1335]),

			.SELF(gen[1274]),
			.cell_state(gen[1274])
		); 

/******************* CELL 1275 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1275 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1214]),
			.N(gen[1215]),
			.NE(gen[1216]),

			.O(gen[1274]),
			.E(gen[1276]),

			.SO(gen[1334]),
			.S(gen[1335]),
			.SE(gen[1336]),

			.SELF(gen[1275]),
			.cell_state(gen[1275])
		); 

/******************* CELL 1276 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1276 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1215]),
			.N(gen[1216]),
			.NE(gen[1217]),

			.O(gen[1275]),
			.E(gen[1277]),

			.SO(gen[1335]),
			.S(gen[1336]),
			.SE(gen[1337]),

			.SELF(gen[1276]),
			.cell_state(gen[1276])
		); 

/******************* CELL 1277 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1277 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1216]),
			.N(gen[1217]),
			.NE(gen[1218]),

			.O(gen[1276]),
			.E(gen[1278]),

			.SO(gen[1336]),
			.S(gen[1337]),
			.SE(gen[1338]),

			.SELF(gen[1277]),
			.cell_state(gen[1277])
		); 

/******************* CELL 1278 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1278 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1217]),
			.N(gen[1218]),
			.NE(gen[1219]),

			.O(gen[1277]),
			.E(gen[1279]),

			.SO(gen[1337]),
			.S(gen[1338]),
			.SE(gen[1339]),

			.SELF(gen[1278]),
			.cell_state(gen[1278])
		); 

/******************* CELL 1279 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1279 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1218]),
			.N(gen[1219]),
			.NE(gen[1220]),

			.O(gen[1278]),
			.E(gen[1280]),

			.SO(gen[1338]),
			.S(gen[1339]),
			.SE(gen[1340]),

			.SELF(gen[1279]),
			.cell_state(gen[1279])
		); 

/******************* CELL 1280 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1280 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1219]),
			.N(gen[1220]),
			.NE(gen[1221]),

			.O(gen[1279]),
			.E(gen[1281]),

			.SO(gen[1339]),
			.S(gen[1340]),
			.SE(gen[1341]),

			.SELF(gen[1280]),
			.cell_state(gen[1280])
		); 

/******************* CELL 1281 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1281 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1220]),
			.N(gen[1221]),
			.NE(gen[1222]),

			.O(gen[1280]),
			.E(gen[1282]),

			.SO(gen[1340]),
			.S(gen[1341]),
			.SE(gen[1342]),

			.SELF(gen[1281]),
			.cell_state(gen[1281])
		); 

/******************* CELL 1282 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1282 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1221]),
			.N(gen[1222]),
			.NE(gen[1223]),

			.O(gen[1281]),
			.E(gen[1283]),

			.SO(gen[1341]),
			.S(gen[1342]),
			.SE(gen[1343]),

			.SELF(gen[1282]),
			.cell_state(gen[1282])
		); 

/******************* CELL 1283 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1283 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1222]),
			.N(gen[1223]),
			.NE(gen[1224]),

			.O(gen[1282]),
			.E(gen[1284]),

			.SO(gen[1342]),
			.S(gen[1343]),
			.SE(gen[1344]),

			.SELF(gen[1283]),
			.cell_state(gen[1283])
		); 

/******************* CELL 1284 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1284 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1223]),
			.N(gen[1224]),
			.NE(gen[1225]),

			.O(gen[1283]),
			.E(gen[1285]),

			.SO(gen[1343]),
			.S(gen[1344]),
			.SE(gen[1345]),

			.SELF(gen[1284]),
			.cell_state(gen[1284])
		); 

/******************* CELL 1285 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1285 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1224]),
			.N(gen[1225]),
			.NE(gen[1226]),

			.O(gen[1284]),
			.E(gen[1286]),

			.SO(gen[1344]),
			.S(gen[1345]),
			.SE(gen[1346]),

			.SELF(gen[1285]),
			.cell_state(gen[1285])
		); 

/******************* CELL 1286 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1286 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1225]),
			.N(gen[1226]),
			.NE(gen[1227]),

			.O(gen[1285]),
			.E(gen[1287]),

			.SO(gen[1345]),
			.S(gen[1346]),
			.SE(gen[1347]),

			.SELF(gen[1286]),
			.cell_state(gen[1286])
		); 

/******************* CELL 1287 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1287 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1226]),
			.N(gen[1227]),
			.NE(gen[1228]),

			.O(gen[1286]),
			.E(gen[1288]),

			.SO(gen[1346]),
			.S(gen[1347]),
			.SE(gen[1348]),

			.SELF(gen[1287]),
			.cell_state(gen[1287])
		); 

/******************* CELL 1288 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1288 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1227]),
			.N(gen[1228]),
			.NE(gen[1229]),

			.O(gen[1287]),
			.E(gen[1289]),

			.SO(gen[1347]),
			.S(gen[1348]),
			.SE(gen[1349]),

			.SELF(gen[1288]),
			.cell_state(gen[1288])
		); 

/******************* CELL 1289 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1289 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1228]),
			.N(gen[1229]),
			.NE(gen[1230]),

			.O(gen[1288]),
			.E(gen[1290]),

			.SO(gen[1348]),
			.S(gen[1349]),
			.SE(gen[1350]),

			.SELF(gen[1289]),
			.cell_state(gen[1289])
		); 

/******************* CELL 1290 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1290 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1229]),
			.N(gen[1230]),
			.NE(gen[1231]),

			.O(gen[1289]),
			.E(gen[1291]),

			.SO(gen[1349]),
			.S(gen[1350]),
			.SE(gen[1351]),

			.SELF(gen[1290]),
			.cell_state(gen[1290])
		); 

/******************* CELL 1291 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1291 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1230]),
			.N(gen[1231]),
			.NE(gen[1232]),

			.O(gen[1290]),
			.E(gen[1292]),

			.SO(gen[1350]),
			.S(gen[1351]),
			.SE(gen[1352]),

			.SELF(gen[1291]),
			.cell_state(gen[1291])
		); 

/******************* CELL 1292 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1292 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1231]),
			.N(gen[1232]),
			.NE(gen[1233]),

			.O(gen[1291]),
			.E(gen[1293]),

			.SO(gen[1351]),
			.S(gen[1352]),
			.SE(gen[1353]),

			.SELF(gen[1292]),
			.cell_state(gen[1292])
		); 

/******************* CELL 1293 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1293 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1232]),
			.N(gen[1233]),
			.NE(gen[1234]),

			.O(gen[1292]),
			.E(gen[1294]),

			.SO(gen[1352]),
			.S(gen[1353]),
			.SE(gen[1354]),

			.SELF(gen[1293]),
			.cell_state(gen[1293])
		); 

/******************* CELL 1294 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1294 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1233]),
			.N(gen[1234]),
			.NE(gen[1235]),

			.O(gen[1293]),
			.E(gen[1295]),

			.SO(gen[1353]),
			.S(gen[1354]),
			.SE(gen[1355]),

			.SELF(gen[1294]),
			.cell_state(gen[1294])
		); 

/******************* CELL 1295 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1295 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1234]),
			.N(gen[1235]),
			.NE(gen[1236]),

			.O(gen[1294]),
			.E(gen[1296]),

			.SO(gen[1354]),
			.S(gen[1355]),
			.SE(gen[1356]),

			.SELF(gen[1295]),
			.cell_state(gen[1295])
		); 

/******************* CELL 1296 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1296 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1235]),
			.N(gen[1236]),
			.NE(gen[1237]),

			.O(gen[1295]),
			.E(gen[1297]),

			.SO(gen[1355]),
			.S(gen[1356]),
			.SE(gen[1357]),

			.SELF(gen[1296]),
			.cell_state(gen[1296])
		); 

/******************* CELL 1297 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1297 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1236]),
			.N(gen[1237]),
			.NE(gen[1238]),

			.O(gen[1296]),
			.E(gen[1298]),

			.SO(gen[1356]),
			.S(gen[1357]),
			.SE(gen[1358]),

			.SELF(gen[1297]),
			.cell_state(gen[1297])
		); 

/******************* CELL 1298 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1298 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1237]),
			.N(gen[1238]),
			.NE(gen[1239]),

			.O(gen[1297]),
			.E(gen[1299]),

			.SO(gen[1357]),
			.S(gen[1358]),
			.SE(gen[1359]),

			.SELF(gen[1298]),
			.cell_state(gen[1298])
		); 

/******************* CELL 1299 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1299 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1238]),
			.N(gen[1239]),
			.NE(gen[1240]),

			.O(gen[1298]),
			.E(gen[1300]),

			.SO(gen[1358]),
			.S(gen[1359]),
			.SE(gen[1360]),

			.SELF(gen[1299]),
			.cell_state(gen[1299])
		); 

/******************* CELL 1300 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1300 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1239]),
			.N(gen[1240]),
			.NE(gen[1241]),

			.O(gen[1299]),
			.E(gen[1301]),

			.SO(gen[1359]),
			.S(gen[1360]),
			.SE(gen[1361]),

			.SELF(gen[1300]),
			.cell_state(gen[1300])
		); 

/******************* CELL 1301 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1301 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1240]),
			.N(gen[1241]),
			.NE(gen[1242]),

			.O(gen[1300]),
			.E(gen[1302]),

			.SO(gen[1360]),
			.S(gen[1361]),
			.SE(gen[1362]),

			.SELF(gen[1301]),
			.cell_state(gen[1301])
		); 

/******************* CELL 1302 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1302 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1241]),
			.N(gen[1242]),
			.NE(gen[1243]),

			.O(gen[1301]),
			.E(gen[1303]),

			.SO(gen[1361]),
			.S(gen[1362]),
			.SE(gen[1363]),

			.SELF(gen[1302]),
			.cell_state(gen[1302])
		); 

/******************* CELL 1303 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1303 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1242]),
			.N(gen[1243]),
			.NE(gen[1244]),

			.O(gen[1302]),
			.E(gen[1304]),

			.SO(gen[1362]),
			.S(gen[1363]),
			.SE(gen[1364]),

			.SELF(gen[1303]),
			.cell_state(gen[1303])
		); 

/******************* CELL 1304 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1304 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1243]),
			.N(gen[1244]),
			.NE(gen[1245]),

			.O(gen[1303]),
			.E(gen[1305]),

			.SO(gen[1363]),
			.S(gen[1364]),
			.SE(gen[1365]),

			.SELF(gen[1304]),
			.cell_state(gen[1304])
		); 

/******************* CELL 1305 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1305 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1244]),
			.N(gen[1245]),
			.NE(gen[1246]),

			.O(gen[1304]),
			.E(gen[1306]),

			.SO(gen[1364]),
			.S(gen[1365]),
			.SE(gen[1366]),

			.SELF(gen[1305]),
			.cell_state(gen[1305])
		); 

/******************* CELL 1306 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1306 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1245]),
			.N(gen[1246]),
			.NE(gen[1247]),

			.O(gen[1305]),
			.E(gen[1307]),

			.SO(gen[1365]),
			.S(gen[1366]),
			.SE(gen[1367]),

			.SELF(gen[1306]),
			.cell_state(gen[1306])
		); 

/******************* CELL 1307 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1307 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1246]),
			.N(gen[1247]),
			.NE(gen[1248]),

			.O(gen[1306]),
			.E(gen[1308]),

			.SO(gen[1366]),
			.S(gen[1367]),
			.SE(gen[1368]),

			.SELF(gen[1307]),
			.cell_state(gen[1307])
		); 

/******************* CELL 1308 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1308 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1247]),
			.N(gen[1248]),
			.NE(gen[1249]),

			.O(gen[1307]),
			.E(gen[1309]),

			.SO(gen[1367]),
			.S(gen[1368]),
			.SE(gen[1369]),

			.SELF(gen[1308]),
			.cell_state(gen[1308])
		); 

/******************* CELL 1309 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1309 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1248]),
			.N(gen[1249]),
			.NE(gen[1250]),

			.O(gen[1308]),
			.E(gen[1310]),

			.SO(gen[1368]),
			.S(gen[1369]),
			.SE(gen[1370]),

			.SELF(gen[1309]),
			.cell_state(gen[1309])
		); 

/******************* CELL 1310 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1310 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1249]),
			.N(gen[1250]),
			.NE(gen[1251]),

			.O(gen[1309]),
			.E(gen[1311]),

			.SO(gen[1369]),
			.S(gen[1370]),
			.SE(gen[1371]),

			.SELF(gen[1310]),
			.cell_state(gen[1310])
		); 

/******************* CELL 1311 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1311 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1250]),
			.N(gen[1251]),
			.NE(gen[1252]),

			.O(gen[1310]),
			.E(gen[1312]),

			.SO(gen[1370]),
			.S(gen[1371]),
			.SE(gen[1372]),

			.SELF(gen[1311]),
			.cell_state(gen[1311])
		); 

/******************* CELL 1312 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1312 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1251]),
			.N(gen[1252]),
			.NE(gen[1253]),

			.O(gen[1311]),
			.E(gen[1313]),

			.SO(gen[1371]),
			.S(gen[1372]),
			.SE(gen[1373]),

			.SELF(gen[1312]),
			.cell_state(gen[1312])
		); 

/******************* CELL 1313 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1313 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1252]),
			.N(gen[1253]),
			.NE(gen[1254]),

			.O(gen[1312]),
			.E(gen[1314]),

			.SO(gen[1372]),
			.S(gen[1373]),
			.SE(gen[1374]),

			.SELF(gen[1313]),
			.cell_state(gen[1313])
		); 

/******************* CELL 1314 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1314 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1253]),
			.N(gen[1254]),
			.NE(gen[1255]),

			.O(gen[1313]),
			.E(gen[1315]),

			.SO(gen[1373]),
			.S(gen[1374]),
			.SE(gen[1375]),

			.SELF(gen[1314]),
			.cell_state(gen[1314])
		); 

/******************* CELL 1315 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1315 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1254]),
			.N(gen[1255]),
			.NE(gen[1256]),

			.O(gen[1314]),
			.E(gen[1316]),

			.SO(gen[1374]),
			.S(gen[1375]),
			.SE(gen[1376]),

			.SELF(gen[1315]),
			.cell_state(gen[1315])
		); 

/******************* CELL 1316 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1316 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1255]),
			.N(gen[1256]),
			.NE(gen[1257]),

			.O(gen[1315]),
			.E(gen[1317]),

			.SO(gen[1375]),
			.S(gen[1376]),
			.SE(gen[1377]),

			.SELF(gen[1316]),
			.cell_state(gen[1316])
		); 

/******************* CELL 1317 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1317 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1256]),
			.N(gen[1257]),
			.NE(gen[1258]),

			.O(gen[1316]),
			.E(gen[1318]),

			.SO(gen[1376]),
			.S(gen[1377]),
			.SE(gen[1378]),

			.SELF(gen[1317]),
			.cell_state(gen[1317])
		); 

/******************* CELL 1318 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1318 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1257]),
			.N(gen[1258]),
			.NE(gen[1259]),

			.O(gen[1317]),
			.E(gen[1319]),

			.SO(gen[1377]),
			.S(gen[1378]),
			.SE(gen[1379]),

			.SELF(gen[1318]),
			.cell_state(gen[1318])
		); 

/******************* CELL 1319 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1319 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1258]),
			.N(gen[1259]),
			.NE(gen[1258]),

			.O(gen[1318]),
			.E(gen[1318]),

			.SO(gen[1378]),
			.S(gen[1379]),
			.SE(gen[1378]),

			.SELF(gen[1319]),
			.cell_state(gen[1319])
		); 

/******************* CELL 1320 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1320 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1261]),
			.N(gen[1260]),
			.NE(gen[1261]),

			.O(gen[1321]),
			.E(gen[1321]),

			.SO(gen[1381]),
			.S(gen[1380]),
			.SE(gen[1381]),

			.SELF(gen[1320]),
			.cell_state(gen[1320])
		); 

/******************* CELL 1321 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1321 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1260]),
			.N(gen[1261]),
			.NE(gen[1262]),

			.O(gen[1320]),
			.E(gen[1322]),

			.SO(gen[1380]),
			.S(gen[1381]),
			.SE(gen[1382]),

			.SELF(gen[1321]),
			.cell_state(gen[1321])
		); 

/******************* CELL 1322 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1322 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1261]),
			.N(gen[1262]),
			.NE(gen[1263]),

			.O(gen[1321]),
			.E(gen[1323]),

			.SO(gen[1381]),
			.S(gen[1382]),
			.SE(gen[1383]),

			.SELF(gen[1322]),
			.cell_state(gen[1322])
		); 

/******************* CELL 1323 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1323 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1262]),
			.N(gen[1263]),
			.NE(gen[1264]),

			.O(gen[1322]),
			.E(gen[1324]),

			.SO(gen[1382]),
			.S(gen[1383]),
			.SE(gen[1384]),

			.SELF(gen[1323]),
			.cell_state(gen[1323])
		); 

/******************* CELL 1324 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1324 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1263]),
			.N(gen[1264]),
			.NE(gen[1265]),

			.O(gen[1323]),
			.E(gen[1325]),

			.SO(gen[1383]),
			.S(gen[1384]),
			.SE(gen[1385]),

			.SELF(gen[1324]),
			.cell_state(gen[1324])
		); 

/******************* CELL 1325 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1325 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1264]),
			.N(gen[1265]),
			.NE(gen[1266]),

			.O(gen[1324]),
			.E(gen[1326]),

			.SO(gen[1384]),
			.S(gen[1385]),
			.SE(gen[1386]),

			.SELF(gen[1325]),
			.cell_state(gen[1325])
		); 

/******************* CELL 1326 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1326 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1265]),
			.N(gen[1266]),
			.NE(gen[1267]),

			.O(gen[1325]),
			.E(gen[1327]),

			.SO(gen[1385]),
			.S(gen[1386]),
			.SE(gen[1387]),

			.SELF(gen[1326]),
			.cell_state(gen[1326])
		); 

/******************* CELL 1327 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1327 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1266]),
			.N(gen[1267]),
			.NE(gen[1268]),

			.O(gen[1326]),
			.E(gen[1328]),

			.SO(gen[1386]),
			.S(gen[1387]),
			.SE(gen[1388]),

			.SELF(gen[1327]),
			.cell_state(gen[1327])
		); 

/******************* CELL 1328 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1328 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1267]),
			.N(gen[1268]),
			.NE(gen[1269]),

			.O(gen[1327]),
			.E(gen[1329]),

			.SO(gen[1387]),
			.S(gen[1388]),
			.SE(gen[1389]),

			.SELF(gen[1328]),
			.cell_state(gen[1328])
		); 

/******************* CELL 1329 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1329 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1268]),
			.N(gen[1269]),
			.NE(gen[1270]),

			.O(gen[1328]),
			.E(gen[1330]),

			.SO(gen[1388]),
			.S(gen[1389]),
			.SE(gen[1390]),

			.SELF(gen[1329]),
			.cell_state(gen[1329])
		); 

/******************* CELL 1330 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1330 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1269]),
			.N(gen[1270]),
			.NE(gen[1271]),

			.O(gen[1329]),
			.E(gen[1331]),

			.SO(gen[1389]),
			.S(gen[1390]),
			.SE(gen[1391]),

			.SELF(gen[1330]),
			.cell_state(gen[1330])
		); 

/******************* CELL 1331 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1331 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1270]),
			.N(gen[1271]),
			.NE(gen[1272]),

			.O(gen[1330]),
			.E(gen[1332]),

			.SO(gen[1390]),
			.S(gen[1391]),
			.SE(gen[1392]),

			.SELF(gen[1331]),
			.cell_state(gen[1331])
		); 

/******************* CELL 1332 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1332 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1271]),
			.N(gen[1272]),
			.NE(gen[1273]),

			.O(gen[1331]),
			.E(gen[1333]),

			.SO(gen[1391]),
			.S(gen[1392]),
			.SE(gen[1393]),

			.SELF(gen[1332]),
			.cell_state(gen[1332])
		); 

/******************* CELL 1333 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1333 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1272]),
			.N(gen[1273]),
			.NE(gen[1274]),

			.O(gen[1332]),
			.E(gen[1334]),

			.SO(gen[1392]),
			.S(gen[1393]),
			.SE(gen[1394]),

			.SELF(gen[1333]),
			.cell_state(gen[1333])
		); 

/******************* CELL 1334 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1334 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1273]),
			.N(gen[1274]),
			.NE(gen[1275]),

			.O(gen[1333]),
			.E(gen[1335]),

			.SO(gen[1393]),
			.S(gen[1394]),
			.SE(gen[1395]),

			.SELF(gen[1334]),
			.cell_state(gen[1334])
		); 

/******************* CELL 1335 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1335 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1274]),
			.N(gen[1275]),
			.NE(gen[1276]),

			.O(gen[1334]),
			.E(gen[1336]),

			.SO(gen[1394]),
			.S(gen[1395]),
			.SE(gen[1396]),

			.SELF(gen[1335]),
			.cell_state(gen[1335])
		); 

/******************* CELL 1336 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1336 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1275]),
			.N(gen[1276]),
			.NE(gen[1277]),

			.O(gen[1335]),
			.E(gen[1337]),

			.SO(gen[1395]),
			.S(gen[1396]),
			.SE(gen[1397]),

			.SELF(gen[1336]),
			.cell_state(gen[1336])
		); 

/******************* CELL 1337 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1337 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1276]),
			.N(gen[1277]),
			.NE(gen[1278]),

			.O(gen[1336]),
			.E(gen[1338]),

			.SO(gen[1396]),
			.S(gen[1397]),
			.SE(gen[1398]),

			.SELF(gen[1337]),
			.cell_state(gen[1337])
		); 

/******************* CELL 1338 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1338 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1277]),
			.N(gen[1278]),
			.NE(gen[1279]),

			.O(gen[1337]),
			.E(gen[1339]),

			.SO(gen[1397]),
			.S(gen[1398]),
			.SE(gen[1399]),

			.SELF(gen[1338]),
			.cell_state(gen[1338])
		); 

/******************* CELL 1339 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1339 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1278]),
			.N(gen[1279]),
			.NE(gen[1280]),

			.O(gen[1338]),
			.E(gen[1340]),

			.SO(gen[1398]),
			.S(gen[1399]),
			.SE(gen[1400]),

			.SELF(gen[1339]),
			.cell_state(gen[1339])
		); 

/******************* CELL 1340 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1340 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1279]),
			.N(gen[1280]),
			.NE(gen[1281]),

			.O(gen[1339]),
			.E(gen[1341]),

			.SO(gen[1399]),
			.S(gen[1400]),
			.SE(gen[1401]),

			.SELF(gen[1340]),
			.cell_state(gen[1340])
		); 

/******************* CELL 1341 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1341 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1280]),
			.N(gen[1281]),
			.NE(gen[1282]),

			.O(gen[1340]),
			.E(gen[1342]),

			.SO(gen[1400]),
			.S(gen[1401]),
			.SE(gen[1402]),

			.SELF(gen[1341]),
			.cell_state(gen[1341])
		); 

/******************* CELL 1342 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1342 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1281]),
			.N(gen[1282]),
			.NE(gen[1283]),

			.O(gen[1341]),
			.E(gen[1343]),

			.SO(gen[1401]),
			.S(gen[1402]),
			.SE(gen[1403]),

			.SELF(gen[1342]),
			.cell_state(gen[1342])
		); 

/******************* CELL 1343 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1343 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1282]),
			.N(gen[1283]),
			.NE(gen[1284]),

			.O(gen[1342]),
			.E(gen[1344]),

			.SO(gen[1402]),
			.S(gen[1403]),
			.SE(gen[1404]),

			.SELF(gen[1343]),
			.cell_state(gen[1343])
		); 

/******************* CELL 1344 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1344 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1283]),
			.N(gen[1284]),
			.NE(gen[1285]),

			.O(gen[1343]),
			.E(gen[1345]),

			.SO(gen[1403]),
			.S(gen[1404]),
			.SE(gen[1405]),

			.SELF(gen[1344]),
			.cell_state(gen[1344])
		); 

/******************* CELL 1345 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1345 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1284]),
			.N(gen[1285]),
			.NE(gen[1286]),

			.O(gen[1344]),
			.E(gen[1346]),

			.SO(gen[1404]),
			.S(gen[1405]),
			.SE(gen[1406]),

			.SELF(gen[1345]),
			.cell_state(gen[1345])
		); 

/******************* CELL 1346 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1346 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1285]),
			.N(gen[1286]),
			.NE(gen[1287]),

			.O(gen[1345]),
			.E(gen[1347]),

			.SO(gen[1405]),
			.S(gen[1406]),
			.SE(gen[1407]),

			.SELF(gen[1346]),
			.cell_state(gen[1346])
		); 

/******************* CELL 1347 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1347 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1286]),
			.N(gen[1287]),
			.NE(gen[1288]),

			.O(gen[1346]),
			.E(gen[1348]),

			.SO(gen[1406]),
			.S(gen[1407]),
			.SE(gen[1408]),

			.SELF(gen[1347]),
			.cell_state(gen[1347])
		); 

/******************* CELL 1348 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1348 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1287]),
			.N(gen[1288]),
			.NE(gen[1289]),

			.O(gen[1347]),
			.E(gen[1349]),

			.SO(gen[1407]),
			.S(gen[1408]),
			.SE(gen[1409]),

			.SELF(gen[1348]),
			.cell_state(gen[1348])
		); 

/******************* CELL 1349 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1349 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1288]),
			.N(gen[1289]),
			.NE(gen[1290]),

			.O(gen[1348]),
			.E(gen[1350]),

			.SO(gen[1408]),
			.S(gen[1409]),
			.SE(gen[1410]),

			.SELF(gen[1349]),
			.cell_state(gen[1349])
		); 

/******************* CELL 1350 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1350 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1289]),
			.N(gen[1290]),
			.NE(gen[1291]),

			.O(gen[1349]),
			.E(gen[1351]),

			.SO(gen[1409]),
			.S(gen[1410]),
			.SE(gen[1411]),

			.SELF(gen[1350]),
			.cell_state(gen[1350])
		); 

/******************* CELL 1351 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1351 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1290]),
			.N(gen[1291]),
			.NE(gen[1292]),

			.O(gen[1350]),
			.E(gen[1352]),

			.SO(gen[1410]),
			.S(gen[1411]),
			.SE(gen[1412]),

			.SELF(gen[1351]),
			.cell_state(gen[1351])
		); 

/******************* CELL 1352 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1352 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1291]),
			.N(gen[1292]),
			.NE(gen[1293]),

			.O(gen[1351]),
			.E(gen[1353]),

			.SO(gen[1411]),
			.S(gen[1412]),
			.SE(gen[1413]),

			.SELF(gen[1352]),
			.cell_state(gen[1352])
		); 

/******************* CELL 1353 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1353 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1292]),
			.N(gen[1293]),
			.NE(gen[1294]),

			.O(gen[1352]),
			.E(gen[1354]),

			.SO(gen[1412]),
			.S(gen[1413]),
			.SE(gen[1414]),

			.SELF(gen[1353]),
			.cell_state(gen[1353])
		); 

/******************* CELL 1354 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1354 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1293]),
			.N(gen[1294]),
			.NE(gen[1295]),

			.O(gen[1353]),
			.E(gen[1355]),

			.SO(gen[1413]),
			.S(gen[1414]),
			.SE(gen[1415]),

			.SELF(gen[1354]),
			.cell_state(gen[1354])
		); 

/******************* CELL 1355 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1355 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1294]),
			.N(gen[1295]),
			.NE(gen[1296]),

			.O(gen[1354]),
			.E(gen[1356]),

			.SO(gen[1414]),
			.S(gen[1415]),
			.SE(gen[1416]),

			.SELF(gen[1355]),
			.cell_state(gen[1355])
		); 

/******************* CELL 1356 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1356 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1295]),
			.N(gen[1296]),
			.NE(gen[1297]),

			.O(gen[1355]),
			.E(gen[1357]),

			.SO(gen[1415]),
			.S(gen[1416]),
			.SE(gen[1417]),

			.SELF(gen[1356]),
			.cell_state(gen[1356])
		); 

/******************* CELL 1357 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1357 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1296]),
			.N(gen[1297]),
			.NE(gen[1298]),

			.O(gen[1356]),
			.E(gen[1358]),

			.SO(gen[1416]),
			.S(gen[1417]),
			.SE(gen[1418]),

			.SELF(gen[1357]),
			.cell_state(gen[1357])
		); 

/******************* CELL 1358 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1358 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1297]),
			.N(gen[1298]),
			.NE(gen[1299]),

			.O(gen[1357]),
			.E(gen[1359]),

			.SO(gen[1417]),
			.S(gen[1418]),
			.SE(gen[1419]),

			.SELF(gen[1358]),
			.cell_state(gen[1358])
		); 

/******************* CELL 1359 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1359 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1298]),
			.N(gen[1299]),
			.NE(gen[1300]),

			.O(gen[1358]),
			.E(gen[1360]),

			.SO(gen[1418]),
			.S(gen[1419]),
			.SE(gen[1420]),

			.SELF(gen[1359]),
			.cell_state(gen[1359])
		); 

/******************* CELL 1360 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1360 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1299]),
			.N(gen[1300]),
			.NE(gen[1301]),

			.O(gen[1359]),
			.E(gen[1361]),

			.SO(gen[1419]),
			.S(gen[1420]),
			.SE(gen[1421]),

			.SELF(gen[1360]),
			.cell_state(gen[1360])
		); 

/******************* CELL 1361 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1361 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1300]),
			.N(gen[1301]),
			.NE(gen[1302]),

			.O(gen[1360]),
			.E(gen[1362]),

			.SO(gen[1420]),
			.S(gen[1421]),
			.SE(gen[1422]),

			.SELF(gen[1361]),
			.cell_state(gen[1361])
		); 

/******************* CELL 1362 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1362 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1301]),
			.N(gen[1302]),
			.NE(gen[1303]),

			.O(gen[1361]),
			.E(gen[1363]),

			.SO(gen[1421]),
			.S(gen[1422]),
			.SE(gen[1423]),

			.SELF(gen[1362]),
			.cell_state(gen[1362])
		); 

/******************* CELL 1363 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1363 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1302]),
			.N(gen[1303]),
			.NE(gen[1304]),

			.O(gen[1362]),
			.E(gen[1364]),

			.SO(gen[1422]),
			.S(gen[1423]),
			.SE(gen[1424]),

			.SELF(gen[1363]),
			.cell_state(gen[1363])
		); 

/******************* CELL 1364 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1364 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1303]),
			.N(gen[1304]),
			.NE(gen[1305]),

			.O(gen[1363]),
			.E(gen[1365]),

			.SO(gen[1423]),
			.S(gen[1424]),
			.SE(gen[1425]),

			.SELF(gen[1364]),
			.cell_state(gen[1364])
		); 

/******************* CELL 1365 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1365 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1304]),
			.N(gen[1305]),
			.NE(gen[1306]),

			.O(gen[1364]),
			.E(gen[1366]),

			.SO(gen[1424]),
			.S(gen[1425]),
			.SE(gen[1426]),

			.SELF(gen[1365]),
			.cell_state(gen[1365])
		); 

/******************* CELL 1366 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1366 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1305]),
			.N(gen[1306]),
			.NE(gen[1307]),

			.O(gen[1365]),
			.E(gen[1367]),

			.SO(gen[1425]),
			.S(gen[1426]),
			.SE(gen[1427]),

			.SELF(gen[1366]),
			.cell_state(gen[1366])
		); 

/******************* CELL 1367 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1367 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1306]),
			.N(gen[1307]),
			.NE(gen[1308]),

			.O(gen[1366]),
			.E(gen[1368]),

			.SO(gen[1426]),
			.S(gen[1427]),
			.SE(gen[1428]),

			.SELF(gen[1367]),
			.cell_state(gen[1367])
		); 

/******************* CELL 1368 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1368 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1307]),
			.N(gen[1308]),
			.NE(gen[1309]),

			.O(gen[1367]),
			.E(gen[1369]),

			.SO(gen[1427]),
			.S(gen[1428]),
			.SE(gen[1429]),

			.SELF(gen[1368]),
			.cell_state(gen[1368])
		); 

/******************* CELL 1369 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1369 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1308]),
			.N(gen[1309]),
			.NE(gen[1310]),

			.O(gen[1368]),
			.E(gen[1370]),

			.SO(gen[1428]),
			.S(gen[1429]),
			.SE(gen[1430]),

			.SELF(gen[1369]),
			.cell_state(gen[1369])
		); 

/******************* CELL 1370 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1370 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1309]),
			.N(gen[1310]),
			.NE(gen[1311]),

			.O(gen[1369]),
			.E(gen[1371]),

			.SO(gen[1429]),
			.S(gen[1430]),
			.SE(gen[1431]),

			.SELF(gen[1370]),
			.cell_state(gen[1370])
		); 

/******************* CELL 1371 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1371 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1310]),
			.N(gen[1311]),
			.NE(gen[1312]),

			.O(gen[1370]),
			.E(gen[1372]),

			.SO(gen[1430]),
			.S(gen[1431]),
			.SE(gen[1432]),

			.SELF(gen[1371]),
			.cell_state(gen[1371])
		); 

/******************* CELL 1372 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1372 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1311]),
			.N(gen[1312]),
			.NE(gen[1313]),

			.O(gen[1371]),
			.E(gen[1373]),

			.SO(gen[1431]),
			.S(gen[1432]),
			.SE(gen[1433]),

			.SELF(gen[1372]),
			.cell_state(gen[1372])
		); 

/******************* CELL 1373 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1373 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1312]),
			.N(gen[1313]),
			.NE(gen[1314]),

			.O(gen[1372]),
			.E(gen[1374]),

			.SO(gen[1432]),
			.S(gen[1433]),
			.SE(gen[1434]),

			.SELF(gen[1373]),
			.cell_state(gen[1373])
		); 

/******************* CELL 1374 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1374 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1313]),
			.N(gen[1314]),
			.NE(gen[1315]),

			.O(gen[1373]),
			.E(gen[1375]),

			.SO(gen[1433]),
			.S(gen[1434]),
			.SE(gen[1435]),

			.SELF(gen[1374]),
			.cell_state(gen[1374])
		); 

/******************* CELL 1375 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1375 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1314]),
			.N(gen[1315]),
			.NE(gen[1316]),

			.O(gen[1374]),
			.E(gen[1376]),

			.SO(gen[1434]),
			.S(gen[1435]),
			.SE(gen[1436]),

			.SELF(gen[1375]),
			.cell_state(gen[1375])
		); 

/******************* CELL 1376 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1376 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1315]),
			.N(gen[1316]),
			.NE(gen[1317]),

			.O(gen[1375]),
			.E(gen[1377]),

			.SO(gen[1435]),
			.S(gen[1436]),
			.SE(gen[1437]),

			.SELF(gen[1376]),
			.cell_state(gen[1376])
		); 

/******************* CELL 1377 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1377 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1316]),
			.N(gen[1317]),
			.NE(gen[1318]),

			.O(gen[1376]),
			.E(gen[1378]),

			.SO(gen[1436]),
			.S(gen[1437]),
			.SE(gen[1438]),

			.SELF(gen[1377]),
			.cell_state(gen[1377])
		); 

/******************* CELL 1378 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1378 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1317]),
			.N(gen[1318]),
			.NE(gen[1319]),

			.O(gen[1377]),
			.E(gen[1379]),

			.SO(gen[1437]),
			.S(gen[1438]),
			.SE(gen[1439]),

			.SELF(gen[1378]),
			.cell_state(gen[1378])
		); 

/******************* CELL 1379 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1379 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1318]),
			.N(gen[1319]),
			.NE(gen[1318]),

			.O(gen[1378]),
			.E(gen[1378]),

			.SO(gen[1438]),
			.S(gen[1439]),
			.SE(gen[1438]),

			.SELF(gen[1379]),
			.cell_state(gen[1379])
		); 

/******************* CELL 1380 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1380 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1321]),
			.N(gen[1320]),
			.NE(gen[1321]),

			.O(gen[1381]),
			.E(gen[1381]),

			.SO(gen[1441]),
			.S(gen[1440]),
			.SE(gen[1441]),

			.SELF(gen[1380]),
			.cell_state(gen[1380])
		); 

/******************* CELL 1381 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1381 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1320]),
			.N(gen[1321]),
			.NE(gen[1322]),

			.O(gen[1380]),
			.E(gen[1382]),

			.SO(gen[1440]),
			.S(gen[1441]),
			.SE(gen[1442]),

			.SELF(gen[1381]),
			.cell_state(gen[1381])
		); 

/******************* CELL 1382 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1382 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1321]),
			.N(gen[1322]),
			.NE(gen[1323]),

			.O(gen[1381]),
			.E(gen[1383]),

			.SO(gen[1441]),
			.S(gen[1442]),
			.SE(gen[1443]),

			.SELF(gen[1382]),
			.cell_state(gen[1382])
		); 

/******************* CELL 1383 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1383 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1322]),
			.N(gen[1323]),
			.NE(gen[1324]),

			.O(gen[1382]),
			.E(gen[1384]),

			.SO(gen[1442]),
			.S(gen[1443]),
			.SE(gen[1444]),

			.SELF(gen[1383]),
			.cell_state(gen[1383])
		); 

/******************* CELL 1384 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1384 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1323]),
			.N(gen[1324]),
			.NE(gen[1325]),

			.O(gen[1383]),
			.E(gen[1385]),

			.SO(gen[1443]),
			.S(gen[1444]),
			.SE(gen[1445]),

			.SELF(gen[1384]),
			.cell_state(gen[1384])
		); 

/******************* CELL 1385 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1385 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1324]),
			.N(gen[1325]),
			.NE(gen[1326]),

			.O(gen[1384]),
			.E(gen[1386]),

			.SO(gen[1444]),
			.S(gen[1445]),
			.SE(gen[1446]),

			.SELF(gen[1385]),
			.cell_state(gen[1385])
		); 

/******************* CELL 1386 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1386 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1325]),
			.N(gen[1326]),
			.NE(gen[1327]),

			.O(gen[1385]),
			.E(gen[1387]),

			.SO(gen[1445]),
			.S(gen[1446]),
			.SE(gen[1447]),

			.SELF(gen[1386]),
			.cell_state(gen[1386])
		); 

/******************* CELL 1387 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1387 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1326]),
			.N(gen[1327]),
			.NE(gen[1328]),

			.O(gen[1386]),
			.E(gen[1388]),

			.SO(gen[1446]),
			.S(gen[1447]),
			.SE(gen[1448]),

			.SELF(gen[1387]),
			.cell_state(gen[1387])
		); 

/******************* CELL 1388 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1388 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1327]),
			.N(gen[1328]),
			.NE(gen[1329]),

			.O(gen[1387]),
			.E(gen[1389]),

			.SO(gen[1447]),
			.S(gen[1448]),
			.SE(gen[1449]),

			.SELF(gen[1388]),
			.cell_state(gen[1388])
		); 

/******************* CELL 1389 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1389 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1328]),
			.N(gen[1329]),
			.NE(gen[1330]),

			.O(gen[1388]),
			.E(gen[1390]),

			.SO(gen[1448]),
			.S(gen[1449]),
			.SE(gen[1450]),

			.SELF(gen[1389]),
			.cell_state(gen[1389])
		); 

/******************* CELL 1390 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1390 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1329]),
			.N(gen[1330]),
			.NE(gen[1331]),

			.O(gen[1389]),
			.E(gen[1391]),

			.SO(gen[1449]),
			.S(gen[1450]),
			.SE(gen[1451]),

			.SELF(gen[1390]),
			.cell_state(gen[1390])
		); 

/******************* CELL 1391 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1391 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1330]),
			.N(gen[1331]),
			.NE(gen[1332]),

			.O(gen[1390]),
			.E(gen[1392]),

			.SO(gen[1450]),
			.S(gen[1451]),
			.SE(gen[1452]),

			.SELF(gen[1391]),
			.cell_state(gen[1391])
		); 

/******************* CELL 1392 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1392 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1331]),
			.N(gen[1332]),
			.NE(gen[1333]),

			.O(gen[1391]),
			.E(gen[1393]),

			.SO(gen[1451]),
			.S(gen[1452]),
			.SE(gen[1453]),

			.SELF(gen[1392]),
			.cell_state(gen[1392])
		); 

/******************* CELL 1393 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1393 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1332]),
			.N(gen[1333]),
			.NE(gen[1334]),

			.O(gen[1392]),
			.E(gen[1394]),

			.SO(gen[1452]),
			.S(gen[1453]),
			.SE(gen[1454]),

			.SELF(gen[1393]),
			.cell_state(gen[1393])
		); 

/******************* CELL 1394 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1394 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1333]),
			.N(gen[1334]),
			.NE(gen[1335]),

			.O(gen[1393]),
			.E(gen[1395]),

			.SO(gen[1453]),
			.S(gen[1454]),
			.SE(gen[1455]),

			.SELF(gen[1394]),
			.cell_state(gen[1394])
		); 

/******************* CELL 1395 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1395 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1334]),
			.N(gen[1335]),
			.NE(gen[1336]),

			.O(gen[1394]),
			.E(gen[1396]),

			.SO(gen[1454]),
			.S(gen[1455]),
			.SE(gen[1456]),

			.SELF(gen[1395]),
			.cell_state(gen[1395])
		); 

/******************* CELL 1396 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1396 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1335]),
			.N(gen[1336]),
			.NE(gen[1337]),

			.O(gen[1395]),
			.E(gen[1397]),

			.SO(gen[1455]),
			.S(gen[1456]),
			.SE(gen[1457]),

			.SELF(gen[1396]),
			.cell_state(gen[1396])
		); 

/******************* CELL 1397 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1397 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1336]),
			.N(gen[1337]),
			.NE(gen[1338]),

			.O(gen[1396]),
			.E(gen[1398]),

			.SO(gen[1456]),
			.S(gen[1457]),
			.SE(gen[1458]),

			.SELF(gen[1397]),
			.cell_state(gen[1397])
		); 

/******************* CELL 1398 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1398 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1337]),
			.N(gen[1338]),
			.NE(gen[1339]),

			.O(gen[1397]),
			.E(gen[1399]),

			.SO(gen[1457]),
			.S(gen[1458]),
			.SE(gen[1459]),

			.SELF(gen[1398]),
			.cell_state(gen[1398])
		); 

/******************* CELL 1399 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1399 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1338]),
			.N(gen[1339]),
			.NE(gen[1340]),

			.O(gen[1398]),
			.E(gen[1400]),

			.SO(gen[1458]),
			.S(gen[1459]),
			.SE(gen[1460]),

			.SELF(gen[1399]),
			.cell_state(gen[1399])
		); 

/******************* CELL 1400 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1400 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1339]),
			.N(gen[1340]),
			.NE(gen[1341]),

			.O(gen[1399]),
			.E(gen[1401]),

			.SO(gen[1459]),
			.S(gen[1460]),
			.SE(gen[1461]),

			.SELF(gen[1400]),
			.cell_state(gen[1400])
		); 

/******************* CELL 1401 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1401 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1340]),
			.N(gen[1341]),
			.NE(gen[1342]),

			.O(gen[1400]),
			.E(gen[1402]),

			.SO(gen[1460]),
			.S(gen[1461]),
			.SE(gen[1462]),

			.SELF(gen[1401]),
			.cell_state(gen[1401])
		); 

/******************* CELL 1402 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1402 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1341]),
			.N(gen[1342]),
			.NE(gen[1343]),

			.O(gen[1401]),
			.E(gen[1403]),

			.SO(gen[1461]),
			.S(gen[1462]),
			.SE(gen[1463]),

			.SELF(gen[1402]),
			.cell_state(gen[1402])
		); 

/******************* CELL 1403 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1403 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1342]),
			.N(gen[1343]),
			.NE(gen[1344]),

			.O(gen[1402]),
			.E(gen[1404]),

			.SO(gen[1462]),
			.S(gen[1463]),
			.SE(gen[1464]),

			.SELF(gen[1403]),
			.cell_state(gen[1403])
		); 

/******************* CELL 1404 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1404 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1343]),
			.N(gen[1344]),
			.NE(gen[1345]),

			.O(gen[1403]),
			.E(gen[1405]),

			.SO(gen[1463]),
			.S(gen[1464]),
			.SE(gen[1465]),

			.SELF(gen[1404]),
			.cell_state(gen[1404])
		); 

/******************* CELL 1405 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1405 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1344]),
			.N(gen[1345]),
			.NE(gen[1346]),

			.O(gen[1404]),
			.E(gen[1406]),

			.SO(gen[1464]),
			.S(gen[1465]),
			.SE(gen[1466]),

			.SELF(gen[1405]),
			.cell_state(gen[1405])
		); 

/******************* CELL 1406 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1406 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1345]),
			.N(gen[1346]),
			.NE(gen[1347]),

			.O(gen[1405]),
			.E(gen[1407]),

			.SO(gen[1465]),
			.S(gen[1466]),
			.SE(gen[1467]),

			.SELF(gen[1406]),
			.cell_state(gen[1406])
		); 

/******************* CELL 1407 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1407 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1346]),
			.N(gen[1347]),
			.NE(gen[1348]),

			.O(gen[1406]),
			.E(gen[1408]),

			.SO(gen[1466]),
			.S(gen[1467]),
			.SE(gen[1468]),

			.SELF(gen[1407]),
			.cell_state(gen[1407])
		); 

/******************* CELL 1408 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1408 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1347]),
			.N(gen[1348]),
			.NE(gen[1349]),

			.O(gen[1407]),
			.E(gen[1409]),

			.SO(gen[1467]),
			.S(gen[1468]),
			.SE(gen[1469]),

			.SELF(gen[1408]),
			.cell_state(gen[1408])
		); 

/******************* CELL 1409 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1409 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1348]),
			.N(gen[1349]),
			.NE(gen[1350]),

			.O(gen[1408]),
			.E(gen[1410]),

			.SO(gen[1468]),
			.S(gen[1469]),
			.SE(gen[1470]),

			.SELF(gen[1409]),
			.cell_state(gen[1409])
		); 

/******************* CELL 1410 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1410 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1349]),
			.N(gen[1350]),
			.NE(gen[1351]),

			.O(gen[1409]),
			.E(gen[1411]),

			.SO(gen[1469]),
			.S(gen[1470]),
			.SE(gen[1471]),

			.SELF(gen[1410]),
			.cell_state(gen[1410])
		); 

/******************* CELL 1411 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1411 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1350]),
			.N(gen[1351]),
			.NE(gen[1352]),

			.O(gen[1410]),
			.E(gen[1412]),

			.SO(gen[1470]),
			.S(gen[1471]),
			.SE(gen[1472]),

			.SELF(gen[1411]),
			.cell_state(gen[1411])
		); 

/******************* CELL 1412 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1412 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1351]),
			.N(gen[1352]),
			.NE(gen[1353]),

			.O(gen[1411]),
			.E(gen[1413]),

			.SO(gen[1471]),
			.S(gen[1472]),
			.SE(gen[1473]),

			.SELF(gen[1412]),
			.cell_state(gen[1412])
		); 

/******************* CELL 1413 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1413 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1352]),
			.N(gen[1353]),
			.NE(gen[1354]),

			.O(gen[1412]),
			.E(gen[1414]),

			.SO(gen[1472]),
			.S(gen[1473]),
			.SE(gen[1474]),

			.SELF(gen[1413]),
			.cell_state(gen[1413])
		); 

/******************* CELL 1414 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1414 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1353]),
			.N(gen[1354]),
			.NE(gen[1355]),

			.O(gen[1413]),
			.E(gen[1415]),

			.SO(gen[1473]),
			.S(gen[1474]),
			.SE(gen[1475]),

			.SELF(gen[1414]),
			.cell_state(gen[1414])
		); 

/******************* CELL 1415 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1415 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1354]),
			.N(gen[1355]),
			.NE(gen[1356]),

			.O(gen[1414]),
			.E(gen[1416]),

			.SO(gen[1474]),
			.S(gen[1475]),
			.SE(gen[1476]),

			.SELF(gen[1415]),
			.cell_state(gen[1415])
		); 

/******************* CELL 1416 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1416 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1355]),
			.N(gen[1356]),
			.NE(gen[1357]),

			.O(gen[1415]),
			.E(gen[1417]),

			.SO(gen[1475]),
			.S(gen[1476]),
			.SE(gen[1477]),

			.SELF(gen[1416]),
			.cell_state(gen[1416])
		); 

/******************* CELL 1417 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1417 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1356]),
			.N(gen[1357]),
			.NE(gen[1358]),

			.O(gen[1416]),
			.E(gen[1418]),

			.SO(gen[1476]),
			.S(gen[1477]),
			.SE(gen[1478]),

			.SELF(gen[1417]),
			.cell_state(gen[1417])
		); 

/******************* CELL 1418 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1418 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1357]),
			.N(gen[1358]),
			.NE(gen[1359]),

			.O(gen[1417]),
			.E(gen[1419]),

			.SO(gen[1477]),
			.S(gen[1478]),
			.SE(gen[1479]),

			.SELF(gen[1418]),
			.cell_state(gen[1418])
		); 

/******************* CELL 1419 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1419 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1358]),
			.N(gen[1359]),
			.NE(gen[1360]),

			.O(gen[1418]),
			.E(gen[1420]),

			.SO(gen[1478]),
			.S(gen[1479]),
			.SE(gen[1480]),

			.SELF(gen[1419]),
			.cell_state(gen[1419])
		); 

/******************* CELL 1420 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1420 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1359]),
			.N(gen[1360]),
			.NE(gen[1361]),

			.O(gen[1419]),
			.E(gen[1421]),

			.SO(gen[1479]),
			.S(gen[1480]),
			.SE(gen[1481]),

			.SELF(gen[1420]),
			.cell_state(gen[1420])
		); 

/******************* CELL 1421 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1421 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1360]),
			.N(gen[1361]),
			.NE(gen[1362]),

			.O(gen[1420]),
			.E(gen[1422]),

			.SO(gen[1480]),
			.S(gen[1481]),
			.SE(gen[1482]),

			.SELF(gen[1421]),
			.cell_state(gen[1421])
		); 

/******************* CELL 1422 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1422 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1361]),
			.N(gen[1362]),
			.NE(gen[1363]),

			.O(gen[1421]),
			.E(gen[1423]),

			.SO(gen[1481]),
			.S(gen[1482]),
			.SE(gen[1483]),

			.SELF(gen[1422]),
			.cell_state(gen[1422])
		); 

/******************* CELL 1423 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1423 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1362]),
			.N(gen[1363]),
			.NE(gen[1364]),

			.O(gen[1422]),
			.E(gen[1424]),

			.SO(gen[1482]),
			.S(gen[1483]),
			.SE(gen[1484]),

			.SELF(gen[1423]),
			.cell_state(gen[1423])
		); 

/******************* CELL 1424 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1424 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1363]),
			.N(gen[1364]),
			.NE(gen[1365]),

			.O(gen[1423]),
			.E(gen[1425]),

			.SO(gen[1483]),
			.S(gen[1484]),
			.SE(gen[1485]),

			.SELF(gen[1424]),
			.cell_state(gen[1424])
		); 

/******************* CELL 1425 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1425 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1364]),
			.N(gen[1365]),
			.NE(gen[1366]),

			.O(gen[1424]),
			.E(gen[1426]),

			.SO(gen[1484]),
			.S(gen[1485]),
			.SE(gen[1486]),

			.SELF(gen[1425]),
			.cell_state(gen[1425])
		); 

/******************* CELL 1426 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1426 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1365]),
			.N(gen[1366]),
			.NE(gen[1367]),

			.O(gen[1425]),
			.E(gen[1427]),

			.SO(gen[1485]),
			.S(gen[1486]),
			.SE(gen[1487]),

			.SELF(gen[1426]),
			.cell_state(gen[1426])
		); 

/******************* CELL 1427 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1427 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1366]),
			.N(gen[1367]),
			.NE(gen[1368]),

			.O(gen[1426]),
			.E(gen[1428]),

			.SO(gen[1486]),
			.S(gen[1487]),
			.SE(gen[1488]),

			.SELF(gen[1427]),
			.cell_state(gen[1427])
		); 

/******************* CELL 1428 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1428 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1367]),
			.N(gen[1368]),
			.NE(gen[1369]),

			.O(gen[1427]),
			.E(gen[1429]),

			.SO(gen[1487]),
			.S(gen[1488]),
			.SE(gen[1489]),

			.SELF(gen[1428]),
			.cell_state(gen[1428])
		); 

/******************* CELL 1429 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1429 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1368]),
			.N(gen[1369]),
			.NE(gen[1370]),

			.O(gen[1428]),
			.E(gen[1430]),

			.SO(gen[1488]),
			.S(gen[1489]),
			.SE(gen[1490]),

			.SELF(gen[1429]),
			.cell_state(gen[1429])
		); 

/******************* CELL 1430 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1430 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1369]),
			.N(gen[1370]),
			.NE(gen[1371]),

			.O(gen[1429]),
			.E(gen[1431]),

			.SO(gen[1489]),
			.S(gen[1490]),
			.SE(gen[1491]),

			.SELF(gen[1430]),
			.cell_state(gen[1430])
		); 

/******************* CELL 1431 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1431 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1370]),
			.N(gen[1371]),
			.NE(gen[1372]),

			.O(gen[1430]),
			.E(gen[1432]),

			.SO(gen[1490]),
			.S(gen[1491]),
			.SE(gen[1492]),

			.SELF(gen[1431]),
			.cell_state(gen[1431])
		); 

/******************* CELL 1432 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1432 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1371]),
			.N(gen[1372]),
			.NE(gen[1373]),

			.O(gen[1431]),
			.E(gen[1433]),

			.SO(gen[1491]),
			.S(gen[1492]),
			.SE(gen[1493]),

			.SELF(gen[1432]),
			.cell_state(gen[1432])
		); 

/******************* CELL 1433 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1433 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1372]),
			.N(gen[1373]),
			.NE(gen[1374]),

			.O(gen[1432]),
			.E(gen[1434]),

			.SO(gen[1492]),
			.S(gen[1493]),
			.SE(gen[1494]),

			.SELF(gen[1433]),
			.cell_state(gen[1433])
		); 

/******************* CELL 1434 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1434 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1373]),
			.N(gen[1374]),
			.NE(gen[1375]),

			.O(gen[1433]),
			.E(gen[1435]),

			.SO(gen[1493]),
			.S(gen[1494]),
			.SE(gen[1495]),

			.SELF(gen[1434]),
			.cell_state(gen[1434])
		); 

/******************* CELL 1435 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1435 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1374]),
			.N(gen[1375]),
			.NE(gen[1376]),

			.O(gen[1434]),
			.E(gen[1436]),

			.SO(gen[1494]),
			.S(gen[1495]),
			.SE(gen[1496]),

			.SELF(gen[1435]),
			.cell_state(gen[1435])
		); 

/******************* CELL 1436 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1436 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1375]),
			.N(gen[1376]),
			.NE(gen[1377]),

			.O(gen[1435]),
			.E(gen[1437]),

			.SO(gen[1495]),
			.S(gen[1496]),
			.SE(gen[1497]),

			.SELF(gen[1436]),
			.cell_state(gen[1436])
		); 

/******************* CELL 1437 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1437 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1376]),
			.N(gen[1377]),
			.NE(gen[1378]),

			.O(gen[1436]),
			.E(gen[1438]),

			.SO(gen[1496]),
			.S(gen[1497]),
			.SE(gen[1498]),

			.SELF(gen[1437]),
			.cell_state(gen[1437])
		); 

/******************* CELL 1438 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1438 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1377]),
			.N(gen[1378]),
			.NE(gen[1379]),

			.O(gen[1437]),
			.E(gen[1439]),

			.SO(gen[1497]),
			.S(gen[1498]),
			.SE(gen[1499]),

			.SELF(gen[1438]),
			.cell_state(gen[1438])
		); 

/******************* CELL 1439 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1439 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1378]),
			.N(gen[1379]),
			.NE(gen[1378]),

			.O(gen[1438]),
			.E(gen[1438]),

			.SO(gen[1498]),
			.S(gen[1499]),
			.SE(gen[1498]),

			.SELF(gen[1439]),
			.cell_state(gen[1439])
		); 

/******************* CELL 1440 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1440 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1381]),
			.N(gen[1380]),
			.NE(gen[1381]),

			.O(gen[1441]),
			.E(gen[1441]),

			.SO(gen[1501]),
			.S(gen[1500]),
			.SE(gen[1501]),

			.SELF(gen[1440]),
			.cell_state(gen[1440])
		); 

/******************* CELL 1441 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1441 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1380]),
			.N(gen[1381]),
			.NE(gen[1382]),

			.O(gen[1440]),
			.E(gen[1442]),

			.SO(gen[1500]),
			.S(gen[1501]),
			.SE(gen[1502]),

			.SELF(gen[1441]),
			.cell_state(gen[1441])
		); 

/******************* CELL 1442 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1442 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1381]),
			.N(gen[1382]),
			.NE(gen[1383]),

			.O(gen[1441]),
			.E(gen[1443]),

			.SO(gen[1501]),
			.S(gen[1502]),
			.SE(gen[1503]),

			.SELF(gen[1442]),
			.cell_state(gen[1442])
		); 

/******************* CELL 1443 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1443 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1382]),
			.N(gen[1383]),
			.NE(gen[1384]),

			.O(gen[1442]),
			.E(gen[1444]),

			.SO(gen[1502]),
			.S(gen[1503]),
			.SE(gen[1504]),

			.SELF(gen[1443]),
			.cell_state(gen[1443])
		); 

/******************* CELL 1444 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1444 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1383]),
			.N(gen[1384]),
			.NE(gen[1385]),

			.O(gen[1443]),
			.E(gen[1445]),

			.SO(gen[1503]),
			.S(gen[1504]),
			.SE(gen[1505]),

			.SELF(gen[1444]),
			.cell_state(gen[1444])
		); 

/******************* CELL 1445 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1445 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1384]),
			.N(gen[1385]),
			.NE(gen[1386]),

			.O(gen[1444]),
			.E(gen[1446]),

			.SO(gen[1504]),
			.S(gen[1505]),
			.SE(gen[1506]),

			.SELF(gen[1445]),
			.cell_state(gen[1445])
		); 

/******************* CELL 1446 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1446 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1385]),
			.N(gen[1386]),
			.NE(gen[1387]),

			.O(gen[1445]),
			.E(gen[1447]),

			.SO(gen[1505]),
			.S(gen[1506]),
			.SE(gen[1507]),

			.SELF(gen[1446]),
			.cell_state(gen[1446])
		); 

/******************* CELL 1447 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1447 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1386]),
			.N(gen[1387]),
			.NE(gen[1388]),

			.O(gen[1446]),
			.E(gen[1448]),

			.SO(gen[1506]),
			.S(gen[1507]),
			.SE(gen[1508]),

			.SELF(gen[1447]),
			.cell_state(gen[1447])
		); 

/******************* CELL 1448 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1448 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1387]),
			.N(gen[1388]),
			.NE(gen[1389]),

			.O(gen[1447]),
			.E(gen[1449]),

			.SO(gen[1507]),
			.S(gen[1508]),
			.SE(gen[1509]),

			.SELF(gen[1448]),
			.cell_state(gen[1448])
		); 

/******************* CELL 1449 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1449 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1388]),
			.N(gen[1389]),
			.NE(gen[1390]),

			.O(gen[1448]),
			.E(gen[1450]),

			.SO(gen[1508]),
			.S(gen[1509]),
			.SE(gen[1510]),

			.SELF(gen[1449]),
			.cell_state(gen[1449])
		); 

/******************* CELL 1450 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1450 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1389]),
			.N(gen[1390]),
			.NE(gen[1391]),

			.O(gen[1449]),
			.E(gen[1451]),

			.SO(gen[1509]),
			.S(gen[1510]),
			.SE(gen[1511]),

			.SELF(gen[1450]),
			.cell_state(gen[1450])
		); 

/******************* CELL 1451 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1451 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1390]),
			.N(gen[1391]),
			.NE(gen[1392]),

			.O(gen[1450]),
			.E(gen[1452]),

			.SO(gen[1510]),
			.S(gen[1511]),
			.SE(gen[1512]),

			.SELF(gen[1451]),
			.cell_state(gen[1451])
		); 

/******************* CELL 1452 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1452 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1391]),
			.N(gen[1392]),
			.NE(gen[1393]),

			.O(gen[1451]),
			.E(gen[1453]),

			.SO(gen[1511]),
			.S(gen[1512]),
			.SE(gen[1513]),

			.SELF(gen[1452]),
			.cell_state(gen[1452])
		); 

/******************* CELL 1453 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1453 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1392]),
			.N(gen[1393]),
			.NE(gen[1394]),

			.O(gen[1452]),
			.E(gen[1454]),

			.SO(gen[1512]),
			.S(gen[1513]),
			.SE(gen[1514]),

			.SELF(gen[1453]),
			.cell_state(gen[1453])
		); 

/******************* CELL 1454 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1454 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1393]),
			.N(gen[1394]),
			.NE(gen[1395]),

			.O(gen[1453]),
			.E(gen[1455]),

			.SO(gen[1513]),
			.S(gen[1514]),
			.SE(gen[1515]),

			.SELF(gen[1454]),
			.cell_state(gen[1454])
		); 

/******************* CELL 1455 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1455 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1394]),
			.N(gen[1395]),
			.NE(gen[1396]),

			.O(gen[1454]),
			.E(gen[1456]),

			.SO(gen[1514]),
			.S(gen[1515]),
			.SE(gen[1516]),

			.SELF(gen[1455]),
			.cell_state(gen[1455])
		); 

/******************* CELL 1456 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1456 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1395]),
			.N(gen[1396]),
			.NE(gen[1397]),

			.O(gen[1455]),
			.E(gen[1457]),

			.SO(gen[1515]),
			.S(gen[1516]),
			.SE(gen[1517]),

			.SELF(gen[1456]),
			.cell_state(gen[1456])
		); 

/******************* CELL 1457 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1457 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1396]),
			.N(gen[1397]),
			.NE(gen[1398]),

			.O(gen[1456]),
			.E(gen[1458]),

			.SO(gen[1516]),
			.S(gen[1517]),
			.SE(gen[1518]),

			.SELF(gen[1457]),
			.cell_state(gen[1457])
		); 

/******************* CELL 1458 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1458 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1397]),
			.N(gen[1398]),
			.NE(gen[1399]),

			.O(gen[1457]),
			.E(gen[1459]),

			.SO(gen[1517]),
			.S(gen[1518]),
			.SE(gen[1519]),

			.SELF(gen[1458]),
			.cell_state(gen[1458])
		); 

/******************* CELL 1459 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1459 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1398]),
			.N(gen[1399]),
			.NE(gen[1400]),

			.O(gen[1458]),
			.E(gen[1460]),

			.SO(gen[1518]),
			.S(gen[1519]),
			.SE(gen[1520]),

			.SELF(gen[1459]),
			.cell_state(gen[1459])
		); 

/******************* CELL 1460 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1460 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1399]),
			.N(gen[1400]),
			.NE(gen[1401]),

			.O(gen[1459]),
			.E(gen[1461]),

			.SO(gen[1519]),
			.S(gen[1520]),
			.SE(gen[1521]),

			.SELF(gen[1460]),
			.cell_state(gen[1460])
		); 

/******************* CELL 1461 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1461 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1400]),
			.N(gen[1401]),
			.NE(gen[1402]),

			.O(gen[1460]),
			.E(gen[1462]),

			.SO(gen[1520]),
			.S(gen[1521]),
			.SE(gen[1522]),

			.SELF(gen[1461]),
			.cell_state(gen[1461])
		); 

/******************* CELL 1462 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1462 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1401]),
			.N(gen[1402]),
			.NE(gen[1403]),

			.O(gen[1461]),
			.E(gen[1463]),

			.SO(gen[1521]),
			.S(gen[1522]),
			.SE(gen[1523]),

			.SELF(gen[1462]),
			.cell_state(gen[1462])
		); 

/******************* CELL 1463 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1463 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1402]),
			.N(gen[1403]),
			.NE(gen[1404]),

			.O(gen[1462]),
			.E(gen[1464]),

			.SO(gen[1522]),
			.S(gen[1523]),
			.SE(gen[1524]),

			.SELF(gen[1463]),
			.cell_state(gen[1463])
		); 

/******************* CELL 1464 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1464 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1403]),
			.N(gen[1404]),
			.NE(gen[1405]),

			.O(gen[1463]),
			.E(gen[1465]),

			.SO(gen[1523]),
			.S(gen[1524]),
			.SE(gen[1525]),

			.SELF(gen[1464]),
			.cell_state(gen[1464])
		); 

/******************* CELL 1465 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1465 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1404]),
			.N(gen[1405]),
			.NE(gen[1406]),

			.O(gen[1464]),
			.E(gen[1466]),

			.SO(gen[1524]),
			.S(gen[1525]),
			.SE(gen[1526]),

			.SELF(gen[1465]),
			.cell_state(gen[1465])
		); 

/******************* CELL 1466 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1466 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1405]),
			.N(gen[1406]),
			.NE(gen[1407]),

			.O(gen[1465]),
			.E(gen[1467]),

			.SO(gen[1525]),
			.S(gen[1526]),
			.SE(gen[1527]),

			.SELF(gen[1466]),
			.cell_state(gen[1466])
		); 

/******************* CELL 1467 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1467 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1406]),
			.N(gen[1407]),
			.NE(gen[1408]),

			.O(gen[1466]),
			.E(gen[1468]),

			.SO(gen[1526]),
			.S(gen[1527]),
			.SE(gen[1528]),

			.SELF(gen[1467]),
			.cell_state(gen[1467])
		); 

/******************* CELL 1468 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1468 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1407]),
			.N(gen[1408]),
			.NE(gen[1409]),

			.O(gen[1467]),
			.E(gen[1469]),

			.SO(gen[1527]),
			.S(gen[1528]),
			.SE(gen[1529]),

			.SELF(gen[1468]),
			.cell_state(gen[1468])
		); 

/******************* CELL 1469 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1469 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1408]),
			.N(gen[1409]),
			.NE(gen[1410]),

			.O(gen[1468]),
			.E(gen[1470]),

			.SO(gen[1528]),
			.S(gen[1529]),
			.SE(gen[1530]),

			.SELF(gen[1469]),
			.cell_state(gen[1469])
		); 

/******************* CELL 1470 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1470 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1409]),
			.N(gen[1410]),
			.NE(gen[1411]),

			.O(gen[1469]),
			.E(gen[1471]),

			.SO(gen[1529]),
			.S(gen[1530]),
			.SE(gen[1531]),

			.SELF(gen[1470]),
			.cell_state(gen[1470])
		); 

/******************* CELL 1471 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1471 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1410]),
			.N(gen[1411]),
			.NE(gen[1412]),

			.O(gen[1470]),
			.E(gen[1472]),

			.SO(gen[1530]),
			.S(gen[1531]),
			.SE(gen[1532]),

			.SELF(gen[1471]),
			.cell_state(gen[1471])
		); 

/******************* CELL 1472 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1472 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1411]),
			.N(gen[1412]),
			.NE(gen[1413]),

			.O(gen[1471]),
			.E(gen[1473]),

			.SO(gen[1531]),
			.S(gen[1532]),
			.SE(gen[1533]),

			.SELF(gen[1472]),
			.cell_state(gen[1472])
		); 

/******************* CELL 1473 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1473 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1412]),
			.N(gen[1413]),
			.NE(gen[1414]),

			.O(gen[1472]),
			.E(gen[1474]),

			.SO(gen[1532]),
			.S(gen[1533]),
			.SE(gen[1534]),

			.SELF(gen[1473]),
			.cell_state(gen[1473])
		); 

/******************* CELL 1474 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1474 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1413]),
			.N(gen[1414]),
			.NE(gen[1415]),

			.O(gen[1473]),
			.E(gen[1475]),

			.SO(gen[1533]),
			.S(gen[1534]),
			.SE(gen[1535]),

			.SELF(gen[1474]),
			.cell_state(gen[1474])
		); 

/******************* CELL 1475 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1475 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1414]),
			.N(gen[1415]),
			.NE(gen[1416]),

			.O(gen[1474]),
			.E(gen[1476]),

			.SO(gen[1534]),
			.S(gen[1535]),
			.SE(gen[1536]),

			.SELF(gen[1475]),
			.cell_state(gen[1475])
		); 

/******************* CELL 1476 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1476 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1415]),
			.N(gen[1416]),
			.NE(gen[1417]),

			.O(gen[1475]),
			.E(gen[1477]),

			.SO(gen[1535]),
			.S(gen[1536]),
			.SE(gen[1537]),

			.SELF(gen[1476]),
			.cell_state(gen[1476])
		); 

/******************* CELL 1477 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1477 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1416]),
			.N(gen[1417]),
			.NE(gen[1418]),

			.O(gen[1476]),
			.E(gen[1478]),

			.SO(gen[1536]),
			.S(gen[1537]),
			.SE(gen[1538]),

			.SELF(gen[1477]),
			.cell_state(gen[1477])
		); 

/******************* CELL 1478 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1478 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1417]),
			.N(gen[1418]),
			.NE(gen[1419]),

			.O(gen[1477]),
			.E(gen[1479]),

			.SO(gen[1537]),
			.S(gen[1538]),
			.SE(gen[1539]),

			.SELF(gen[1478]),
			.cell_state(gen[1478])
		); 

/******************* CELL 1479 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1479 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1418]),
			.N(gen[1419]),
			.NE(gen[1420]),

			.O(gen[1478]),
			.E(gen[1480]),

			.SO(gen[1538]),
			.S(gen[1539]),
			.SE(gen[1540]),

			.SELF(gen[1479]),
			.cell_state(gen[1479])
		); 

/******************* CELL 1480 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1480 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1419]),
			.N(gen[1420]),
			.NE(gen[1421]),

			.O(gen[1479]),
			.E(gen[1481]),

			.SO(gen[1539]),
			.S(gen[1540]),
			.SE(gen[1541]),

			.SELF(gen[1480]),
			.cell_state(gen[1480])
		); 

/******************* CELL 1481 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1481 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1420]),
			.N(gen[1421]),
			.NE(gen[1422]),

			.O(gen[1480]),
			.E(gen[1482]),

			.SO(gen[1540]),
			.S(gen[1541]),
			.SE(gen[1542]),

			.SELF(gen[1481]),
			.cell_state(gen[1481])
		); 

/******************* CELL 1482 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1482 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1421]),
			.N(gen[1422]),
			.NE(gen[1423]),

			.O(gen[1481]),
			.E(gen[1483]),

			.SO(gen[1541]),
			.S(gen[1542]),
			.SE(gen[1543]),

			.SELF(gen[1482]),
			.cell_state(gen[1482])
		); 

/******************* CELL 1483 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1483 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1422]),
			.N(gen[1423]),
			.NE(gen[1424]),

			.O(gen[1482]),
			.E(gen[1484]),

			.SO(gen[1542]),
			.S(gen[1543]),
			.SE(gen[1544]),

			.SELF(gen[1483]),
			.cell_state(gen[1483])
		); 

/******************* CELL 1484 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1484 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1423]),
			.N(gen[1424]),
			.NE(gen[1425]),

			.O(gen[1483]),
			.E(gen[1485]),

			.SO(gen[1543]),
			.S(gen[1544]),
			.SE(gen[1545]),

			.SELF(gen[1484]),
			.cell_state(gen[1484])
		); 

/******************* CELL 1485 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1485 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1424]),
			.N(gen[1425]),
			.NE(gen[1426]),

			.O(gen[1484]),
			.E(gen[1486]),

			.SO(gen[1544]),
			.S(gen[1545]),
			.SE(gen[1546]),

			.SELF(gen[1485]),
			.cell_state(gen[1485])
		); 

/******************* CELL 1486 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1486 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1425]),
			.N(gen[1426]),
			.NE(gen[1427]),

			.O(gen[1485]),
			.E(gen[1487]),

			.SO(gen[1545]),
			.S(gen[1546]),
			.SE(gen[1547]),

			.SELF(gen[1486]),
			.cell_state(gen[1486])
		); 

/******************* CELL 1487 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1487 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1426]),
			.N(gen[1427]),
			.NE(gen[1428]),

			.O(gen[1486]),
			.E(gen[1488]),

			.SO(gen[1546]),
			.S(gen[1547]),
			.SE(gen[1548]),

			.SELF(gen[1487]),
			.cell_state(gen[1487])
		); 

/******************* CELL 1488 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1488 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1427]),
			.N(gen[1428]),
			.NE(gen[1429]),

			.O(gen[1487]),
			.E(gen[1489]),

			.SO(gen[1547]),
			.S(gen[1548]),
			.SE(gen[1549]),

			.SELF(gen[1488]),
			.cell_state(gen[1488])
		); 

/******************* CELL 1489 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1489 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1428]),
			.N(gen[1429]),
			.NE(gen[1430]),

			.O(gen[1488]),
			.E(gen[1490]),

			.SO(gen[1548]),
			.S(gen[1549]),
			.SE(gen[1550]),

			.SELF(gen[1489]),
			.cell_state(gen[1489])
		); 

/******************* CELL 1490 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1490 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1429]),
			.N(gen[1430]),
			.NE(gen[1431]),

			.O(gen[1489]),
			.E(gen[1491]),

			.SO(gen[1549]),
			.S(gen[1550]),
			.SE(gen[1551]),

			.SELF(gen[1490]),
			.cell_state(gen[1490])
		); 

/******************* CELL 1491 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1491 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1430]),
			.N(gen[1431]),
			.NE(gen[1432]),

			.O(gen[1490]),
			.E(gen[1492]),

			.SO(gen[1550]),
			.S(gen[1551]),
			.SE(gen[1552]),

			.SELF(gen[1491]),
			.cell_state(gen[1491])
		); 

/******************* CELL 1492 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1492 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1431]),
			.N(gen[1432]),
			.NE(gen[1433]),

			.O(gen[1491]),
			.E(gen[1493]),

			.SO(gen[1551]),
			.S(gen[1552]),
			.SE(gen[1553]),

			.SELF(gen[1492]),
			.cell_state(gen[1492])
		); 

/******************* CELL 1493 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1493 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1432]),
			.N(gen[1433]),
			.NE(gen[1434]),

			.O(gen[1492]),
			.E(gen[1494]),

			.SO(gen[1552]),
			.S(gen[1553]),
			.SE(gen[1554]),

			.SELF(gen[1493]),
			.cell_state(gen[1493])
		); 

/******************* CELL 1494 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1494 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1433]),
			.N(gen[1434]),
			.NE(gen[1435]),

			.O(gen[1493]),
			.E(gen[1495]),

			.SO(gen[1553]),
			.S(gen[1554]),
			.SE(gen[1555]),

			.SELF(gen[1494]),
			.cell_state(gen[1494])
		); 

/******************* CELL 1495 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1495 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1434]),
			.N(gen[1435]),
			.NE(gen[1436]),

			.O(gen[1494]),
			.E(gen[1496]),

			.SO(gen[1554]),
			.S(gen[1555]),
			.SE(gen[1556]),

			.SELF(gen[1495]),
			.cell_state(gen[1495])
		); 

/******************* CELL 1496 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1496 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1435]),
			.N(gen[1436]),
			.NE(gen[1437]),

			.O(gen[1495]),
			.E(gen[1497]),

			.SO(gen[1555]),
			.S(gen[1556]),
			.SE(gen[1557]),

			.SELF(gen[1496]),
			.cell_state(gen[1496])
		); 

/******************* CELL 1497 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1497 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1436]),
			.N(gen[1437]),
			.NE(gen[1438]),

			.O(gen[1496]),
			.E(gen[1498]),

			.SO(gen[1556]),
			.S(gen[1557]),
			.SE(gen[1558]),

			.SELF(gen[1497]),
			.cell_state(gen[1497])
		); 

/******************* CELL 1498 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1498 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1437]),
			.N(gen[1438]),
			.NE(gen[1439]),

			.O(gen[1497]),
			.E(gen[1499]),

			.SO(gen[1557]),
			.S(gen[1558]),
			.SE(gen[1559]),

			.SELF(gen[1498]),
			.cell_state(gen[1498])
		); 

/******************* CELL 1499 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1499 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1438]),
			.N(gen[1439]),
			.NE(gen[1438]),

			.O(gen[1498]),
			.E(gen[1498]),

			.SO(gen[1558]),
			.S(gen[1559]),
			.SE(gen[1558]),

			.SELF(gen[1499]),
			.cell_state(gen[1499])
		); 

/******************* CELL 1500 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1500 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1441]),
			.N(gen[1440]),
			.NE(gen[1441]),

			.O(gen[1501]),
			.E(gen[1501]),

			.SO(gen[1561]),
			.S(gen[1560]),
			.SE(gen[1561]),

			.SELF(gen[1500]),
			.cell_state(gen[1500])
		); 

/******************* CELL 1501 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1501 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1440]),
			.N(gen[1441]),
			.NE(gen[1442]),

			.O(gen[1500]),
			.E(gen[1502]),

			.SO(gen[1560]),
			.S(gen[1561]),
			.SE(gen[1562]),

			.SELF(gen[1501]),
			.cell_state(gen[1501])
		); 

/******************* CELL 1502 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1502 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1441]),
			.N(gen[1442]),
			.NE(gen[1443]),

			.O(gen[1501]),
			.E(gen[1503]),

			.SO(gen[1561]),
			.S(gen[1562]),
			.SE(gen[1563]),

			.SELF(gen[1502]),
			.cell_state(gen[1502])
		); 

/******************* CELL 1503 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1503 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1442]),
			.N(gen[1443]),
			.NE(gen[1444]),

			.O(gen[1502]),
			.E(gen[1504]),

			.SO(gen[1562]),
			.S(gen[1563]),
			.SE(gen[1564]),

			.SELF(gen[1503]),
			.cell_state(gen[1503])
		); 

/******************* CELL 1504 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1504 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1443]),
			.N(gen[1444]),
			.NE(gen[1445]),

			.O(gen[1503]),
			.E(gen[1505]),

			.SO(gen[1563]),
			.S(gen[1564]),
			.SE(gen[1565]),

			.SELF(gen[1504]),
			.cell_state(gen[1504])
		); 

/******************* CELL 1505 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1505 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1444]),
			.N(gen[1445]),
			.NE(gen[1446]),

			.O(gen[1504]),
			.E(gen[1506]),

			.SO(gen[1564]),
			.S(gen[1565]),
			.SE(gen[1566]),

			.SELF(gen[1505]),
			.cell_state(gen[1505])
		); 

/******************* CELL 1506 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1506 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1445]),
			.N(gen[1446]),
			.NE(gen[1447]),

			.O(gen[1505]),
			.E(gen[1507]),

			.SO(gen[1565]),
			.S(gen[1566]),
			.SE(gen[1567]),

			.SELF(gen[1506]),
			.cell_state(gen[1506])
		); 

/******************* CELL 1507 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1507 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1446]),
			.N(gen[1447]),
			.NE(gen[1448]),

			.O(gen[1506]),
			.E(gen[1508]),

			.SO(gen[1566]),
			.S(gen[1567]),
			.SE(gen[1568]),

			.SELF(gen[1507]),
			.cell_state(gen[1507])
		); 

/******************* CELL 1508 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1508 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1447]),
			.N(gen[1448]),
			.NE(gen[1449]),

			.O(gen[1507]),
			.E(gen[1509]),

			.SO(gen[1567]),
			.S(gen[1568]),
			.SE(gen[1569]),

			.SELF(gen[1508]),
			.cell_state(gen[1508])
		); 

/******************* CELL 1509 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1509 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1448]),
			.N(gen[1449]),
			.NE(gen[1450]),

			.O(gen[1508]),
			.E(gen[1510]),

			.SO(gen[1568]),
			.S(gen[1569]),
			.SE(gen[1570]),

			.SELF(gen[1509]),
			.cell_state(gen[1509])
		); 

/******************* CELL 1510 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1510 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1449]),
			.N(gen[1450]),
			.NE(gen[1451]),

			.O(gen[1509]),
			.E(gen[1511]),

			.SO(gen[1569]),
			.S(gen[1570]),
			.SE(gen[1571]),

			.SELF(gen[1510]),
			.cell_state(gen[1510])
		); 

/******************* CELL 1511 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1511 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1450]),
			.N(gen[1451]),
			.NE(gen[1452]),

			.O(gen[1510]),
			.E(gen[1512]),

			.SO(gen[1570]),
			.S(gen[1571]),
			.SE(gen[1572]),

			.SELF(gen[1511]),
			.cell_state(gen[1511])
		); 

/******************* CELL 1512 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1512 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1451]),
			.N(gen[1452]),
			.NE(gen[1453]),

			.O(gen[1511]),
			.E(gen[1513]),

			.SO(gen[1571]),
			.S(gen[1572]),
			.SE(gen[1573]),

			.SELF(gen[1512]),
			.cell_state(gen[1512])
		); 

/******************* CELL 1513 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1513 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1452]),
			.N(gen[1453]),
			.NE(gen[1454]),

			.O(gen[1512]),
			.E(gen[1514]),

			.SO(gen[1572]),
			.S(gen[1573]),
			.SE(gen[1574]),

			.SELF(gen[1513]),
			.cell_state(gen[1513])
		); 

/******************* CELL 1514 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1514 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1453]),
			.N(gen[1454]),
			.NE(gen[1455]),

			.O(gen[1513]),
			.E(gen[1515]),

			.SO(gen[1573]),
			.S(gen[1574]),
			.SE(gen[1575]),

			.SELF(gen[1514]),
			.cell_state(gen[1514])
		); 

/******************* CELL 1515 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1515 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1454]),
			.N(gen[1455]),
			.NE(gen[1456]),

			.O(gen[1514]),
			.E(gen[1516]),

			.SO(gen[1574]),
			.S(gen[1575]),
			.SE(gen[1576]),

			.SELF(gen[1515]),
			.cell_state(gen[1515])
		); 

/******************* CELL 1516 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1516 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1455]),
			.N(gen[1456]),
			.NE(gen[1457]),

			.O(gen[1515]),
			.E(gen[1517]),

			.SO(gen[1575]),
			.S(gen[1576]),
			.SE(gen[1577]),

			.SELF(gen[1516]),
			.cell_state(gen[1516])
		); 

/******************* CELL 1517 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1517 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1456]),
			.N(gen[1457]),
			.NE(gen[1458]),

			.O(gen[1516]),
			.E(gen[1518]),

			.SO(gen[1576]),
			.S(gen[1577]),
			.SE(gen[1578]),

			.SELF(gen[1517]),
			.cell_state(gen[1517])
		); 

/******************* CELL 1518 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1518 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1457]),
			.N(gen[1458]),
			.NE(gen[1459]),

			.O(gen[1517]),
			.E(gen[1519]),

			.SO(gen[1577]),
			.S(gen[1578]),
			.SE(gen[1579]),

			.SELF(gen[1518]),
			.cell_state(gen[1518])
		); 

/******************* CELL 1519 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1519 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1458]),
			.N(gen[1459]),
			.NE(gen[1460]),

			.O(gen[1518]),
			.E(gen[1520]),

			.SO(gen[1578]),
			.S(gen[1579]),
			.SE(gen[1580]),

			.SELF(gen[1519]),
			.cell_state(gen[1519])
		); 

/******************* CELL 1520 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1520 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1459]),
			.N(gen[1460]),
			.NE(gen[1461]),

			.O(gen[1519]),
			.E(gen[1521]),

			.SO(gen[1579]),
			.S(gen[1580]),
			.SE(gen[1581]),

			.SELF(gen[1520]),
			.cell_state(gen[1520])
		); 

/******************* CELL 1521 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1521 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1460]),
			.N(gen[1461]),
			.NE(gen[1462]),

			.O(gen[1520]),
			.E(gen[1522]),

			.SO(gen[1580]),
			.S(gen[1581]),
			.SE(gen[1582]),

			.SELF(gen[1521]),
			.cell_state(gen[1521])
		); 

/******************* CELL 1522 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1522 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1461]),
			.N(gen[1462]),
			.NE(gen[1463]),

			.O(gen[1521]),
			.E(gen[1523]),

			.SO(gen[1581]),
			.S(gen[1582]),
			.SE(gen[1583]),

			.SELF(gen[1522]),
			.cell_state(gen[1522])
		); 

/******************* CELL 1523 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1523 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1462]),
			.N(gen[1463]),
			.NE(gen[1464]),

			.O(gen[1522]),
			.E(gen[1524]),

			.SO(gen[1582]),
			.S(gen[1583]),
			.SE(gen[1584]),

			.SELF(gen[1523]),
			.cell_state(gen[1523])
		); 

/******************* CELL 1524 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1524 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1463]),
			.N(gen[1464]),
			.NE(gen[1465]),

			.O(gen[1523]),
			.E(gen[1525]),

			.SO(gen[1583]),
			.S(gen[1584]),
			.SE(gen[1585]),

			.SELF(gen[1524]),
			.cell_state(gen[1524])
		); 

/******************* CELL 1525 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1525 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1464]),
			.N(gen[1465]),
			.NE(gen[1466]),

			.O(gen[1524]),
			.E(gen[1526]),

			.SO(gen[1584]),
			.S(gen[1585]),
			.SE(gen[1586]),

			.SELF(gen[1525]),
			.cell_state(gen[1525])
		); 

/******************* CELL 1526 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1526 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1465]),
			.N(gen[1466]),
			.NE(gen[1467]),

			.O(gen[1525]),
			.E(gen[1527]),

			.SO(gen[1585]),
			.S(gen[1586]),
			.SE(gen[1587]),

			.SELF(gen[1526]),
			.cell_state(gen[1526])
		); 

/******************* CELL 1527 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1527 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1466]),
			.N(gen[1467]),
			.NE(gen[1468]),

			.O(gen[1526]),
			.E(gen[1528]),

			.SO(gen[1586]),
			.S(gen[1587]),
			.SE(gen[1588]),

			.SELF(gen[1527]),
			.cell_state(gen[1527])
		); 

/******************* CELL 1528 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1528 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1467]),
			.N(gen[1468]),
			.NE(gen[1469]),

			.O(gen[1527]),
			.E(gen[1529]),

			.SO(gen[1587]),
			.S(gen[1588]),
			.SE(gen[1589]),

			.SELF(gen[1528]),
			.cell_state(gen[1528])
		); 

/******************* CELL 1529 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1529 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1468]),
			.N(gen[1469]),
			.NE(gen[1470]),

			.O(gen[1528]),
			.E(gen[1530]),

			.SO(gen[1588]),
			.S(gen[1589]),
			.SE(gen[1590]),

			.SELF(gen[1529]),
			.cell_state(gen[1529])
		); 

/******************* CELL 1530 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1530 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1469]),
			.N(gen[1470]),
			.NE(gen[1471]),

			.O(gen[1529]),
			.E(gen[1531]),

			.SO(gen[1589]),
			.S(gen[1590]),
			.SE(gen[1591]),

			.SELF(gen[1530]),
			.cell_state(gen[1530])
		); 

/******************* CELL 1531 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1531 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1470]),
			.N(gen[1471]),
			.NE(gen[1472]),

			.O(gen[1530]),
			.E(gen[1532]),

			.SO(gen[1590]),
			.S(gen[1591]),
			.SE(gen[1592]),

			.SELF(gen[1531]),
			.cell_state(gen[1531])
		); 

/******************* CELL 1532 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1532 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1471]),
			.N(gen[1472]),
			.NE(gen[1473]),

			.O(gen[1531]),
			.E(gen[1533]),

			.SO(gen[1591]),
			.S(gen[1592]),
			.SE(gen[1593]),

			.SELF(gen[1532]),
			.cell_state(gen[1532])
		); 

/******************* CELL 1533 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1533 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1472]),
			.N(gen[1473]),
			.NE(gen[1474]),

			.O(gen[1532]),
			.E(gen[1534]),

			.SO(gen[1592]),
			.S(gen[1593]),
			.SE(gen[1594]),

			.SELF(gen[1533]),
			.cell_state(gen[1533])
		); 

/******************* CELL 1534 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1534 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1473]),
			.N(gen[1474]),
			.NE(gen[1475]),

			.O(gen[1533]),
			.E(gen[1535]),

			.SO(gen[1593]),
			.S(gen[1594]),
			.SE(gen[1595]),

			.SELF(gen[1534]),
			.cell_state(gen[1534])
		); 

/******************* CELL 1535 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1535 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1474]),
			.N(gen[1475]),
			.NE(gen[1476]),

			.O(gen[1534]),
			.E(gen[1536]),

			.SO(gen[1594]),
			.S(gen[1595]),
			.SE(gen[1596]),

			.SELF(gen[1535]),
			.cell_state(gen[1535])
		); 

/******************* CELL 1536 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1536 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1475]),
			.N(gen[1476]),
			.NE(gen[1477]),

			.O(gen[1535]),
			.E(gen[1537]),

			.SO(gen[1595]),
			.S(gen[1596]),
			.SE(gen[1597]),

			.SELF(gen[1536]),
			.cell_state(gen[1536])
		); 

/******************* CELL 1537 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1537 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1476]),
			.N(gen[1477]),
			.NE(gen[1478]),

			.O(gen[1536]),
			.E(gen[1538]),

			.SO(gen[1596]),
			.S(gen[1597]),
			.SE(gen[1598]),

			.SELF(gen[1537]),
			.cell_state(gen[1537])
		); 

/******************* CELL 1538 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1538 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1477]),
			.N(gen[1478]),
			.NE(gen[1479]),

			.O(gen[1537]),
			.E(gen[1539]),

			.SO(gen[1597]),
			.S(gen[1598]),
			.SE(gen[1599]),

			.SELF(gen[1538]),
			.cell_state(gen[1538])
		); 

/******************* CELL 1539 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1539 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1478]),
			.N(gen[1479]),
			.NE(gen[1480]),

			.O(gen[1538]),
			.E(gen[1540]),

			.SO(gen[1598]),
			.S(gen[1599]),
			.SE(gen[1600]),

			.SELF(gen[1539]),
			.cell_state(gen[1539])
		); 

/******************* CELL 1540 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1540 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1479]),
			.N(gen[1480]),
			.NE(gen[1481]),

			.O(gen[1539]),
			.E(gen[1541]),

			.SO(gen[1599]),
			.S(gen[1600]),
			.SE(gen[1601]),

			.SELF(gen[1540]),
			.cell_state(gen[1540])
		); 

/******************* CELL 1541 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1541 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1480]),
			.N(gen[1481]),
			.NE(gen[1482]),

			.O(gen[1540]),
			.E(gen[1542]),

			.SO(gen[1600]),
			.S(gen[1601]),
			.SE(gen[1602]),

			.SELF(gen[1541]),
			.cell_state(gen[1541])
		); 

/******************* CELL 1542 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1542 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1481]),
			.N(gen[1482]),
			.NE(gen[1483]),

			.O(gen[1541]),
			.E(gen[1543]),

			.SO(gen[1601]),
			.S(gen[1602]),
			.SE(gen[1603]),

			.SELF(gen[1542]),
			.cell_state(gen[1542])
		); 

/******************* CELL 1543 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1543 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1482]),
			.N(gen[1483]),
			.NE(gen[1484]),

			.O(gen[1542]),
			.E(gen[1544]),

			.SO(gen[1602]),
			.S(gen[1603]),
			.SE(gen[1604]),

			.SELF(gen[1543]),
			.cell_state(gen[1543])
		); 

/******************* CELL 1544 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1544 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1483]),
			.N(gen[1484]),
			.NE(gen[1485]),

			.O(gen[1543]),
			.E(gen[1545]),

			.SO(gen[1603]),
			.S(gen[1604]),
			.SE(gen[1605]),

			.SELF(gen[1544]),
			.cell_state(gen[1544])
		); 

/******************* CELL 1545 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1545 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1484]),
			.N(gen[1485]),
			.NE(gen[1486]),

			.O(gen[1544]),
			.E(gen[1546]),

			.SO(gen[1604]),
			.S(gen[1605]),
			.SE(gen[1606]),

			.SELF(gen[1545]),
			.cell_state(gen[1545])
		); 

/******************* CELL 1546 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1546 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1485]),
			.N(gen[1486]),
			.NE(gen[1487]),

			.O(gen[1545]),
			.E(gen[1547]),

			.SO(gen[1605]),
			.S(gen[1606]),
			.SE(gen[1607]),

			.SELF(gen[1546]),
			.cell_state(gen[1546])
		); 

/******************* CELL 1547 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1547 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1486]),
			.N(gen[1487]),
			.NE(gen[1488]),

			.O(gen[1546]),
			.E(gen[1548]),

			.SO(gen[1606]),
			.S(gen[1607]),
			.SE(gen[1608]),

			.SELF(gen[1547]),
			.cell_state(gen[1547])
		); 

/******************* CELL 1548 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1548 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1487]),
			.N(gen[1488]),
			.NE(gen[1489]),

			.O(gen[1547]),
			.E(gen[1549]),

			.SO(gen[1607]),
			.S(gen[1608]),
			.SE(gen[1609]),

			.SELF(gen[1548]),
			.cell_state(gen[1548])
		); 

/******************* CELL 1549 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1549 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1488]),
			.N(gen[1489]),
			.NE(gen[1490]),

			.O(gen[1548]),
			.E(gen[1550]),

			.SO(gen[1608]),
			.S(gen[1609]),
			.SE(gen[1610]),

			.SELF(gen[1549]),
			.cell_state(gen[1549])
		); 

/******************* CELL 1550 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1550 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1489]),
			.N(gen[1490]),
			.NE(gen[1491]),

			.O(gen[1549]),
			.E(gen[1551]),

			.SO(gen[1609]),
			.S(gen[1610]),
			.SE(gen[1611]),

			.SELF(gen[1550]),
			.cell_state(gen[1550])
		); 

/******************* CELL 1551 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1551 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1490]),
			.N(gen[1491]),
			.NE(gen[1492]),

			.O(gen[1550]),
			.E(gen[1552]),

			.SO(gen[1610]),
			.S(gen[1611]),
			.SE(gen[1612]),

			.SELF(gen[1551]),
			.cell_state(gen[1551])
		); 

/******************* CELL 1552 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1552 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1491]),
			.N(gen[1492]),
			.NE(gen[1493]),

			.O(gen[1551]),
			.E(gen[1553]),

			.SO(gen[1611]),
			.S(gen[1612]),
			.SE(gen[1613]),

			.SELF(gen[1552]),
			.cell_state(gen[1552])
		); 

/******************* CELL 1553 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1553 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1492]),
			.N(gen[1493]),
			.NE(gen[1494]),

			.O(gen[1552]),
			.E(gen[1554]),

			.SO(gen[1612]),
			.S(gen[1613]),
			.SE(gen[1614]),

			.SELF(gen[1553]),
			.cell_state(gen[1553])
		); 

/******************* CELL 1554 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1554 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1493]),
			.N(gen[1494]),
			.NE(gen[1495]),

			.O(gen[1553]),
			.E(gen[1555]),

			.SO(gen[1613]),
			.S(gen[1614]),
			.SE(gen[1615]),

			.SELF(gen[1554]),
			.cell_state(gen[1554])
		); 

/******************* CELL 1555 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1555 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1494]),
			.N(gen[1495]),
			.NE(gen[1496]),

			.O(gen[1554]),
			.E(gen[1556]),

			.SO(gen[1614]),
			.S(gen[1615]),
			.SE(gen[1616]),

			.SELF(gen[1555]),
			.cell_state(gen[1555])
		); 

/******************* CELL 1556 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1556 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1495]),
			.N(gen[1496]),
			.NE(gen[1497]),

			.O(gen[1555]),
			.E(gen[1557]),

			.SO(gen[1615]),
			.S(gen[1616]),
			.SE(gen[1617]),

			.SELF(gen[1556]),
			.cell_state(gen[1556])
		); 

/******************* CELL 1557 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1557 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1496]),
			.N(gen[1497]),
			.NE(gen[1498]),

			.O(gen[1556]),
			.E(gen[1558]),

			.SO(gen[1616]),
			.S(gen[1617]),
			.SE(gen[1618]),

			.SELF(gen[1557]),
			.cell_state(gen[1557])
		); 

/******************* CELL 1558 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1558 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1497]),
			.N(gen[1498]),
			.NE(gen[1499]),

			.O(gen[1557]),
			.E(gen[1559]),

			.SO(gen[1617]),
			.S(gen[1618]),
			.SE(gen[1619]),

			.SELF(gen[1558]),
			.cell_state(gen[1558])
		); 

/******************* CELL 1559 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1559 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1498]),
			.N(gen[1499]),
			.NE(gen[1498]),

			.O(gen[1558]),
			.E(gen[1558]),

			.SO(gen[1618]),
			.S(gen[1619]),
			.SE(gen[1618]),

			.SELF(gen[1559]),
			.cell_state(gen[1559])
		); 

/******************* CELL 1560 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1560 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1501]),
			.N(gen[1500]),
			.NE(gen[1501]),

			.O(gen[1561]),
			.E(gen[1561]),

			.SO(gen[1621]),
			.S(gen[1620]),
			.SE(gen[1621]),

			.SELF(gen[1560]),
			.cell_state(gen[1560])
		); 

/******************* CELL 1561 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1561 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1500]),
			.N(gen[1501]),
			.NE(gen[1502]),

			.O(gen[1560]),
			.E(gen[1562]),

			.SO(gen[1620]),
			.S(gen[1621]),
			.SE(gen[1622]),

			.SELF(gen[1561]),
			.cell_state(gen[1561])
		); 

/******************* CELL 1562 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1562 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1501]),
			.N(gen[1502]),
			.NE(gen[1503]),

			.O(gen[1561]),
			.E(gen[1563]),

			.SO(gen[1621]),
			.S(gen[1622]),
			.SE(gen[1623]),

			.SELF(gen[1562]),
			.cell_state(gen[1562])
		); 

/******************* CELL 1563 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1563 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1502]),
			.N(gen[1503]),
			.NE(gen[1504]),

			.O(gen[1562]),
			.E(gen[1564]),

			.SO(gen[1622]),
			.S(gen[1623]),
			.SE(gen[1624]),

			.SELF(gen[1563]),
			.cell_state(gen[1563])
		); 

/******************* CELL 1564 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1564 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1503]),
			.N(gen[1504]),
			.NE(gen[1505]),

			.O(gen[1563]),
			.E(gen[1565]),

			.SO(gen[1623]),
			.S(gen[1624]),
			.SE(gen[1625]),

			.SELF(gen[1564]),
			.cell_state(gen[1564])
		); 

/******************* CELL 1565 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1565 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1504]),
			.N(gen[1505]),
			.NE(gen[1506]),

			.O(gen[1564]),
			.E(gen[1566]),

			.SO(gen[1624]),
			.S(gen[1625]),
			.SE(gen[1626]),

			.SELF(gen[1565]),
			.cell_state(gen[1565])
		); 

/******************* CELL 1566 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1566 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1505]),
			.N(gen[1506]),
			.NE(gen[1507]),

			.O(gen[1565]),
			.E(gen[1567]),

			.SO(gen[1625]),
			.S(gen[1626]),
			.SE(gen[1627]),

			.SELF(gen[1566]),
			.cell_state(gen[1566])
		); 

/******************* CELL 1567 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1567 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1506]),
			.N(gen[1507]),
			.NE(gen[1508]),

			.O(gen[1566]),
			.E(gen[1568]),

			.SO(gen[1626]),
			.S(gen[1627]),
			.SE(gen[1628]),

			.SELF(gen[1567]),
			.cell_state(gen[1567])
		); 

/******************* CELL 1568 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1568 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1507]),
			.N(gen[1508]),
			.NE(gen[1509]),

			.O(gen[1567]),
			.E(gen[1569]),

			.SO(gen[1627]),
			.S(gen[1628]),
			.SE(gen[1629]),

			.SELF(gen[1568]),
			.cell_state(gen[1568])
		); 

/******************* CELL 1569 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1569 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1508]),
			.N(gen[1509]),
			.NE(gen[1510]),

			.O(gen[1568]),
			.E(gen[1570]),

			.SO(gen[1628]),
			.S(gen[1629]),
			.SE(gen[1630]),

			.SELF(gen[1569]),
			.cell_state(gen[1569])
		); 

/******************* CELL 1570 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1570 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1509]),
			.N(gen[1510]),
			.NE(gen[1511]),

			.O(gen[1569]),
			.E(gen[1571]),

			.SO(gen[1629]),
			.S(gen[1630]),
			.SE(gen[1631]),

			.SELF(gen[1570]),
			.cell_state(gen[1570])
		); 

/******************* CELL 1571 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1571 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1510]),
			.N(gen[1511]),
			.NE(gen[1512]),

			.O(gen[1570]),
			.E(gen[1572]),

			.SO(gen[1630]),
			.S(gen[1631]),
			.SE(gen[1632]),

			.SELF(gen[1571]),
			.cell_state(gen[1571])
		); 

/******************* CELL 1572 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1572 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1511]),
			.N(gen[1512]),
			.NE(gen[1513]),

			.O(gen[1571]),
			.E(gen[1573]),

			.SO(gen[1631]),
			.S(gen[1632]),
			.SE(gen[1633]),

			.SELF(gen[1572]),
			.cell_state(gen[1572])
		); 

/******************* CELL 1573 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1573 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1512]),
			.N(gen[1513]),
			.NE(gen[1514]),

			.O(gen[1572]),
			.E(gen[1574]),

			.SO(gen[1632]),
			.S(gen[1633]),
			.SE(gen[1634]),

			.SELF(gen[1573]),
			.cell_state(gen[1573])
		); 

/******************* CELL 1574 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1574 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1513]),
			.N(gen[1514]),
			.NE(gen[1515]),

			.O(gen[1573]),
			.E(gen[1575]),

			.SO(gen[1633]),
			.S(gen[1634]),
			.SE(gen[1635]),

			.SELF(gen[1574]),
			.cell_state(gen[1574])
		); 

/******************* CELL 1575 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1575 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1514]),
			.N(gen[1515]),
			.NE(gen[1516]),

			.O(gen[1574]),
			.E(gen[1576]),

			.SO(gen[1634]),
			.S(gen[1635]),
			.SE(gen[1636]),

			.SELF(gen[1575]),
			.cell_state(gen[1575])
		); 

/******************* CELL 1576 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1576 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1515]),
			.N(gen[1516]),
			.NE(gen[1517]),

			.O(gen[1575]),
			.E(gen[1577]),

			.SO(gen[1635]),
			.S(gen[1636]),
			.SE(gen[1637]),

			.SELF(gen[1576]),
			.cell_state(gen[1576])
		); 

/******************* CELL 1577 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1577 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1516]),
			.N(gen[1517]),
			.NE(gen[1518]),

			.O(gen[1576]),
			.E(gen[1578]),

			.SO(gen[1636]),
			.S(gen[1637]),
			.SE(gen[1638]),

			.SELF(gen[1577]),
			.cell_state(gen[1577])
		); 

/******************* CELL 1578 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1578 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1517]),
			.N(gen[1518]),
			.NE(gen[1519]),

			.O(gen[1577]),
			.E(gen[1579]),

			.SO(gen[1637]),
			.S(gen[1638]),
			.SE(gen[1639]),

			.SELF(gen[1578]),
			.cell_state(gen[1578])
		); 

/******************* CELL 1579 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1579 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1518]),
			.N(gen[1519]),
			.NE(gen[1520]),

			.O(gen[1578]),
			.E(gen[1580]),

			.SO(gen[1638]),
			.S(gen[1639]),
			.SE(gen[1640]),

			.SELF(gen[1579]),
			.cell_state(gen[1579])
		); 

/******************* CELL 1580 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1580 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1519]),
			.N(gen[1520]),
			.NE(gen[1521]),

			.O(gen[1579]),
			.E(gen[1581]),

			.SO(gen[1639]),
			.S(gen[1640]),
			.SE(gen[1641]),

			.SELF(gen[1580]),
			.cell_state(gen[1580])
		); 

/******************* CELL 1581 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1581 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1520]),
			.N(gen[1521]),
			.NE(gen[1522]),

			.O(gen[1580]),
			.E(gen[1582]),

			.SO(gen[1640]),
			.S(gen[1641]),
			.SE(gen[1642]),

			.SELF(gen[1581]),
			.cell_state(gen[1581])
		); 

/******************* CELL 1582 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1582 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1521]),
			.N(gen[1522]),
			.NE(gen[1523]),

			.O(gen[1581]),
			.E(gen[1583]),

			.SO(gen[1641]),
			.S(gen[1642]),
			.SE(gen[1643]),

			.SELF(gen[1582]),
			.cell_state(gen[1582])
		); 

/******************* CELL 1583 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1583 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1522]),
			.N(gen[1523]),
			.NE(gen[1524]),

			.O(gen[1582]),
			.E(gen[1584]),

			.SO(gen[1642]),
			.S(gen[1643]),
			.SE(gen[1644]),

			.SELF(gen[1583]),
			.cell_state(gen[1583])
		); 

/******************* CELL 1584 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1584 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1523]),
			.N(gen[1524]),
			.NE(gen[1525]),

			.O(gen[1583]),
			.E(gen[1585]),

			.SO(gen[1643]),
			.S(gen[1644]),
			.SE(gen[1645]),

			.SELF(gen[1584]),
			.cell_state(gen[1584])
		); 

/******************* CELL 1585 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1585 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1524]),
			.N(gen[1525]),
			.NE(gen[1526]),

			.O(gen[1584]),
			.E(gen[1586]),

			.SO(gen[1644]),
			.S(gen[1645]),
			.SE(gen[1646]),

			.SELF(gen[1585]),
			.cell_state(gen[1585])
		); 

/******************* CELL 1586 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1586 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1525]),
			.N(gen[1526]),
			.NE(gen[1527]),

			.O(gen[1585]),
			.E(gen[1587]),

			.SO(gen[1645]),
			.S(gen[1646]),
			.SE(gen[1647]),

			.SELF(gen[1586]),
			.cell_state(gen[1586])
		); 

/******************* CELL 1587 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1587 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1526]),
			.N(gen[1527]),
			.NE(gen[1528]),

			.O(gen[1586]),
			.E(gen[1588]),

			.SO(gen[1646]),
			.S(gen[1647]),
			.SE(gen[1648]),

			.SELF(gen[1587]),
			.cell_state(gen[1587])
		); 

/******************* CELL 1588 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1588 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1527]),
			.N(gen[1528]),
			.NE(gen[1529]),

			.O(gen[1587]),
			.E(gen[1589]),

			.SO(gen[1647]),
			.S(gen[1648]),
			.SE(gen[1649]),

			.SELF(gen[1588]),
			.cell_state(gen[1588])
		); 

/******************* CELL 1589 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1589 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1528]),
			.N(gen[1529]),
			.NE(gen[1530]),

			.O(gen[1588]),
			.E(gen[1590]),

			.SO(gen[1648]),
			.S(gen[1649]),
			.SE(gen[1650]),

			.SELF(gen[1589]),
			.cell_state(gen[1589])
		); 

/******************* CELL 1590 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1590 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1529]),
			.N(gen[1530]),
			.NE(gen[1531]),

			.O(gen[1589]),
			.E(gen[1591]),

			.SO(gen[1649]),
			.S(gen[1650]),
			.SE(gen[1651]),

			.SELF(gen[1590]),
			.cell_state(gen[1590])
		); 

/******************* CELL 1591 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1591 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1530]),
			.N(gen[1531]),
			.NE(gen[1532]),

			.O(gen[1590]),
			.E(gen[1592]),

			.SO(gen[1650]),
			.S(gen[1651]),
			.SE(gen[1652]),

			.SELF(gen[1591]),
			.cell_state(gen[1591])
		); 

/******************* CELL 1592 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1592 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1531]),
			.N(gen[1532]),
			.NE(gen[1533]),

			.O(gen[1591]),
			.E(gen[1593]),

			.SO(gen[1651]),
			.S(gen[1652]),
			.SE(gen[1653]),

			.SELF(gen[1592]),
			.cell_state(gen[1592])
		); 

/******************* CELL 1593 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1593 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1532]),
			.N(gen[1533]),
			.NE(gen[1534]),

			.O(gen[1592]),
			.E(gen[1594]),

			.SO(gen[1652]),
			.S(gen[1653]),
			.SE(gen[1654]),

			.SELF(gen[1593]),
			.cell_state(gen[1593])
		); 

/******************* CELL 1594 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1594 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1533]),
			.N(gen[1534]),
			.NE(gen[1535]),

			.O(gen[1593]),
			.E(gen[1595]),

			.SO(gen[1653]),
			.S(gen[1654]),
			.SE(gen[1655]),

			.SELF(gen[1594]),
			.cell_state(gen[1594])
		); 

/******************* CELL 1595 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1595 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1534]),
			.N(gen[1535]),
			.NE(gen[1536]),

			.O(gen[1594]),
			.E(gen[1596]),

			.SO(gen[1654]),
			.S(gen[1655]),
			.SE(gen[1656]),

			.SELF(gen[1595]),
			.cell_state(gen[1595])
		); 

/******************* CELL 1596 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1596 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1535]),
			.N(gen[1536]),
			.NE(gen[1537]),

			.O(gen[1595]),
			.E(gen[1597]),

			.SO(gen[1655]),
			.S(gen[1656]),
			.SE(gen[1657]),

			.SELF(gen[1596]),
			.cell_state(gen[1596])
		); 

/******************* CELL 1597 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1597 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1536]),
			.N(gen[1537]),
			.NE(gen[1538]),

			.O(gen[1596]),
			.E(gen[1598]),

			.SO(gen[1656]),
			.S(gen[1657]),
			.SE(gen[1658]),

			.SELF(gen[1597]),
			.cell_state(gen[1597])
		); 

/******************* CELL 1598 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1598 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1537]),
			.N(gen[1538]),
			.NE(gen[1539]),

			.O(gen[1597]),
			.E(gen[1599]),

			.SO(gen[1657]),
			.S(gen[1658]),
			.SE(gen[1659]),

			.SELF(gen[1598]),
			.cell_state(gen[1598])
		); 

/******************* CELL 1599 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1599 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1538]),
			.N(gen[1539]),
			.NE(gen[1540]),

			.O(gen[1598]),
			.E(gen[1600]),

			.SO(gen[1658]),
			.S(gen[1659]),
			.SE(gen[1660]),

			.SELF(gen[1599]),
			.cell_state(gen[1599])
		); 

/******************* CELL 1600 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1600 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1539]),
			.N(gen[1540]),
			.NE(gen[1541]),

			.O(gen[1599]),
			.E(gen[1601]),

			.SO(gen[1659]),
			.S(gen[1660]),
			.SE(gen[1661]),

			.SELF(gen[1600]),
			.cell_state(gen[1600])
		); 

/******************* CELL 1601 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1601 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1540]),
			.N(gen[1541]),
			.NE(gen[1542]),

			.O(gen[1600]),
			.E(gen[1602]),

			.SO(gen[1660]),
			.S(gen[1661]),
			.SE(gen[1662]),

			.SELF(gen[1601]),
			.cell_state(gen[1601])
		); 

/******************* CELL 1602 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1602 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1541]),
			.N(gen[1542]),
			.NE(gen[1543]),

			.O(gen[1601]),
			.E(gen[1603]),

			.SO(gen[1661]),
			.S(gen[1662]),
			.SE(gen[1663]),

			.SELF(gen[1602]),
			.cell_state(gen[1602])
		); 

/******************* CELL 1603 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1603 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1542]),
			.N(gen[1543]),
			.NE(gen[1544]),

			.O(gen[1602]),
			.E(gen[1604]),

			.SO(gen[1662]),
			.S(gen[1663]),
			.SE(gen[1664]),

			.SELF(gen[1603]),
			.cell_state(gen[1603])
		); 

/******************* CELL 1604 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1604 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1543]),
			.N(gen[1544]),
			.NE(gen[1545]),

			.O(gen[1603]),
			.E(gen[1605]),

			.SO(gen[1663]),
			.S(gen[1664]),
			.SE(gen[1665]),

			.SELF(gen[1604]),
			.cell_state(gen[1604])
		); 

/******************* CELL 1605 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1605 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1544]),
			.N(gen[1545]),
			.NE(gen[1546]),

			.O(gen[1604]),
			.E(gen[1606]),

			.SO(gen[1664]),
			.S(gen[1665]),
			.SE(gen[1666]),

			.SELF(gen[1605]),
			.cell_state(gen[1605])
		); 

/******************* CELL 1606 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1606 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1545]),
			.N(gen[1546]),
			.NE(gen[1547]),

			.O(gen[1605]),
			.E(gen[1607]),

			.SO(gen[1665]),
			.S(gen[1666]),
			.SE(gen[1667]),

			.SELF(gen[1606]),
			.cell_state(gen[1606])
		); 

/******************* CELL 1607 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1607 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1546]),
			.N(gen[1547]),
			.NE(gen[1548]),

			.O(gen[1606]),
			.E(gen[1608]),

			.SO(gen[1666]),
			.S(gen[1667]),
			.SE(gen[1668]),

			.SELF(gen[1607]),
			.cell_state(gen[1607])
		); 

/******************* CELL 1608 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1608 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1547]),
			.N(gen[1548]),
			.NE(gen[1549]),

			.O(gen[1607]),
			.E(gen[1609]),

			.SO(gen[1667]),
			.S(gen[1668]),
			.SE(gen[1669]),

			.SELF(gen[1608]),
			.cell_state(gen[1608])
		); 

/******************* CELL 1609 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1609 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1548]),
			.N(gen[1549]),
			.NE(gen[1550]),

			.O(gen[1608]),
			.E(gen[1610]),

			.SO(gen[1668]),
			.S(gen[1669]),
			.SE(gen[1670]),

			.SELF(gen[1609]),
			.cell_state(gen[1609])
		); 

/******************* CELL 1610 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1610 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1549]),
			.N(gen[1550]),
			.NE(gen[1551]),

			.O(gen[1609]),
			.E(gen[1611]),

			.SO(gen[1669]),
			.S(gen[1670]),
			.SE(gen[1671]),

			.SELF(gen[1610]),
			.cell_state(gen[1610])
		); 

/******************* CELL 1611 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1611 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1550]),
			.N(gen[1551]),
			.NE(gen[1552]),

			.O(gen[1610]),
			.E(gen[1612]),

			.SO(gen[1670]),
			.S(gen[1671]),
			.SE(gen[1672]),

			.SELF(gen[1611]),
			.cell_state(gen[1611])
		); 

/******************* CELL 1612 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1612 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1551]),
			.N(gen[1552]),
			.NE(gen[1553]),

			.O(gen[1611]),
			.E(gen[1613]),

			.SO(gen[1671]),
			.S(gen[1672]),
			.SE(gen[1673]),

			.SELF(gen[1612]),
			.cell_state(gen[1612])
		); 

/******************* CELL 1613 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1613 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1552]),
			.N(gen[1553]),
			.NE(gen[1554]),

			.O(gen[1612]),
			.E(gen[1614]),

			.SO(gen[1672]),
			.S(gen[1673]),
			.SE(gen[1674]),

			.SELF(gen[1613]),
			.cell_state(gen[1613])
		); 

/******************* CELL 1614 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1614 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1553]),
			.N(gen[1554]),
			.NE(gen[1555]),

			.O(gen[1613]),
			.E(gen[1615]),

			.SO(gen[1673]),
			.S(gen[1674]),
			.SE(gen[1675]),

			.SELF(gen[1614]),
			.cell_state(gen[1614])
		); 

/******************* CELL 1615 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1615 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1554]),
			.N(gen[1555]),
			.NE(gen[1556]),

			.O(gen[1614]),
			.E(gen[1616]),

			.SO(gen[1674]),
			.S(gen[1675]),
			.SE(gen[1676]),

			.SELF(gen[1615]),
			.cell_state(gen[1615])
		); 

/******************* CELL 1616 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1616 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1555]),
			.N(gen[1556]),
			.NE(gen[1557]),

			.O(gen[1615]),
			.E(gen[1617]),

			.SO(gen[1675]),
			.S(gen[1676]),
			.SE(gen[1677]),

			.SELF(gen[1616]),
			.cell_state(gen[1616])
		); 

/******************* CELL 1617 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1617 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1556]),
			.N(gen[1557]),
			.NE(gen[1558]),

			.O(gen[1616]),
			.E(gen[1618]),

			.SO(gen[1676]),
			.S(gen[1677]),
			.SE(gen[1678]),

			.SELF(gen[1617]),
			.cell_state(gen[1617])
		); 

/******************* CELL 1618 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1618 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1557]),
			.N(gen[1558]),
			.NE(gen[1559]),

			.O(gen[1617]),
			.E(gen[1619]),

			.SO(gen[1677]),
			.S(gen[1678]),
			.SE(gen[1679]),

			.SELF(gen[1618]),
			.cell_state(gen[1618])
		); 

/******************* CELL 1619 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1619 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1558]),
			.N(gen[1559]),
			.NE(gen[1558]),

			.O(gen[1618]),
			.E(gen[1618]),

			.SO(gen[1678]),
			.S(gen[1679]),
			.SE(gen[1678]),

			.SELF(gen[1619]),
			.cell_state(gen[1619])
		); 

/******************* CELL 1620 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1620 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1561]),
			.N(gen[1560]),
			.NE(gen[1561]),

			.O(gen[1621]),
			.E(gen[1621]),

			.SO(gen[1681]),
			.S(gen[1680]),
			.SE(gen[1681]),

			.SELF(gen[1620]),
			.cell_state(gen[1620])
		); 

/******************* CELL 1621 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1621 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1560]),
			.N(gen[1561]),
			.NE(gen[1562]),

			.O(gen[1620]),
			.E(gen[1622]),

			.SO(gen[1680]),
			.S(gen[1681]),
			.SE(gen[1682]),

			.SELF(gen[1621]),
			.cell_state(gen[1621])
		); 

/******************* CELL 1622 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1622 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1561]),
			.N(gen[1562]),
			.NE(gen[1563]),

			.O(gen[1621]),
			.E(gen[1623]),

			.SO(gen[1681]),
			.S(gen[1682]),
			.SE(gen[1683]),

			.SELF(gen[1622]),
			.cell_state(gen[1622])
		); 

/******************* CELL 1623 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1623 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1562]),
			.N(gen[1563]),
			.NE(gen[1564]),

			.O(gen[1622]),
			.E(gen[1624]),

			.SO(gen[1682]),
			.S(gen[1683]),
			.SE(gen[1684]),

			.SELF(gen[1623]),
			.cell_state(gen[1623])
		); 

/******************* CELL 1624 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1624 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1563]),
			.N(gen[1564]),
			.NE(gen[1565]),

			.O(gen[1623]),
			.E(gen[1625]),

			.SO(gen[1683]),
			.S(gen[1684]),
			.SE(gen[1685]),

			.SELF(gen[1624]),
			.cell_state(gen[1624])
		); 

/******************* CELL 1625 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1625 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1564]),
			.N(gen[1565]),
			.NE(gen[1566]),

			.O(gen[1624]),
			.E(gen[1626]),

			.SO(gen[1684]),
			.S(gen[1685]),
			.SE(gen[1686]),

			.SELF(gen[1625]),
			.cell_state(gen[1625])
		); 

/******************* CELL 1626 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1626 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1565]),
			.N(gen[1566]),
			.NE(gen[1567]),

			.O(gen[1625]),
			.E(gen[1627]),

			.SO(gen[1685]),
			.S(gen[1686]),
			.SE(gen[1687]),

			.SELF(gen[1626]),
			.cell_state(gen[1626])
		); 

/******************* CELL 1627 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1627 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1566]),
			.N(gen[1567]),
			.NE(gen[1568]),

			.O(gen[1626]),
			.E(gen[1628]),

			.SO(gen[1686]),
			.S(gen[1687]),
			.SE(gen[1688]),

			.SELF(gen[1627]),
			.cell_state(gen[1627])
		); 

/******************* CELL 1628 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1628 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1567]),
			.N(gen[1568]),
			.NE(gen[1569]),

			.O(gen[1627]),
			.E(gen[1629]),

			.SO(gen[1687]),
			.S(gen[1688]),
			.SE(gen[1689]),

			.SELF(gen[1628]),
			.cell_state(gen[1628])
		); 

/******************* CELL 1629 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1629 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1568]),
			.N(gen[1569]),
			.NE(gen[1570]),

			.O(gen[1628]),
			.E(gen[1630]),

			.SO(gen[1688]),
			.S(gen[1689]),
			.SE(gen[1690]),

			.SELF(gen[1629]),
			.cell_state(gen[1629])
		); 

/******************* CELL 1630 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1630 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1569]),
			.N(gen[1570]),
			.NE(gen[1571]),

			.O(gen[1629]),
			.E(gen[1631]),

			.SO(gen[1689]),
			.S(gen[1690]),
			.SE(gen[1691]),

			.SELF(gen[1630]),
			.cell_state(gen[1630])
		); 

/******************* CELL 1631 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1631 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1570]),
			.N(gen[1571]),
			.NE(gen[1572]),

			.O(gen[1630]),
			.E(gen[1632]),

			.SO(gen[1690]),
			.S(gen[1691]),
			.SE(gen[1692]),

			.SELF(gen[1631]),
			.cell_state(gen[1631])
		); 

/******************* CELL 1632 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1632 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1571]),
			.N(gen[1572]),
			.NE(gen[1573]),

			.O(gen[1631]),
			.E(gen[1633]),

			.SO(gen[1691]),
			.S(gen[1692]),
			.SE(gen[1693]),

			.SELF(gen[1632]),
			.cell_state(gen[1632])
		); 

/******************* CELL 1633 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1633 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1572]),
			.N(gen[1573]),
			.NE(gen[1574]),

			.O(gen[1632]),
			.E(gen[1634]),

			.SO(gen[1692]),
			.S(gen[1693]),
			.SE(gen[1694]),

			.SELF(gen[1633]),
			.cell_state(gen[1633])
		); 

/******************* CELL 1634 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1634 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1573]),
			.N(gen[1574]),
			.NE(gen[1575]),

			.O(gen[1633]),
			.E(gen[1635]),

			.SO(gen[1693]),
			.S(gen[1694]),
			.SE(gen[1695]),

			.SELF(gen[1634]),
			.cell_state(gen[1634])
		); 

/******************* CELL 1635 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1635 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1574]),
			.N(gen[1575]),
			.NE(gen[1576]),

			.O(gen[1634]),
			.E(gen[1636]),

			.SO(gen[1694]),
			.S(gen[1695]),
			.SE(gen[1696]),

			.SELF(gen[1635]),
			.cell_state(gen[1635])
		); 

/******************* CELL 1636 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1636 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1575]),
			.N(gen[1576]),
			.NE(gen[1577]),

			.O(gen[1635]),
			.E(gen[1637]),

			.SO(gen[1695]),
			.S(gen[1696]),
			.SE(gen[1697]),

			.SELF(gen[1636]),
			.cell_state(gen[1636])
		); 

/******************* CELL 1637 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1637 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1576]),
			.N(gen[1577]),
			.NE(gen[1578]),

			.O(gen[1636]),
			.E(gen[1638]),

			.SO(gen[1696]),
			.S(gen[1697]),
			.SE(gen[1698]),

			.SELF(gen[1637]),
			.cell_state(gen[1637])
		); 

/******************* CELL 1638 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1638 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1577]),
			.N(gen[1578]),
			.NE(gen[1579]),

			.O(gen[1637]),
			.E(gen[1639]),

			.SO(gen[1697]),
			.S(gen[1698]),
			.SE(gen[1699]),

			.SELF(gen[1638]),
			.cell_state(gen[1638])
		); 

/******************* CELL 1639 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1639 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1578]),
			.N(gen[1579]),
			.NE(gen[1580]),

			.O(gen[1638]),
			.E(gen[1640]),

			.SO(gen[1698]),
			.S(gen[1699]),
			.SE(gen[1700]),

			.SELF(gen[1639]),
			.cell_state(gen[1639])
		); 

/******************* CELL 1640 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1640 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1579]),
			.N(gen[1580]),
			.NE(gen[1581]),

			.O(gen[1639]),
			.E(gen[1641]),

			.SO(gen[1699]),
			.S(gen[1700]),
			.SE(gen[1701]),

			.SELF(gen[1640]),
			.cell_state(gen[1640])
		); 

/******************* CELL 1641 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1641 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1580]),
			.N(gen[1581]),
			.NE(gen[1582]),

			.O(gen[1640]),
			.E(gen[1642]),

			.SO(gen[1700]),
			.S(gen[1701]),
			.SE(gen[1702]),

			.SELF(gen[1641]),
			.cell_state(gen[1641])
		); 

/******************* CELL 1642 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1642 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1581]),
			.N(gen[1582]),
			.NE(gen[1583]),

			.O(gen[1641]),
			.E(gen[1643]),

			.SO(gen[1701]),
			.S(gen[1702]),
			.SE(gen[1703]),

			.SELF(gen[1642]),
			.cell_state(gen[1642])
		); 

/******************* CELL 1643 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1643 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1582]),
			.N(gen[1583]),
			.NE(gen[1584]),

			.O(gen[1642]),
			.E(gen[1644]),

			.SO(gen[1702]),
			.S(gen[1703]),
			.SE(gen[1704]),

			.SELF(gen[1643]),
			.cell_state(gen[1643])
		); 

/******************* CELL 1644 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1644 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1583]),
			.N(gen[1584]),
			.NE(gen[1585]),

			.O(gen[1643]),
			.E(gen[1645]),

			.SO(gen[1703]),
			.S(gen[1704]),
			.SE(gen[1705]),

			.SELF(gen[1644]),
			.cell_state(gen[1644])
		); 

/******************* CELL 1645 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1645 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1584]),
			.N(gen[1585]),
			.NE(gen[1586]),

			.O(gen[1644]),
			.E(gen[1646]),

			.SO(gen[1704]),
			.S(gen[1705]),
			.SE(gen[1706]),

			.SELF(gen[1645]),
			.cell_state(gen[1645])
		); 

/******************* CELL 1646 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1646 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1585]),
			.N(gen[1586]),
			.NE(gen[1587]),

			.O(gen[1645]),
			.E(gen[1647]),

			.SO(gen[1705]),
			.S(gen[1706]),
			.SE(gen[1707]),

			.SELF(gen[1646]),
			.cell_state(gen[1646])
		); 

/******************* CELL 1647 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1647 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1586]),
			.N(gen[1587]),
			.NE(gen[1588]),

			.O(gen[1646]),
			.E(gen[1648]),

			.SO(gen[1706]),
			.S(gen[1707]),
			.SE(gen[1708]),

			.SELF(gen[1647]),
			.cell_state(gen[1647])
		); 

/******************* CELL 1648 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1648 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1587]),
			.N(gen[1588]),
			.NE(gen[1589]),

			.O(gen[1647]),
			.E(gen[1649]),

			.SO(gen[1707]),
			.S(gen[1708]),
			.SE(gen[1709]),

			.SELF(gen[1648]),
			.cell_state(gen[1648])
		); 

/******************* CELL 1649 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1649 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1588]),
			.N(gen[1589]),
			.NE(gen[1590]),

			.O(gen[1648]),
			.E(gen[1650]),

			.SO(gen[1708]),
			.S(gen[1709]),
			.SE(gen[1710]),

			.SELF(gen[1649]),
			.cell_state(gen[1649])
		); 

/******************* CELL 1650 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1650 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1589]),
			.N(gen[1590]),
			.NE(gen[1591]),

			.O(gen[1649]),
			.E(gen[1651]),

			.SO(gen[1709]),
			.S(gen[1710]),
			.SE(gen[1711]),

			.SELF(gen[1650]),
			.cell_state(gen[1650])
		); 

/******************* CELL 1651 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1651 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1590]),
			.N(gen[1591]),
			.NE(gen[1592]),

			.O(gen[1650]),
			.E(gen[1652]),

			.SO(gen[1710]),
			.S(gen[1711]),
			.SE(gen[1712]),

			.SELF(gen[1651]),
			.cell_state(gen[1651])
		); 

/******************* CELL 1652 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1652 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1591]),
			.N(gen[1592]),
			.NE(gen[1593]),

			.O(gen[1651]),
			.E(gen[1653]),

			.SO(gen[1711]),
			.S(gen[1712]),
			.SE(gen[1713]),

			.SELF(gen[1652]),
			.cell_state(gen[1652])
		); 

/******************* CELL 1653 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1653 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1592]),
			.N(gen[1593]),
			.NE(gen[1594]),

			.O(gen[1652]),
			.E(gen[1654]),

			.SO(gen[1712]),
			.S(gen[1713]),
			.SE(gen[1714]),

			.SELF(gen[1653]),
			.cell_state(gen[1653])
		); 

/******************* CELL 1654 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1654 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1593]),
			.N(gen[1594]),
			.NE(gen[1595]),

			.O(gen[1653]),
			.E(gen[1655]),

			.SO(gen[1713]),
			.S(gen[1714]),
			.SE(gen[1715]),

			.SELF(gen[1654]),
			.cell_state(gen[1654])
		); 

/******************* CELL 1655 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1655 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1594]),
			.N(gen[1595]),
			.NE(gen[1596]),

			.O(gen[1654]),
			.E(gen[1656]),

			.SO(gen[1714]),
			.S(gen[1715]),
			.SE(gen[1716]),

			.SELF(gen[1655]),
			.cell_state(gen[1655])
		); 

/******************* CELL 1656 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1656 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1595]),
			.N(gen[1596]),
			.NE(gen[1597]),

			.O(gen[1655]),
			.E(gen[1657]),

			.SO(gen[1715]),
			.S(gen[1716]),
			.SE(gen[1717]),

			.SELF(gen[1656]),
			.cell_state(gen[1656])
		); 

/******************* CELL 1657 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1657 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1596]),
			.N(gen[1597]),
			.NE(gen[1598]),

			.O(gen[1656]),
			.E(gen[1658]),

			.SO(gen[1716]),
			.S(gen[1717]),
			.SE(gen[1718]),

			.SELF(gen[1657]),
			.cell_state(gen[1657])
		); 

/******************* CELL 1658 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1658 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1597]),
			.N(gen[1598]),
			.NE(gen[1599]),

			.O(gen[1657]),
			.E(gen[1659]),

			.SO(gen[1717]),
			.S(gen[1718]),
			.SE(gen[1719]),

			.SELF(gen[1658]),
			.cell_state(gen[1658])
		); 

/******************* CELL 1659 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1659 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1598]),
			.N(gen[1599]),
			.NE(gen[1600]),

			.O(gen[1658]),
			.E(gen[1660]),

			.SO(gen[1718]),
			.S(gen[1719]),
			.SE(gen[1720]),

			.SELF(gen[1659]),
			.cell_state(gen[1659])
		); 

/******************* CELL 1660 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1660 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1599]),
			.N(gen[1600]),
			.NE(gen[1601]),

			.O(gen[1659]),
			.E(gen[1661]),

			.SO(gen[1719]),
			.S(gen[1720]),
			.SE(gen[1721]),

			.SELF(gen[1660]),
			.cell_state(gen[1660])
		); 

/******************* CELL 1661 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1661 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1600]),
			.N(gen[1601]),
			.NE(gen[1602]),

			.O(gen[1660]),
			.E(gen[1662]),

			.SO(gen[1720]),
			.S(gen[1721]),
			.SE(gen[1722]),

			.SELF(gen[1661]),
			.cell_state(gen[1661])
		); 

/******************* CELL 1662 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1662 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1601]),
			.N(gen[1602]),
			.NE(gen[1603]),

			.O(gen[1661]),
			.E(gen[1663]),

			.SO(gen[1721]),
			.S(gen[1722]),
			.SE(gen[1723]),

			.SELF(gen[1662]),
			.cell_state(gen[1662])
		); 

/******************* CELL 1663 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1663 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1602]),
			.N(gen[1603]),
			.NE(gen[1604]),

			.O(gen[1662]),
			.E(gen[1664]),

			.SO(gen[1722]),
			.S(gen[1723]),
			.SE(gen[1724]),

			.SELF(gen[1663]),
			.cell_state(gen[1663])
		); 

/******************* CELL 1664 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1664 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1603]),
			.N(gen[1604]),
			.NE(gen[1605]),

			.O(gen[1663]),
			.E(gen[1665]),

			.SO(gen[1723]),
			.S(gen[1724]),
			.SE(gen[1725]),

			.SELF(gen[1664]),
			.cell_state(gen[1664])
		); 

/******************* CELL 1665 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1665 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1604]),
			.N(gen[1605]),
			.NE(gen[1606]),

			.O(gen[1664]),
			.E(gen[1666]),

			.SO(gen[1724]),
			.S(gen[1725]),
			.SE(gen[1726]),

			.SELF(gen[1665]),
			.cell_state(gen[1665])
		); 

/******************* CELL 1666 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1666 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1605]),
			.N(gen[1606]),
			.NE(gen[1607]),

			.O(gen[1665]),
			.E(gen[1667]),

			.SO(gen[1725]),
			.S(gen[1726]),
			.SE(gen[1727]),

			.SELF(gen[1666]),
			.cell_state(gen[1666])
		); 

/******************* CELL 1667 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1667 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1606]),
			.N(gen[1607]),
			.NE(gen[1608]),

			.O(gen[1666]),
			.E(gen[1668]),

			.SO(gen[1726]),
			.S(gen[1727]),
			.SE(gen[1728]),

			.SELF(gen[1667]),
			.cell_state(gen[1667])
		); 

/******************* CELL 1668 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1668 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1607]),
			.N(gen[1608]),
			.NE(gen[1609]),

			.O(gen[1667]),
			.E(gen[1669]),

			.SO(gen[1727]),
			.S(gen[1728]),
			.SE(gen[1729]),

			.SELF(gen[1668]),
			.cell_state(gen[1668])
		); 

/******************* CELL 1669 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1669 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1608]),
			.N(gen[1609]),
			.NE(gen[1610]),

			.O(gen[1668]),
			.E(gen[1670]),

			.SO(gen[1728]),
			.S(gen[1729]),
			.SE(gen[1730]),

			.SELF(gen[1669]),
			.cell_state(gen[1669])
		); 

/******************* CELL 1670 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1670 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1609]),
			.N(gen[1610]),
			.NE(gen[1611]),

			.O(gen[1669]),
			.E(gen[1671]),

			.SO(gen[1729]),
			.S(gen[1730]),
			.SE(gen[1731]),

			.SELF(gen[1670]),
			.cell_state(gen[1670])
		); 

/******************* CELL 1671 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1671 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1610]),
			.N(gen[1611]),
			.NE(gen[1612]),

			.O(gen[1670]),
			.E(gen[1672]),

			.SO(gen[1730]),
			.S(gen[1731]),
			.SE(gen[1732]),

			.SELF(gen[1671]),
			.cell_state(gen[1671])
		); 

/******************* CELL 1672 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1672 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1611]),
			.N(gen[1612]),
			.NE(gen[1613]),

			.O(gen[1671]),
			.E(gen[1673]),

			.SO(gen[1731]),
			.S(gen[1732]),
			.SE(gen[1733]),

			.SELF(gen[1672]),
			.cell_state(gen[1672])
		); 

/******************* CELL 1673 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1673 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1612]),
			.N(gen[1613]),
			.NE(gen[1614]),

			.O(gen[1672]),
			.E(gen[1674]),

			.SO(gen[1732]),
			.S(gen[1733]),
			.SE(gen[1734]),

			.SELF(gen[1673]),
			.cell_state(gen[1673])
		); 

/******************* CELL 1674 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1674 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1613]),
			.N(gen[1614]),
			.NE(gen[1615]),

			.O(gen[1673]),
			.E(gen[1675]),

			.SO(gen[1733]),
			.S(gen[1734]),
			.SE(gen[1735]),

			.SELF(gen[1674]),
			.cell_state(gen[1674])
		); 

/******************* CELL 1675 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1675 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1614]),
			.N(gen[1615]),
			.NE(gen[1616]),

			.O(gen[1674]),
			.E(gen[1676]),

			.SO(gen[1734]),
			.S(gen[1735]),
			.SE(gen[1736]),

			.SELF(gen[1675]),
			.cell_state(gen[1675])
		); 

/******************* CELL 1676 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1676 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1615]),
			.N(gen[1616]),
			.NE(gen[1617]),

			.O(gen[1675]),
			.E(gen[1677]),

			.SO(gen[1735]),
			.S(gen[1736]),
			.SE(gen[1737]),

			.SELF(gen[1676]),
			.cell_state(gen[1676])
		); 

/******************* CELL 1677 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1677 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1616]),
			.N(gen[1617]),
			.NE(gen[1618]),

			.O(gen[1676]),
			.E(gen[1678]),

			.SO(gen[1736]),
			.S(gen[1737]),
			.SE(gen[1738]),

			.SELF(gen[1677]),
			.cell_state(gen[1677])
		); 

/******************* CELL 1678 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1678 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1617]),
			.N(gen[1618]),
			.NE(gen[1619]),

			.O(gen[1677]),
			.E(gen[1679]),

			.SO(gen[1737]),
			.S(gen[1738]),
			.SE(gen[1739]),

			.SELF(gen[1678]),
			.cell_state(gen[1678])
		); 

/******************* CELL 1679 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1679 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1618]),
			.N(gen[1619]),
			.NE(gen[1618]),

			.O(gen[1678]),
			.E(gen[1678]),

			.SO(gen[1738]),
			.S(gen[1739]),
			.SE(gen[1738]),

			.SELF(gen[1679]),
			.cell_state(gen[1679])
		); 

/******************* CELL 1680 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1680 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1621]),
			.N(gen[1620]),
			.NE(gen[1621]),

			.O(gen[1681]),
			.E(gen[1681]),

			.SO(gen[1741]),
			.S(gen[1740]),
			.SE(gen[1741]),

			.SELF(gen[1680]),
			.cell_state(gen[1680])
		); 

/******************* CELL 1681 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1681 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1620]),
			.N(gen[1621]),
			.NE(gen[1622]),

			.O(gen[1680]),
			.E(gen[1682]),

			.SO(gen[1740]),
			.S(gen[1741]),
			.SE(gen[1742]),

			.SELF(gen[1681]),
			.cell_state(gen[1681])
		); 

/******************* CELL 1682 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1682 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1621]),
			.N(gen[1622]),
			.NE(gen[1623]),

			.O(gen[1681]),
			.E(gen[1683]),

			.SO(gen[1741]),
			.S(gen[1742]),
			.SE(gen[1743]),

			.SELF(gen[1682]),
			.cell_state(gen[1682])
		); 

/******************* CELL 1683 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1683 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1622]),
			.N(gen[1623]),
			.NE(gen[1624]),

			.O(gen[1682]),
			.E(gen[1684]),

			.SO(gen[1742]),
			.S(gen[1743]),
			.SE(gen[1744]),

			.SELF(gen[1683]),
			.cell_state(gen[1683])
		); 

/******************* CELL 1684 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1684 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1623]),
			.N(gen[1624]),
			.NE(gen[1625]),

			.O(gen[1683]),
			.E(gen[1685]),

			.SO(gen[1743]),
			.S(gen[1744]),
			.SE(gen[1745]),

			.SELF(gen[1684]),
			.cell_state(gen[1684])
		); 

/******************* CELL 1685 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1685 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1624]),
			.N(gen[1625]),
			.NE(gen[1626]),

			.O(gen[1684]),
			.E(gen[1686]),

			.SO(gen[1744]),
			.S(gen[1745]),
			.SE(gen[1746]),

			.SELF(gen[1685]),
			.cell_state(gen[1685])
		); 

/******************* CELL 1686 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1686 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1625]),
			.N(gen[1626]),
			.NE(gen[1627]),

			.O(gen[1685]),
			.E(gen[1687]),

			.SO(gen[1745]),
			.S(gen[1746]),
			.SE(gen[1747]),

			.SELF(gen[1686]),
			.cell_state(gen[1686])
		); 

/******************* CELL 1687 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1687 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1626]),
			.N(gen[1627]),
			.NE(gen[1628]),

			.O(gen[1686]),
			.E(gen[1688]),

			.SO(gen[1746]),
			.S(gen[1747]),
			.SE(gen[1748]),

			.SELF(gen[1687]),
			.cell_state(gen[1687])
		); 

/******************* CELL 1688 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1688 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1627]),
			.N(gen[1628]),
			.NE(gen[1629]),

			.O(gen[1687]),
			.E(gen[1689]),

			.SO(gen[1747]),
			.S(gen[1748]),
			.SE(gen[1749]),

			.SELF(gen[1688]),
			.cell_state(gen[1688])
		); 

/******************* CELL 1689 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1689 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1628]),
			.N(gen[1629]),
			.NE(gen[1630]),

			.O(gen[1688]),
			.E(gen[1690]),

			.SO(gen[1748]),
			.S(gen[1749]),
			.SE(gen[1750]),

			.SELF(gen[1689]),
			.cell_state(gen[1689])
		); 

/******************* CELL 1690 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1690 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1629]),
			.N(gen[1630]),
			.NE(gen[1631]),

			.O(gen[1689]),
			.E(gen[1691]),

			.SO(gen[1749]),
			.S(gen[1750]),
			.SE(gen[1751]),

			.SELF(gen[1690]),
			.cell_state(gen[1690])
		); 

/******************* CELL 1691 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1691 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1630]),
			.N(gen[1631]),
			.NE(gen[1632]),

			.O(gen[1690]),
			.E(gen[1692]),

			.SO(gen[1750]),
			.S(gen[1751]),
			.SE(gen[1752]),

			.SELF(gen[1691]),
			.cell_state(gen[1691])
		); 

/******************* CELL 1692 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1692 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1631]),
			.N(gen[1632]),
			.NE(gen[1633]),

			.O(gen[1691]),
			.E(gen[1693]),

			.SO(gen[1751]),
			.S(gen[1752]),
			.SE(gen[1753]),

			.SELF(gen[1692]),
			.cell_state(gen[1692])
		); 

/******************* CELL 1693 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1693 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1632]),
			.N(gen[1633]),
			.NE(gen[1634]),

			.O(gen[1692]),
			.E(gen[1694]),

			.SO(gen[1752]),
			.S(gen[1753]),
			.SE(gen[1754]),

			.SELF(gen[1693]),
			.cell_state(gen[1693])
		); 

/******************* CELL 1694 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1694 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1633]),
			.N(gen[1634]),
			.NE(gen[1635]),

			.O(gen[1693]),
			.E(gen[1695]),

			.SO(gen[1753]),
			.S(gen[1754]),
			.SE(gen[1755]),

			.SELF(gen[1694]),
			.cell_state(gen[1694])
		); 

/******************* CELL 1695 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1695 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1634]),
			.N(gen[1635]),
			.NE(gen[1636]),

			.O(gen[1694]),
			.E(gen[1696]),

			.SO(gen[1754]),
			.S(gen[1755]),
			.SE(gen[1756]),

			.SELF(gen[1695]),
			.cell_state(gen[1695])
		); 

/******************* CELL 1696 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1696 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1635]),
			.N(gen[1636]),
			.NE(gen[1637]),

			.O(gen[1695]),
			.E(gen[1697]),

			.SO(gen[1755]),
			.S(gen[1756]),
			.SE(gen[1757]),

			.SELF(gen[1696]),
			.cell_state(gen[1696])
		); 

/******************* CELL 1697 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1697 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1636]),
			.N(gen[1637]),
			.NE(gen[1638]),

			.O(gen[1696]),
			.E(gen[1698]),

			.SO(gen[1756]),
			.S(gen[1757]),
			.SE(gen[1758]),

			.SELF(gen[1697]),
			.cell_state(gen[1697])
		); 

/******************* CELL 1698 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1698 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1637]),
			.N(gen[1638]),
			.NE(gen[1639]),

			.O(gen[1697]),
			.E(gen[1699]),

			.SO(gen[1757]),
			.S(gen[1758]),
			.SE(gen[1759]),

			.SELF(gen[1698]),
			.cell_state(gen[1698])
		); 

/******************* CELL 1699 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1699 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1638]),
			.N(gen[1639]),
			.NE(gen[1640]),

			.O(gen[1698]),
			.E(gen[1700]),

			.SO(gen[1758]),
			.S(gen[1759]),
			.SE(gen[1760]),

			.SELF(gen[1699]),
			.cell_state(gen[1699])
		); 

/******************* CELL 1700 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1700 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1639]),
			.N(gen[1640]),
			.NE(gen[1641]),

			.O(gen[1699]),
			.E(gen[1701]),

			.SO(gen[1759]),
			.S(gen[1760]),
			.SE(gen[1761]),

			.SELF(gen[1700]),
			.cell_state(gen[1700])
		); 

/******************* CELL 1701 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1701 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1640]),
			.N(gen[1641]),
			.NE(gen[1642]),

			.O(gen[1700]),
			.E(gen[1702]),

			.SO(gen[1760]),
			.S(gen[1761]),
			.SE(gen[1762]),

			.SELF(gen[1701]),
			.cell_state(gen[1701])
		); 

/******************* CELL 1702 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1702 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1641]),
			.N(gen[1642]),
			.NE(gen[1643]),

			.O(gen[1701]),
			.E(gen[1703]),

			.SO(gen[1761]),
			.S(gen[1762]),
			.SE(gen[1763]),

			.SELF(gen[1702]),
			.cell_state(gen[1702])
		); 

/******************* CELL 1703 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1703 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1642]),
			.N(gen[1643]),
			.NE(gen[1644]),

			.O(gen[1702]),
			.E(gen[1704]),

			.SO(gen[1762]),
			.S(gen[1763]),
			.SE(gen[1764]),

			.SELF(gen[1703]),
			.cell_state(gen[1703])
		); 

/******************* CELL 1704 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1704 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1643]),
			.N(gen[1644]),
			.NE(gen[1645]),

			.O(gen[1703]),
			.E(gen[1705]),

			.SO(gen[1763]),
			.S(gen[1764]),
			.SE(gen[1765]),

			.SELF(gen[1704]),
			.cell_state(gen[1704])
		); 

/******************* CELL 1705 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1705 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1644]),
			.N(gen[1645]),
			.NE(gen[1646]),

			.O(gen[1704]),
			.E(gen[1706]),

			.SO(gen[1764]),
			.S(gen[1765]),
			.SE(gen[1766]),

			.SELF(gen[1705]),
			.cell_state(gen[1705])
		); 

/******************* CELL 1706 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1706 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1645]),
			.N(gen[1646]),
			.NE(gen[1647]),

			.O(gen[1705]),
			.E(gen[1707]),

			.SO(gen[1765]),
			.S(gen[1766]),
			.SE(gen[1767]),

			.SELF(gen[1706]),
			.cell_state(gen[1706])
		); 

/******************* CELL 1707 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1707 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1646]),
			.N(gen[1647]),
			.NE(gen[1648]),

			.O(gen[1706]),
			.E(gen[1708]),

			.SO(gen[1766]),
			.S(gen[1767]),
			.SE(gen[1768]),

			.SELF(gen[1707]),
			.cell_state(gen[1707])
		); 

/******************* CELL 1708 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1708 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1647]),
			.N(gen[1648]),
			.NE(gen[1649]),

			.O(gen[1707]),
			.E(gen[1709]),

			.SO(gen[1767]),
			.S(gen[1768]),
			.SE(gen[1769]),

			.SELF(gen[1708]),
			.cell_state(gen[1708])
		); 

/******************* CELL 1709 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1709 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1648]),
			.N(gen[1649]),
			.NE(gen[1650]),

			.O(gen[1708]),
			.E(gen[1710]),

			.SO(gen[1768]),
			.S(gen[1769]),
			.SE(gen[1770]),

			.SELF(gen[1709]),
			.cell_state(gen[1709])
		); 

/******************* CELL 1710 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1710 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1649]),
			.N(gen[1650]),
			.NE(gen[1651]),

			.O(gen[1709]),
			.E(gen[1711]),

			.SO(gen[1769]),
			.S(gen[1770]),
			.SE(gen[1771]),

			.SELF(gen[1710]),
			.cell_state(gen[1710])
		); 

/******************* CELL 1711 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1711 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1650]),
			.N(gen[1651]),
			.NE(gen[1652]),

			.O(gen[1710]),
			.E(gen[1712]),

			.SO(gen[1770]),
			.S(gen[1771]),
			.SE(gen[1772]),

			.SELF(gen[1711]),
			.cell_state(gen[1711])
		); 

/******************* CELL 1712 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1712 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1651]),
			.N(gen[1652]),
			.NE(gen[1653]),

			.O(gen[1711]),
			.E(gen[1713]),

			.SO(gen[1771]),
			.S(gen[1772]),
			.SE(gen[1773]),

			.SELF(gen[1712]),
			.cell_state(gen[1712])
		); 

/******************* CELL 1713 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1713 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1652]),
			.N(gen[1653]),
			.NE(gen[1654]),

			.O(gen[1712]),
			.E(gen[1714]),

			.SO(gen[1772]),
			.S(gen[1773]),
			.SE(gen[1774]),

			.SELF(gen[1713]),
			.cell_state(gen[1713])
		); 

/******************* CELL 1714 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1714 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1653]),
			.N(gen[1654]),
			.NE(gen[1655]),

			.O(gen[1713]),
			.E(gen[1715]),

			.SO(gen[1773]),
			.S(gen[1774]),
			.SE(gen[1775]),

			.SELF(gen[1714]),
			.cell_state(gen[1714])
		); 

/******************* CELL 1715 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1715 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1654]),
			.N(gen[1655]),
			.NE(gen[1656]),

			.O(gen[1714]),
			.E(gen[1716]),

			.SO(gen[1774]),
			.S(gen[1775]),
			.SE(gen[1776]),

			.SELF(gen[1715]),
			.cell_state(gen[1715])
		); 

/******************* CELL 1716 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1716 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1655]),
			.N(gen[1656]),
			.NE(gen[1657]),

			.O(gen[1715]),
			.E(gen[1717]),

			.SO(gen[1775]),
			.S(gen[1776]),
			.SE(gen[1777]),

			.SELF(gen[1716]),
			.cell_state(gen[1716])
		); 

/******************* CELL 1717 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1717 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1656]),
			.N(gen[1657]),
			.NE(gen[1658]),

			.O(gen[1716]),
			.E(gen[1718]),

			.SO(gen[1776]),
			.S(gen[1777]),
			.SE(gen[1778]),

			.SELF(gen[1717]),
			.cell_state(gen[1717])
		); 

/******************* CELL 1718 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1718 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1657]),
			.N(gen[1658]),
			.NE(gen[1659]),

			.O(gen[1717]),
			.E(gen[1719]),

			.SO(gen[1777]),
			.S(gen[1778]),
			.SE(gen[1779]),

			.SELF(gen[1718]),
			.cell_state(gen[1718])
		); 

/******************* CELL 1719 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1719 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1658]),
			.N(gen[1659]),
			.NE(gen[1660]),

			.O(gen[1718]),
			.E(gen[1720]),

			.SO(gen[1778]),
			.S(gen[1779]),
			.SE(gen[1780]),

			.SELF(gen[1719]),
			.cell_state(gen[1719])
		); 

/******************* CELL 1720 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1720 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1659]),
			.N(gen[1660]),
			.NE(gen[1661]),

			.O(gen[1719]),
			.E(gen[1721]),

			.SO(gen[1779]),
			.S(gen[1780]),
			.SE(gen[1781]),

			.SELF(gen[1720]),
			.cell_state(gen[1720])
		); 

/******************* CELL 1721 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1721 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1660]),
			.N(gen[1661]),
			.NE(gen[1662]),

			.O(gen[1720]),
			.E(gen[1722]),

			.SO(gen[1780]),
			.S(gen[1781]),
			.SE(gen[1782]),

			.SELF(gen[1721]),
			.cell_state(gen[1721])
		); 

/******************* CELL 1722 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1722 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1661]),
			.N(gen[1662]),
			.NE(gen[1663]),

			.O(gen[1721]),
			.E(gen[1723]),

			.SO(gen[1781]),
			.S(gen[1782]),
			.SE(gen[1783]),

			.SELF(gen[1722]),
			.cell_state(gen[1722])
		); 

/******************* CELL 1723 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1723 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1662]),
			.N(gen[1663]),
			.NE(gen[1664]),

			.O(gen[1722]),
			.E(gen[1724]),

			.SO(gen[1782]),
			.S(gen[1783]),
			.SE(gen[1784]),

			.SELF(gen[1723]),
			.cell_state(gen[1723])
		); 

/******************* CELL 1724 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1724 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1663]),
			.N(gen[1664]),
			.NE(gen[1665]),

			.O(gen[1723]),
			.E(gen[1725]),

			.SO(gen[1783]),
			.S(gen[1784]),
			.SE(gen[1785]),

			.SELF(gen[1724]),
			.cell_state(gen[1724])
		); 

/******************* CELL 1725 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1725 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1664]),
			.N(gen[1665]),
			.NE(gen[1666]),

			.O(gen[1724]),
			.E(gen[1726]),

			.SO(gen[1784]),
			.S(gen[1785]),
			.SE(gen[1786]),

			.SELF(gen[1725]),
			.cell_state(gen[1725])
		); 

/******************* CELL 1726 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1726 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1665]),
			.N(gen[1666]),
			.NE(gen[1667]),

			.O(gen[1725]),
			.E(gen[1727]),

			.SO(gen[1785]),
			.S(gen[1786]),
			.SE(gen[1787]),

			.SELF(gen[1726]),
			.cell_state(gen[1726])
		); 

/******************* CELL 1727 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1727 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1666]),
			.N(gen[1667]),
			.NE(gen[1668]),

			.O(gen[1726]),
			.E(gen[1728]),

			.SO(gen[1786]),
			.S(gen[1787]),
			.SE(gen[1788]),

			.SELF(gen[1727]),
			.cell_state(gen[1727])
		); 

/******************* CELL 1728 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1728 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1667]),
			.N(gen[1668]),
			.NE(gen[1669]),

			.O(gen[1727]),
			.E(gen[1729]),

			.SO(gen[1787]),
			.S(gen[1788]),
			.SE(gen[1789]),

			.SELF(gen[1728]),
			.cell_state(gen[1728])
		); 

/******************* CELL 1729 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1729 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1668]),
			.N(gen[1669]),
			.NE(gen[1670]),

			.O(gen[1728]),
			.E(gen[1730]),

			.SO(gen[1788]),
			.S(gen[1789]),
			.SE(gen[1790]),

			.SELF(gen[1729]),
			.cell_state(gen[1729])
		); 

/******************* CELL 1730 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1730 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1669]),
			.N(gen[1670]),
			.NE(gen[1671]),

			.O(gen[1729]),
			.E(gen[1731]),

			.SO(gen[1789]),
			.S(gen[1790]),
			.SE(gen[1791]),

			.SELF(gen[1730]),
			.cell_state(gen[1730])
		); 

/******************* CELL 1731 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1731 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1670]),
			.N(gen[1671]),
			.NE(gen[1672]),

			.O(gen[1730]),
			.E(gen[1732]),

			.SO(gen[1790]),
			.S(gen[1791]),
			.SE(gen[1792]),

			.SELF(gen[1731]),
			.cell_state(gen[1731])
		); 

/******************* CELL 1732 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1732 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1671]),
			.N(gen[1672]),
			.NE(gen[1673]),

			.O(gen[1731]),
			.E(gen[1733]),

			.SO(gen[1791]),
			.S(gen[1792]),
			.SE(gen[1793]),

			.SELF(gen[1732]),
			.cell_state(gen[1732])
		); 

/******************* CELL 1733 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1733 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1672]),
			.N(gen[1673]),
			.NE(gen[1674]),

			.O(gen[1732]),
			.E(gen[1734]),

			.SO(gen[1792]),
			.S(gen[1793]),
			.SE(gen[1794]),

			.SELF(gen[1733]),
			.cell_state(gen[1733])
		); 

/******************* CELL 1734 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1734 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1673]),
			.N(gen[1674]),
			.NE(gen[1675]),

			.O(gen[1733]),
			.E(gen[1735]),

			.SO(gen[1793]),
			.S(gen[1794]),
			.SE(gen[1795]),

			.SELF(gen[1734]),
			.cell_state(gen[1734])
		); 

/******************* CELL 1735 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1735 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1674]),
			.N(gen[1675]),
			.NE(gen[1676]),

			.O(gen[1734]),
			.E(gen[1736]),

			.SO(gen[1794]),
			.S(gen[1795]),
			.SE(gen[1796]),

			.SELF(gen[1735]),
			.cell_state(gen[1735])
		); 

/******************* CELL 1736 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1736 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1675]),
			.N(gen[1676]),
			.NE(gen[1677]),

			.O(gen[1735]),
			.E(gen[1737]),

			.SO(gen[1795]),
			.S(gen[1796]),
			.SE(gen[1797]),

			.SELF(gen[1736]),
			.cell_state(gen[1736])
		); 

/******************* CELL 1737 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1737 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1676]),
			.N(gen[1677]),
			.NE(gen[1678]),

			.O(gen[1736]),
			.E(gen[1738]),

			.SO(gen[1796]),
			.S(gen[1797]),
			.SE(gen[1798]),

			.SELF(gen[1737]),
			.cell_state(gen[1737])
		); 

/******************* CELL 1738 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1738 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1677]),
			.N(gen[1678]),
			.NE(gen[1679]),

			.O(gen[1737]),
			.E(gen[1739]),

			.SO(gen[1797]),
			.S(gen[1798]),
			.SE(gen[1799]),

			.SELF(gen[1738]),
			.cell_state(gen[1738])
		); 

/******************* CELL 1739 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1739 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1678]),
			.N(gen[1679]),
			.NE(gen[1678]),

			.O(gen[1738]),
			.E(gen[1738]),

			.SO(gen[1798]),
			.S(gen[1799]),
			.SE(gen[1798]),

			.SELF(gen[1739]),
			.cell_state(gen[1739])
		); 

/******************* CELL 1740 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1740 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1681]),
			.N(gen[1680]),
			.NE(gen[1681]),

			.O(gen[1741]),
			.E(gen[1741]),

			.SO(gen[1801]),
			.S(gen[1800]),
			.SE(gen[1801]),

			.SELF(gen[1740]),
			.cell_state(gen[1740])
		); 

/******************* CELL 1741 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1741 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1680]),
			.N(gen[1681]),
			.NE(gen[1682]),

			.O(gen[1740]),
			.E(gen[1742]),

			.SO(gen[1800]),
			.S(gen[1801]),
			.SE(gen[1802]),

			.SELF(gen[1741]),
			.cell_state(gen[1741])
		); 

/******************* CELL 1742 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1742 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1681]),
			.N(gen[1682]),
			.NE(gen[1683]),

			.O(gen[1741]),
			.E(gen[1743]),

			.SO(gen[1801]),
			.S(gen[1802]),
			.SE(gen[1803]),

			.SELF(gen[1742]),
			.cell_state(gen[1742])
		); 

/******************* CELL 1743 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1743 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1682]),
			.N(gen[1683]),
			.NE(gen[1684]),

			.O(gen[1742]),
			.E(gen[1744]),

			.SO(gen[1802]),
			.S(gen[1803]),
			.SE(gen[1804]),

			.SELF(gen[1743]),
			.cell_state(gen[1743])
		); 

/******************* CELL 1744 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1744 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1683]),
			.N(gen[1684]),
			.NE(gen[1685]),

			.O(gen[1743]),
			.E(gen[1745]),

			.SO(gen[1803]),
			.S(gen[1804]),
			.SE(gen[1805]),

			.SELF(gen[1744]),
			.cell_state(gen[1744])
		); 

/******************* CELL 1745 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1745 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1684]),
			.N(gen[1685]),
			.NE(gen[1686]),

			.O(gen[1744]),
			.E(gen[1746]),

			.SO(gen[1804]),
			.S(gen[1805]),
			.SE(gen[1806]),

			.SELF(gen[1745]),
			.cell_state(gen[1745])
		); 

/******************* CELL 1746 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1746 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1685]),
			.N(gen[1686]),
			.NE(gen[1687]),

			.O(gen[1745]),
			.E(gen[1747]),

			.SO(gen[1805]),
			.S(gen[1806]),
			.SE(gen[1807]),

			.SELF(gen[1746]),
			.cell_state(gen[1746])
		); 

/******************* CELL 1747 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1747 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1686]),
			.N(gen[1687]),
			.NE(gen[1688]),

			.O(gen[1746]),
			.E(gen[1748]),

			.SO(gen[1806]),
			.S(gen[1807]),
			.SE(gen[1808]),

			.SELF(gen[1747]),
			.cell_state(gen[1747])
		); 

/******************* CELL 1748 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1748 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1687]),
			.N(gen[1688]),
			.NE(gen[1689]),

			.O(gen[1747]),
			.E(gen[1749]),

			.SO(gen[1807]),
			.S(gen[1808]),
			.SE(gen[1809]),

			.SELF(gen[1748]),
			.cell_state(gen[1748])
		); 

/******************* CELL 1749 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1749 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1688]),
			.N(gen[1689]),
			.NE(gen[1690]),

			.O(gen[1748]),
			.E(gen[1750]),

			.SO(gen[1808]),
			.S(gen[1809]),
			.SE(gen[1810]),

			.SELF(gen[1749]),
			.cell_state(gen[1749])
		); 

/******************* CELL 1750 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1750 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1689]),
			.N(gen[1690]),
			.NE(gen[1691]),

			.O(gen[1749]),
			.E(gen[1751]),

			.SO(gen[1809]),
			.S(gen[1810]),
			.SE(gen[1811]),

			.SELF(gen[1750]),
			.cell_state(gen[1750])
		); 

/******************* CELL 1751 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1751 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1690]),
			.N(gen[1691]),
			.NE(gen[1692]),

			.O(gen[1750]),
			.E(gen[1752]),

			.SO(gen[1810]),
			.S(gen[1811]),
			.SE(gen[1812]),

			.SELF(gen[1751]),
			.cell_state(gen[1751])
		); 

/******************* CELL 1752 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1752 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1691]),
			.N(gen[1692]),
			.NE(gen[1693]),

			.O(gen[1751]),
			.E(gen[1753]),

			.SO(gen[1811]),
			.S(gen[1812]),
			.SE(gen[1813]),

			.SELF(gen[1752]),
			.cell_state(gen[1752])
		); 

/******************* CELL 1753 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1753 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1692]),
			.N(gen[1693]),
			.NE(gen[1694]),

			.O(gen[1752]),
			.E(gen[1754]),

			.SO(gen[1812]),
			.S(gen[1813]),
			.SE(gen[1814]),

			.SELF(gen[1753]),
			.cell_state(gen[1753])
		); 

/******************* CELL 1754 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1754 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1693]),
			.N(gen[1694]),
			.NE(gen[1695]),

			.O(gen[1753]),
			.E(gen[1755]),

			.SO(gen[1813]),
			.S(gen[1814]),
			.SE(gen[1815]),

			.SELF(gen[1754]),
			.cell_state(gen[1754])
		); 

/******************* CELL 1755 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1755 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1694]),
			.N(gen[1695]),
			.NE(gen[1696]),

			.O(gen[1754]),
			.E(gen[1756]),

			.SO(gen[1814]),
			.S(gen[1815]),
			.SE(gen[1816]),

			.SELF(gen[1755]),
			.cell_state(gen[1755])
		); 

/******************* CELL 1756 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1756 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1695]),
			.N(gen[1696]),
			.NE(gen[1697]),

			.O(gen[1755]),
			.E(gen[1757]),

			.SO(gen[1815]),
			.S(gen[1816]),
			.SE(gen[1817]),

			.SELF(gen[1756]),
			.cell_state(gen[1756])
		); 

/******************* CELL 1757 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1757 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1696]),
			.N(gen[1697]),
			.NE(gen[1698]),

			.O(gen[1756]),
			.E(gen[1758]),

			.SO(gen[1816]),
			.S(gen[1817]),
			.SE(gen[1818]),

			.SELF(gen[1757]),
			.cell_state(gen[1757])
		); 

/******************* CELL 1758 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1758 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1697]),
			.N(gen[1698]),
			.NE(gen[1699]),

			.O(gen[1757]),
			.E(gen[1759]),

			.SO(gen[1817]),
			.S(gen[1818]),
			.SE(gen[1819]),

			.SELF(gen[1758]),
			.cell_state(gen[1758])
		); 

/******************* CELL 1759 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1759 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1698]),
			.N(gen[1699]),
			.NE(gen[1700]),

			.O(gen[1758]),
			.E(gen[1760]),

			.SO(gen[1818]),
			.S(gen[1819]),
			.SE(gen[1820]),

			.SELF(gen[1759]),
			.cell_state(gen[1759])
		); 

/******************* CELL 1760 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1760 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1699]),
			.N(gen[1700]),
			.NE(gen[1701]),

			.O(gen[1759]),
			.E(gen[1761]),

			.SO(gen[1819]),
			.S(gen[1820]),
			.SE(gen[1821]),

			.SELF(gen[1760]),
			.cell_state(gen[1760])
		); 

/******************* CELL 1761 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1761 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1700]),
			.N(gen[1701]),
			.NE(gen[1702]),

			.O(gen[1760]),
			.E(gen[1762]),

			.SO(gen[1820]),
			.S(gen[1821]),
			.SE(gen[1822]),

			.SELF(gen[1761]),
			.cell_state(gen[1761])
		); 

/******************* CELL 1762 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1762 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1701]),
			.N(gen[1702]),
			.NE(gen[1703]),

			.O(gen[1761]),
			.E(gen[1763]),

			.SO(gen[1821]),
			.S(gen[1822]),
			.SE(gen[1823]),

			.SELF(gen[1762]),
			.cell_state(gen[1762])
		); 

/******************* CELL 1763 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1763 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1702]),
			.N(gen[1703]),
			.NE(gen[1704]),

			.O(gen[1762]),
			.E(gen[1764]),

			.SO(gen[1822]),
			.S(gen[1823]),
			.SE(gen[1824]),

			.SELF(gen[1763]),
			.cell_state(gen[1763])
		); 

/******************* CELL 1764 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1764 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1703]),
			.N(gen[1704]),
			.NE(gen[1705]),

			.O(gen[1763]),
			.E(gen[1765]),

			.SO(gen[1823]),
			.S(gen[1824]),
			.SE(gen[1825]),

			.SELF(gen[1764]),
			.cell_state(gen[1764])
		); 

/******************* CELL 1765 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1765 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1704]),
			.N(gen[1705]),
			.NE(gen[1706]),

			.O(gen[1764]),
			.E(gen[1766]),

			.SO(gen[1824]),
			.S(gen[1825]),
			.SE(gen[1826]),

			.SELF(gen[1765]),
			.cell_state(gen[1765])
		); 

/******************* CELL 1766 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1766 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1705]),
			.N(gen[1706]),
			.NE(gen[1707]),

			.O(gen[1765]),
			.E(gen[1767]),

			.SO(gen[1825]),
			.S(gen[1826]),
			.SE(gen[1827]),

			.SELF(gen[1766]),
			.cell_state(gen[1766])
		); 

/******************* CELL 1767 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1767 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1706]),
			.N(gen[1707]),
			.NE(gen[1708]),

			.O(gen[1766]),
			.E(gen[1768]),

			.SO(gen[1826]),
			.S(gen[1827]),
			.SE(gen[1828]),

			.SELF(gen[1767]),
			.cell_state(gen[1767])
		); 

/******************* CELL 1768 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1768 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1707]),
			.N(gen[1708]),
			.NE(gen[1709]),

			.O(gen[1767]),
			.E(gen[1769]),

			.SO(gen[1827]),
			.S(gen[1828]),
			.SE(gen[1829]),

			.SELF(gen[1768]),
			.cell_state(gen[1768])
		); 

/******************* CELL 1769 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1769 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1708]),
			.N(gen[1709]),
			.NE(gen[1710]),

			.O(gen[1768]),
			.E(gen[1770]),

			.SO(gen[1828]),
			.S(gen[1829]),
			.SE(gen[1830]),

			.SELF(gen[1769]),
			.cell_state(gen[1769])
		); 

/******************* CELL 1770 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1770 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1709]),
			.N(gen[1710]),
			.NE(gen[1711]),

			.O(gen[1769]),
			.E(gen[1771]),

			.SO(gen[1829]),
			.S(gen[1830]),
			.SE(gen[1831]),

			.SELF(gen[1770]),
			.cell_state(gen[1770])
		); 

/******************* CELL 1771 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1771 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1710]),
			.N(gen[1711]),
			.NE(gen[1712]),

			.O(gen[1770]),
			.E(gen[1772]),

			.SO(gen[1830]),
			.S(gen[1831]),
			.SE(gen[1832]),

			.SELF(gen[1771]),
			.cell_state(gen[1771])
		); 

/******************* CELL 1772 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1772 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1711]),
			.N(gen[1712]),
			.NE(gen[1713]),

			.O(gen[1771]),
			.E(gen[1773]),

			.SO(gen[1831]),
			.S(gen[1832]),
			.SE(gen[1833]),

			.SELF(gen[1772]),
			.cell_state(gen[1772])
		); 

/******************* CELL 1773 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1773 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1712]),
			.N(gen[1713]),
			.NE(gen[1714]),

			.O(gen[1772]),
			.E(gen[1774]),

			.SO(gen[1832]),
			.S(gen[1833]),
			.SE(gen[1834]),

			.SELF(gen[1773]),
			.cell_state(gen[1773])
		); 

/******************* CELL 1774 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1774 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1713]),
			.N(gen[1714]),
			.NE(gen[1715]),

			.O(gen[1773]),
			.E(gen[1775]),

			.SO(gen[1833]),
			.S(gen[1834]),
			.SE(gen[1835]),

			.SELF(gen[1774]),
			.cell_state(gen[1774])
		); 

/******************* CELL 1775 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1775 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1714]),
			.N(gen[1715]),
			.NE(gen[1716]),

			.O(gen[1774]),
			.E(gen[1776]),

			.SO(gen[1834]),
			.S(gen[1835]),
			.SE(gen[1836]),

			.SELF(gen[1775]),
			.cell_state(gen[1775])
		); 

/******************* CELL 1776 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1776 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1715]),
			.N(gen[1716]),
			.NE(gen[1717]),

			.O(gen[1775]),
			.E(gen[1777]),

			.SO(gen[1835]),
			.S(gen[1836]),
			.SE(gen[1837]),

			.SELF(gen[1776]),
			.cell_state(gen[1776])
		); 

/******************* CELL 1777 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1777 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1716]),
			.N(gen[1717]),
			.NE(gen[1718]),

			.O(gen[1776]),
			.E(gen[1778]),

			.SO(gen[1836]),
			.S(gen[1837]),
			.SE(gen[1838]),

			.SELF(gen[1777]),
			.cell_state(gen[1777])
		); 

/******************* CELL 1778 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1778 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1717]),
			.N(gen[1718]),
			.NE(gen[1719]),

			.O(gen[1777]),
			.E(gen[1779]),

			.SO(gen[1837]),
			.S(gen[1838]),
			.SE(gen[1839]),

			.SELF(gen[1778]),
			.cell_state(gen[1778])
		); 

/******************* CELL 1779 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1779 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1718]),
			.N(gen[1719]),
			.NE(gen[1720]),

			.O(gen[1778]),
			.E(gen[1780]),

			.SO(gen[1838]),
			.S(gen[1839]),
			.SE(gen[1840]),

			.SELF(gen[1779]),
			.cell_state(gen[1779])
		); 

/******************* CELL 1780 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1780 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1719]),
			.N(gen[1720]),
			.NE(gen[1721]),

			.O(gen[1779]),
			.E(gen[1781]),

			.SO(gen[1839]),
			.S(gen[1840]),
			.SE(gen[1841]),

			.SELF(gen[1780]),
			.cell_state(gen[1780])
		); 

/******************* CELL 1781 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1781 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1720]),
			.N(gen[1721]),
			.NE(gen[1722]),

			.O(gen[1780]),
			.E(gen[1782]),

			.SO(gen[1840]),
			.S(gen[1841]),
			.SE(gen[1842]),

			.SELF(gen[1781]),
			.cell_state(gen[1781])
		); 

/******************* CELL 1782 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1782 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1721]),
			.N(gen[1722]),
			.NE(gen[1723]),

			.O(gen[1781]),
			.E(gen[1783]),

			.SO(gen[1841]),
			.S(gen[1842]),
			.SE(gen[1843]),

			.SELF(gen[1782]),
			.cell_state(gen[1782])
		); 

/******************* CELL 1783 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1783 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1722]),
			.N(gen[1723]),
			.NE(gen[1724]),

			.O(gen[1782]),
			.E(gen[1784]),

			.SO(gen[1842]),
			.S(gen[1843]),
			.SE(gen[1844]),

			.SELF(gen[1783]),
			.cell_state(gen[1783])
		); 

/******************* CELL 1784 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1784 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1723]),
			.N(gen[1724]),
			.NE(gen[1725]),

			.O(gen[1783]),
			.E(gen[1785]),

			.SO(gen[1843]),
			.S(gen[1844]),
			.SE(gen[1845]),

			.SELF(gen[1784]),
			.cell_state(gen[1784])
		); 

/******************* CELL 1785 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1785 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1724]),
			.N(gen[1725]),
			.NE(gen[1726]),

			.O(gen[1784]),
			.E(gen[1786]),

			.SO(gen[1844]),
			.S(gen[1845]),
			.SE(gen[1846]),

			.SELF(gen[1785]),
			.cell_state(gen[1785])
		); 

/******************* CELL 1786 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1786 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1725]),
			.N(gen[1726]),
			.NE(gen[1727]),

			.O(gen[1785]),
			.E(gen[1787]),

			.SO(gen[1845]),
			.S(gen[1846]),
			.SE(gen[1847]),

			.SELF(gen[1786]),
			.cell_state(gen[1786])
		); 

/******************* CELL 1787 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1787 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1726]),
			.N(gen[1727]),
			.NE(gen[1728]),

			.O(gen[1786]),
			.E(gen[1788]),

			.SO(gen[1846]),
			.S(gen[1847]),
			.SE(gen[1848]),

			.SELF(gen[1787]),
			.cell_state(gen[1787])
		); 

/******************* CELL 1788 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1788 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1727]),
			.N(gen[1728]),
			.NE(gen[1729]),

			.O(gen[1787]),
			.E(gen[1789]),

			.SO(gen[1847]),
			.S(gen[1848]),
			.SE(gen[1849]),

			.SELF(gen[1788]),
			.cell_state(gen[1788])
		); 

/******************* CELL 1789 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1789 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1728]),
			.N(gen[1729]),
			.NE(gen[1730]),

			.O(gen[1788]),
			.E(gen[1790]),

			.SO(gen[1848]),
			.S(gen[1849]),
			.SE(gen[1850]),

			.SELF(gen[1789]),
			.cell_state(gen[1789])
		); 

/******************* CELL 1790 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1790 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1729]),
			.N(gen[1730]),
			.NE(gen[1731]),

			.O(gen[1789]),
			.E(gen[1791]),

			.SO(gen[1849]),
			.S(gen[1850]),
			.SE(gen[1851]),

			.SELF(gen[1790]),
			.cell_state(gen[1790])
		); 

/******************* CELL 1791 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1791 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1730]),
			.N(gen[1731]),
			.NE(gen[1732]),

			.O(gen[1790]),
			.E(gen[1792]),

			.SO(gen[1850]),
			.S(gen[1851]),
			.SE(gen[1852]),

			.SELF(gen[1791]),
			.cell_state(gen[1791])
		); 

/******************* CELL 1792 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1792 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1731]),
			.N(gen[1732]),
			.NE(gen[1733]),

			.O(gen[1791]),
			.E(gen[1793]),

			.SO(gen[1851]),
			.S(gen[1852]),
			.SE(gen[1853]),

			.SELF(gen[1792]),
			.cell_state(gen[1792])
		); 

/******************* CELL 1793 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1793 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1732]),
			.N(gen[1733]),
			.NE(gen[1734]),

			.O(gen[1792]),
			.E(gen[1794]),

			.SO(gen[1852]),
			.S(gen[1853]),
			.SE(gen[1854]),

			.SELF(gen[1793]),
			.cell_state(gen[1793])
		); 

/******************* CELL 1794 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1794 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1733]),
			.N(gen[1734]),
			.NE(gen[1735]),

			.O(gen[1793]),
			.E(gen[1795]),

			.SO(gen[1853]),
			.S(gen[1854]),
			.SE(gen[1855]),

			.SELF(gen[1794]),
			.cell_state(gen[1794])
		); 

/******************* CELL 1795 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1795 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1734]),
			.N(gen[1735]),
			.NE(gen[1736]),

			.O(gen[1794]),
			.E(gen[1796]),

			.SO(gen[1854]),
			.S(gen[1855]),
			.SE(gen[1856]),

			.SELF(gen[1795]),
			.cell_state(gen[1795])
		); 

/******************* CELL 1796 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1796 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1735]),
			.N(gen[1736]),
			.NE(gen[1737]),

			.O(gen[1795]),
			.E(gen[1797]),

			.SO(gen[1855]),
			.S(gen[1856]),
			.SE(gen[1857]),

			.SELF(gen[1796]),
			.cell_state(gen[1796])
		); 

/******************* CELL 1797 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1797 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1736]),
			.N(gen[1737]),
			.NE(gen[1738]),

			.O(gen[1796]),
			.E(gen[1798]),

			.SO(gen[1856]),
			.S(gen[1857]),
			.SE(gen[1858]),

			.SELF(gen[1797]),
			.cell_state(gen[1797])
		); 

/******************* CELL 1798 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1798 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1737]),
			.N(gen[1738]),
			.NE(gen[1739]),

			.O(gen[1797]),
			.E(gen[1799]),

			.SO(gen[1857]),
			.S(gen[1858]),
			.SE(gen[1859]),

			.SELF(gen[1798]),
			.cell_state(gen[1798])
		); 

/******************* CELL 1799 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1799 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1738]),
			.N(gen[1739]),
			.NE(gen[1738]),

			.O(gen[1798]),
			.E(gen[1798]),

			.SO(gen[1858]),
			.S(gen[1859]),
			.SE(gen[1858]),

			.SELF(gen[1799]),
			.cell_state(gen[1799])
		); 

/******************* CELL 1800 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1800 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1741]),
			.N(gen[1740]),
			.NE(gen[1741]),

			.O(gen[1801]),
			.E(gen[1801]),

			.SO(gen[1861]),
			.S(gen[1860]),
			.SE(gen[1861]),

			.SELF(gen[1800]),
			.cell_state(gen[1800])
		); 

/******************* CELL 1801 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1801 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1740]),
			.N(gen[1741]),
			.NE(gen[1742]),

			.O(gen[1800]),
			.E(gen[1802]),

			.SO(gen[1860]),
			.S(gen[1861]),
			.SE(gen[1862]),

			.SELF(gen[1801]),
			.cell_state(gen[1801])
		); 

/******************* CELL 1802 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1802 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1741]),
			.N(gen[1742]),
			.NE(gen[1743]),

			.O(gen[1801]),
			.E(gen[1803]),

			.SO(gen[1861]),
			.S(gen[1862]),
			.SE(gen[1863]),

			.SELF(gen[1802]),
			.cell_state(gen[1802])
		); 

/******************* CELL 1803 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1803 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1742]),
			.N(gen[1743]),
			.NE(gen[1744]),

			.O(gen[1802]),
			.E(gen[1804]),

			.SO(gen[1862]),
			.S(gen[1863]),
			.SE(gen[1864]),

			.SELF(gen[1803]),
			.cell_state(gen[1803])
		); 

/******************* CELL 1804 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1804 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1743]),
			.N(gen[1744]),
			.NE(gen[1745]),

			.O(gen[1803]),
			.E(gen[1805]),

			.SO(gen[1863]),
			.S(gen[1864]),
			.SE(gen[1865]),

			.SELF(gen[1804]),
			.cell_state(gen[1804])
		); 

/******************* CELL 1805 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1805 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1744]),
			.N(gen[1745]),
			.NE(gen[1746]),

			.O(gen[1804]),
			.E(gen[1806]),

			.SO(gen[1864]),
			.S(gen[1865]),
			.SE(gen[1866]),

			.SELF(gen[1805]),
			.cell_state(gen[1805])
		); 

/******************* CELL 1806 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1806 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1745]),
			.N(gen[1746]),
			.NE(gen[1747]),

			.O(gen[1805]),
			.E(gen[1807]),

			.SO(gen[1865]),
			.S(gen[1866]),
			.SE(gen[1867]),

			.SELF(gen[1806]),
			.cell_state(gen[1806])
		); 

/******************* CELL 1807 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1807 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1746]),
			.N(gen[1747]),
			.NE(gen[1748]),

			.O(gen[1806]),
			.E(gen[1808]),

			.SO(gen[1866]),
			.S(gen[1867]),
			.SE(gen[1868]),

			.SELF(gen[1807]),
			.cell_state(gen[1807])
		); 

/******************* CELL 1808 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1808 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1747]),
			.N(gen[1748]),
			.NE(gen[1749]),

			.O(gen[1807]),
			.E(gen[1809]),

			.SO(gen[1867]),
			.S(gen[1868]),
			.SE(gen[1869]),

			.SELF(gen[1808]),
			.cell_state(gen[1808])
		); 

/******************* CELL 1809 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1809 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1748]),
			.N(gen[1749]),
			.NE(gen[1750]),

			.O(gen[1808]),
			.E(gen[1810]),

			.SO(gen[1868]),
			.S(gen[1869]),
			.SE(gen[1870]),

			.SELF(gen[1809]),
			.cell_state(gen[1809])
		); 

/******************* CELL 1810 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1810 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1749]),
			.N(gen[1750]),
			.NE(gen[1751]),

			.O(gen[1809]),
			.E(gen[1811]),

			.SO(gen[1869]),
			.S(gen[1870]),
			.SE(gen[1871]),

			.SELF(gen[1810]),
			.cell_state(gen[1810])
		); 

/******************* CELL 1811 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1811 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1750]),
			.N(gen[1751]),
			.NE(gen[1752]),

			.O(gen[1810]),
			.E(gen[1812]),

			.SO(gen[1870]),
			.S(gen[1871]),
			.SE(gen[1872]),

			.SELF(gen[1811]),
			.cell_state(gen[1811])
		); 

/******************* CELL 1812 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1812 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1751]),
			.N(gen[1752]),
			.NE(gen[1753]),

			.O(gen[1811]),
			.E(gen[1813]),

			.SO(gen[1871]),
			.S(gen[1872]),
			.SE(gen[1873]),

			.SELF(gen[1812]),
			.cell_state(gen[1812])
		); 

/******************* CELL 1813 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1813 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1752]),
			.N(gen[1753]),
			.NE(gen[1754]),

			.O(gen[1812]),
			.E(gen[1814]),

			.SO(gen[1872]),
			.S(gen[1873]),
			.SE(gen[1874]),

			.SELF(gen[1813]),
			.cell_state(gen[1813])
		); 

/******************* CELL 1814 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1814 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1753]),
			.N(gen[1754]),
			.NE(gen[1755]),

			.O(gen[1813]),
			.E(gen[1815]),

			.SO(gen[1873]),
			.S(gen[1874]),
			.SE(gen[1875]),

			.SELF(gen[1814]),
			.cell_state(gen[1814])
		); 

/******************* CELL 1815 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1815 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1754]),
			.N(gen[1755]),
			.NE(gen[1756]),

			.O(gen[1814]),
			.E(gen[1816]),

			.SO(gen[1874]),
			.S(gen[1875]),
			.SE(gen[1876]),

			.SELF(gen[1815]),
			.cell_state(gen[1815])
		); 

/******************* CELL 1816 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1816 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1755]),
			.N(gen[1756]),
			.NE(gen[1757]),

			.O(gen[1815]),
			.E(gen[1817]),

			.SO(gen[1875]),
			.S(gen[1876]),
			.SE(gen[1877]),

			.SELF(gen[1816]),
			.cell_state(gen[1816])
		); 

/******************* CELL 1817 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1817 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1756]),
			.N(gen[1757]),
			.NE(gen[1758]),

			.O(gen[1816]),
			.E(gen[1818]),

			.SO(gen[1876]),
			.S(gen[1877]),
			.SE(gen[1878]),

			.SELF(gen[1817]),
			.cell_state(gen[1817])
		); 

/******************* CELL 1818 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1818 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1757]),
			.N(gen[1758]),
			.NE(gen[1759]),

			.O(gen[1817]),
			.E(gen[1819]),

			.SO(gen[1877]),
			.S(gen[1878]),
			.SE(gen[1879]),

			.SELF(gen[1818]),
			.cell_state(gen[1818])
		); 

/******************* CELL 1819 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1819 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1758]),
			.N(gen[1759]),
			.NE(gen[1760]),

			.O(gen[1818]),
			.E(gen[1820]),

			.SO(gen[1878]),
			.S(gen[1879]),
			.SE(gen[1880]),

			.SELF(gen[1819]),
			.cell_state(gen[1819])
		); 

/******************* CELL 1820 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1820 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1759]),
			.N(gen[1760]),
			.NE(gen[1761]),

			.O(gen[1819]),
			.E(gen[1821]),

			.SO(gen[1879]),
			.S(gen[1880]),
			.SE(gen[1881]),

			.SELF(gen[1820]),
			.cell_state(gen[1820])
		); 

/******************* CELL 1821 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1821 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1760]),
			.N(gen[1761]),
			.NE(gen[1762]),

			.O(gen[1820]),
			.E(gen[1822]),

			.SO(gen[1880]),
			.S(gen[1881]),
			.SE(gen[1882]),

			.SELF(gen[1821]),
			.cell_state(gen[1821])
		); 

/******************* CELL 1822 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1822 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1761]),
			.N(gen[1762]),
			.NE(gen[1763]),

			.O(gen[1821]),
			.E(gen[1823]),

			.SO(gen[1881]),
			.S(gen[1882]),
			.SE(gen[1883]),

			.SELF(gen[1822]),
			.cell_state(gen[1822])
		); 

/******************* CELL 1823 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1823 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1762]),
			.N(gen[1763]),
			.NE(gen[1764]),

			.O(gen[1822]),
			.E(gen[1824]),

			.SO(gen[1882]),
			.S(gen[1883]),
			.SE(gen[1884]),

			.SELF(gen[1823]),
			.cell_state(gen[1823])
		); 

/******************* CELL 1824 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1824 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1763]),
			.N(gen[1764]),
			.NE(gen[1765]),

			.O(gen[1823]),
			.E(gen[1825]),

			.SO(gen[1883]),
			.S(gen[1884]),
			.SE(gen[1885]),

			.SELF(gen[1824]),
			.cell_state(gen[1824])
		); 

/******************* CELL 1825 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1825 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1764]),
			.N(gen[1765]),
			.NE(gen[1766]),

			.O(gen[1824]),
			.E(gen[1826]),

			.SO(gen[1884]),
			.S(gen[1885]),
			.SE(gen[1886]),

			.SELF(gen[1825]),
			.cell_state(gen[1825])
		); 

/******************* CELL 1826 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1826 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1765]),
			.N(gen[1766]),
			.NE(gen[1767]),

			.O(gen[1825]),
			.E(gen[1827]),

			.SO(gen[1885]),
			.S(gen[1886]),
			.SE(gen[1887]),

			.SELF(gen[1826]),
			.cell_state(gen[1826])
		); 

/******************* CELL 1827 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1827 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1766]),
			.N(gen[1767]),
			.NE(gen[1768]),

			.O(gen[1826]),
			.E(gen[1828]),

			.SO(gen[1886]),
			.S(gen[1887]),
			.SE(gen[1888]),

			.SELF(gen[1827]),
			.cell_state(gen[1827])
		); 

/******************* CELL 1828 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1828 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1767]),
			.N(gen[1768]),
			.NE(gen[1769]),

			.O(gen[1827]),
			.E(gen[1829]),

			.SO(gen[1887]),
			.S(gen[1888]),
			.SE(gen[1889]),

			.SELF(gen[1828]),
			.cell_state(gen[1828])
		); 

/******************* CELL 1829 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1829 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1768]),
			.N(gen[1769]),
			.NE(gen[1770]),

			.O(gen[1828]),
			.E(gen[1830]),

			.SO(gen[1888]),
			.S(gen[1889]),
			.SE(gen[1890]),

			.SELF(gen[1829]),
			.cell_state(gen[1829])
		); 

/******************* CELL 1830 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1830 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1769]),
			.N(gen[1770]),
			.NE(gen[1771]),

			.O(gen[1829]),
			.E(gen[1831]),

			.SO(gen[1889]),
			.S(gen[1890]),
			.SE(gen[1891]),

			.SELF(gen[1830]),
			.cell_state(gen[1830])
		); 

/******************* CELL 1831 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1831 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1770]),
			.N(gen[1771]),
			.NE(gen[1772]),

			.O(gen[1830]),
			.E(gen[1832]),

			.SO(gen[1890]),
			.S(gen[1891]),
			.SE(gen[1892]),

			.SELF(gen[1831]),
			.cell_state(gen[1831])
		); 

/******************* CELL 1832 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1832 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1771]),
			.N(gen[1772]),
			.NE(gen[1773]),

			.O(gen[1831]),
			.E(gen[1833]),

			.SO(gen[1891]),
			.S(gen[1892]),
			.SE(gen[1893]),

			.SELF(gen[1832]),
			.cell_state(gen[1832])
		); 

/******************* CELL 1833 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1833 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1772]),
			.N(gen[1773]),
			.NE(gen[1774]),

			.O(gen[1832]),
			.E(gen[1834]),

			.SO(gen[1892]),
			.S(gen[1893]),
			.SE(gen[1894]),

			.SELF(gen[1833]),
			.cell_state(gen[1833])
		); 

/******************* CELL 1834 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1834 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1773]),
			.N(gen[1774]),
			.NE(gen[1775]),

			.O(gen[1833]),
			.E(gen[1835]),

			.SO(gen[1893]),
			.S(gen[1894]),
			.SE(gen[1895]),

			.SELF(gen[1834]),
			.cell_state(gen[1834])
		); 

/******************* CELL 1835 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1835 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1774]),
			.N(gen[1775]),
			.NE(gen[1776]),

			.O(gen[1834]),
			.E(gen[1836]),

			.SO(gen[1894]),
			.S(gen[1895]),
			.SE(gen[1896]),

			.SELF(gen[1835]),
			.cell_state(gen[1835])
		); 

/******************* CELL 1836 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1836 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1775]),
			.N(gen[1776]),
			.NE(gen[1777]),

			.O(gen[1835]),
			.E(gen[1837]),

			.SO(gen[1895]),
			.S(gen[1896]),
			.SE(gen[1897]),

			.SELF(gen[1836]),
			.cell_state(gen[1836])
		); 

/******************* CELL 1837 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1837 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1776]),
			.N(gen[1777]),
			.NE(gen[1778]),

			.O(gen[1836]),
			.E(gen[1838]),

			.SO(gen[1896]),
			.S(gen[1897]),
			.SE(gen[1898]),

			.SELF(gen[1837]),
			.cell_state(gen[1837])
		); 

/******************* CELL 1838 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1838 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1777]),
			.N(gen[1778]),
			.NE(gen[1779]),

			.O(gen[1837]),
			.E(gen[1839]),

			.SO(gen[1897]),
			.S(gen[1898]),
			.SE(gen[1899]),

			.SELF(gen[1838]),
			.cell_state(gen[1838])
		); 

/******************* CELL 1839 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1839 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1778]),
			.N(gen[1779]),
			.NE(gen[1780]),

			.O(gen[1838]),
			.E(gen[1840]),

			.SO(gen[1898]),
			.S(gen[1899]),
			.SE(gen[1900]),

			.SELF(gen[1839]),
			.cell_state(gen[1839])
		); 

/******************* CELL 1840 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1840 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1779]),
			.N(gen[1780]),
			.NE(gen[1781]),

			.O(gen[1839]),
			.E(gen[1841]),

			.SO(gen[1899]),
			.S(gen[1900]),
			.SE(gen[1901]),

			.SELF(gen[1840]),
			.cell_state(gen[1840])
		); 

/******************* CELL 1841 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1841 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1780]),
			.N(gen[1781]),
			.NE(gen[1782]),

			.O(gen[1840]),
			.E(gen[1842]),

			.SO(gen[1900]),
			.S(gen[1901]),
			.SE(gen[1902]),

			.SELF(gen[1841]),
			.cell_state(gen[1841])
		); 

/******************* CELL 1842 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1842 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1781]),
			.N(gen[1782]),
			.NE(gen[1783]),

			.O(gen[1841]),
			.E(gen[1843]),

			.SO(gen[1901]),
			.S(gen[1902]),
			.SE(gen[1903]),

			.SELF(gen[1842]),
			.cell_state(gen[1842])
		); 

/******************* CELL 1843 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1843 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1782]),
			.N(gen[1783]),
			.NE(gen[1784]),

			.O(gen[1842]),
			.E(gen[1844]),

			.SO(gen[1902]),
			.S(gen[1903]),
			.SE(gen[1904]),

			.SELF(gen[1843]),
			.cell_state(gen[1843])
		); 

/******************* CELL 1844 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1844 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1783]),
			.N(gen[1784]),
			.NE(gen[1785]),

			.O(gen[1843]),
			.E(gen[1845]),

			.SO(gen[1903]),
			.S(gen[1904]),
			.SE(gen[1905]),

			.SELF(gen[1844]),
			.cell_state(gen[1844])
		); 

/******************* CELL 1845 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1845 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1784]),
			.N(gen[1785]),
			.NE(gen[1786]),

			.O(gen[1844]),
			.E(gen[1846]),

			.SO(gen[1904]),
			.S(gen[1905]),
			.SE(gen[1906]),

			.SELF(gen[1845]),
			.cell_state(gen[1845])
		); 

/******************* CELL 1846 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1846 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1785]),
			.N(gen[1786]),
			.NE(gen[1787]),

			.O(gen[1845]),
			.E(gen[1847]),

			.SO(gen[1905]),
			.S(gen[1906]),
			.SE(gen[1907]),

			.SELF(gen[1846]),
			.cell_state(gen[1846])
		); 

/******************* CELL 1847 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1847 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1786]),
			.N(gen[1787]),
			.NE(gen[1788]),

			.O(gen[1846]),
			.E(gen[1848]),

			.SO(gen[1906]),
			.S(gen[1907]),
			.SE(gen[1908]),

			.SELF(gen[1847]),
			.cell_state(gen[1847])
		); 

/******************* CELL 1848 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1848 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1787]),
			.N(gen[1788]),
			.NE(gen[1789]),

			.O(gen[1847]),
			.E(gen[1849]),

			.SO(gen[1907]),
			.S(gen[1908]),
			.SE(gen[1909]),

			.SELF(gen[1848]),
			.cell_state(gen[1848])
		); 

/******************* CELL 1849 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1849 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1788]),
			.N(gen[1789]),
			.NE(gen[1790]),

			.O(gen[1848]),
			.E(gen[1850]),

			.SO(gen[1908]),
			.S(gen[1909]),
			.SE(gen[1910]),

			.SELF(gen[1849]),
			.cell_state(gen[1849])
		); 

/******************* CELL 1850 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1850 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1789]),
			.N(gen[1790]),
			.NE(gen[1791]),

			.O(gen[1849]),
			.E(gen[1851]),

			.SO(gen[1909]),
			.S(gen[1910]),
			.SE(gen[1911]),

			.SELF(gen[1850]),
			.cell_state(gen[1850])
		); 

/******************* CELL 1851 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1851 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1790]),
			.N(gen[1791]),
			.NE(gen[1792]),

			.O(gen[1850]),
			.E(gen[1852]),

			.SO(gen[1910]),
			.S(gen[1911]),
			.SE(gen[1912]),

			.SELF(gen[1851]),
			.cell_state(gen[1851])
		); 

/******************* CELL 1852 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1852 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1791]),
			.N(gen[1792]),
			.NE(gen[1793]),

			.O(gen[1851]),
			.E(gen[1853]),

			.SO(gen[1911]),
			.S(gen[1912]),
			.SE(gen[1913]),

			.SELF(gen[1852]),
			.cell_state(gen[1852])
		); 

/******************* CELL 1853 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1853 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1792]),
			.N(gen[1793]),
			.NE(gen[1794]),

			.O(gen[1852]),
			.E(gen[1854]),

			.SO(gen[1912]),
			.S(gen[1913]),
			.SE(gen[1914]),

			.SELF(gen[1853]),
			.cell_state(gen[1853])
		); 

/******************* CELL 1854 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1854 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1793]),
			.N(gen[1794]),
			.NE(gen[1795]),

			.O(gen[1853]),
			.E(gen[1855]),

			.SO(gen[1913]),
			.S(gen[1914]),
			.SE(gen[1915]),

			.SELF(gen[1854]),
			.cell_state(gen[1854])
		); 

/******************* CELL 1855 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1855 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1794]),
			.N(gen[1795]),
			.NE(gen[1796]),

			.O(gen[1854]),
			.E(gen[1856]),

			.SO(gen[1914]),
			.S(gen[1915]),
			.SE(gen[1916]),

			.SELF(gen[1855]),
			.cell_state(gen[1855])
		); 

/******************* CELL 1856 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1856 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1795]),
			.N(gen[1796]),
			.NE(gen[1797]),

			.O(gen[1855]),
			.E(gen[1857]),

			.SO(gen[1915]),
			.S(gen[1916]),
			.SE(gen[1917]),

			.SELF(gen[1856]),
			.cell_state(gen[1856])
		); 

/******************* CELL 1857 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1857 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1796]),
			.N(gen[1797]),
			.NE(gen[1798]),

			.O(gen[1856]),
			.E(gen[1858]),

			.SO(gen[1916]),
			.S(gen[1917]),
			.SE(gen[1918]),

			.SELF(gen[1857]),
			.cell_state(gen[1857])
		); 

/******************* CELL 1858 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1858 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1797]),
			.N(gen[1798]),
			.NE(gen[1799]),

			.O(gen[1857]),
			.E(gen[1859]),

			.SO(gen[1917]),
			.S(gen[1918]),
			.SE(gen[1919]),

			.SELF(gen[1858]),
			.cell_state(gen[1858])
		); 

/******************* CELL 1859 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1859 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1798]),
			.N(gen[1799]),
			.NE(gen[1798]),

			.O(gen[1858]),
			.E(gen[1858]),

			.SO(gen[1918]),
			.S(gen[1919]),
			.SE(gen[1918]),

			.SELF(gen[1859]),
			.cell_state(gen[1859])
		); 

/******************* CELL 1860 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1860 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1801]),
			.N(gen[1800]),
			.NE(gen[1801]),

			.O(gen[1861]),
			.E(gen[1861]),

			.SO(gen[1921]),
			.S(gen[1920]),
			.SE(gen[1921]),

			.SELF(gen[1860]),
			.cell_state(gen[1860])
		); 

/******************* CELL 1861 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1861 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1800]),
			.N(gen[1801]),
			.NE(gen[1802]),

			.O(gen[1860]),
			.E(gen[1862]),

			.SO(gen[1920]),
			.S(gen[1921]),
			.SE(gen[1922]),

			.SELF(gen[1861]),
			.cell_state(gen[1861])
		); 

/******************* CELL 1862 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1862 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1801]),
			.N(gen[1802]),
			.NE(gen[1803]),

			.O(gen[1861]),
			.E(gen[1863]),

			.SO(gen[1921]),
			.S(gen[1922]),
			.SE(gen[1923]),

			.SELF(gen[1862]),
			.cell_state(gen[1862])
		); 

/******************* CELL 1863 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1863 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1802]),
			.N(gen[1803]),
			.NE(gen[1804]),

			.O(gen[1862]),
			.E(gen[1864]),

			.SO(gen[1922]),
			.S(gen[1923]),
			.SE(gen[1924]),

			.SELF(gen[1863]),
			.cell_state(gen[1863])
		); 

/******************* CELL 1864 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1864 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1803]),
			.N(gen[1804]),
			.NE(gen[1805]),

			.O(gen[1863]),
			.E(gen[1865]),

			.SO(gen[1923]),
			.S(gen[1924]),
			.SE(gen[1925]),

			.SELF(gen[1864]),
			.cell_state(gen[1864])
		); 

/******************* CELL 1865 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1865 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1804]),
			.N(gen[1805]),
			.NE(gen[1806]),

			.O(gen[1864]),
			.E(gen[1866]),

			.SO(gen[1924]),
			.S(gen[1925]),
			.SE(gen[1926]),

			.SELF(gen[1865]),
			.cell_state(gen[1865])
		); 

/******************* CELL 1866 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1866 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1805]),
			.N(gen[1806]),
			.NE(gen[1807]),

			.O(gen[1865]),
			.E(gen[1867]),

			.SO(gen[1925]),
			.S(gen[1926]),
			.SE(gen[1927]),

			.SELF(gen[1866]),
			.cell_state(gen[1866])
		); 

/******************* CELL 1867 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1867 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1806]),
			.N(gen[1807]),
			.NE(gen[1808]),

			.O(gen[1866]),
			.E(gen[1868]),

			.SO(gen[1926]),
			.S(gen[1927]),
			.SE(gen[1928]),

			.SELF(gen[1867]),
			.cell_state(gen[1867])
		); 

/******************* CELL 1868 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1868 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1807]),
			.N(gen[1808]),
			.NE(gen[1809]),

			.O(gen[1867]),
			.E(gen[1869]),

			.SO(gen[1927]),
			.S(gen[1928]),
			.SE(gen[1929]),

			.SELF(gen[1868]),
			.cell_state(gen[1868])
		); 

/******************* CELL 1869 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1869 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1808]),
			.N(gen[1809]),
			.NE(gen[1810]),

			.O(gen[1868]),
			.E(gen[1870]),

			.SO(gen[1928]),
			.S(gen[1929]),
			.SE(gen[1930]),

			.SELF(gen[1869]),
			.cell_state(gen[1869])
		); 

/******************* CELL 1870 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1870 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1809]),
			.N(gen[1810]),
			.NE(gen[1811]),

			.O(gen[1869]),
			.E(gen[1871]),

			.SO(gen[1929]),
			.S(gen[1930]),
			.SE(gen[1931]),

			.SELF(gen[1870]),
			.cell_state(gen[1870])
		); 

/******************* CELL 1871 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1871 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1810]),
			.N(gen[1811]),
			.NE(gen[1812]),

			.O(gen[1870]),
			.E(gen[1872]),

			.SO(gen[1930]),
			.S(gen[1931]),
			.SE(gen[1932]),

			.SELF(gen[1871]),
			.cell_state(gen[1871])
		); 

/******************* CELL 1872 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1872 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1811]),
			.N(gen[1812]),
			.NE(gen[1813]),

			.O(gen[1871]),
			.E(gen[1873]),

			.SO(gen[1931]),
			.S(gen[1932]),
			.SE(gen[1933]),

			.SELF(gen[1872]),
			.cell_state(gen[1872])
		); 

/******************* CELL 1873 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1873 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1812]),
			.N(gen[1813]),
			.NE(gen[1814]),

			.O(gen[1872]),
			.E(gen[1874]),

			.SO(gen[1932]),
			.S(gen[1933]),
			.SE(gen[1934]),

			.SELF(gen[1873]),
			.cell_state(gen[1873])
		); 

/******************* CELL 1874 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1874 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1813]),
			.N(gen[1814]),
			.NE(gen[1815]),

			.O(gen[1873]),
			.E(gen[1875]),

			.SO(gen[1933]),
			.S(gen[1934]),
			.SE(gen[1935]),

			.SELF(gen[1874]),
			.cell_state(gen[1874])
		); 

/******************* CELL 1875 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1875 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1814]),
			.N(gen[1815]),
			.NE(gen[1816]),

			.O(gen[1874]),
			.E(gen[1876]),

			.SO(gen[1934]),
			.S(gen[1935]),
			.SE(gen[1936]),

			.SELF(gen[1875]),
			.cell_state(gen[1875])
		); 

/******************* CELL 1876 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1876 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1815]),
			.N(gen[1816]),
			.NE(gen[1817]),

			.O(gen[1875]),
			.E(gen[1877]),

			.SO(gen[1935]),
			.S(gen[1936]),
			.SE(gen[1937]),

			.SELF(gen[1876]),
			.cell_state(gen[1876])
		); 

/******************* CELL 1877 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1877 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1816]),
			.N(gen[1817]),
			.NE(gen[1818]),

			.O(gen[1876]),
			.E(gen[1878]),

			.SO(gen[1936]),
			.S(gen[1937]),
			.SE(gen[1938]),

			.SELF(gen[1877]),
			.cell_state(gen[1877])
		); 

/******************* CELL 1878 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1878 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1817]),
			.N(gen[1818]),
			.NE(gen[1819]),

			.O(gen[1877]),
			.E(gen[1879]),

			.SO(gen[1937]),
			.S(gen[1938]),
			.SE(gen[1939]),

			.SELF(gen[1878]),
			.cell_state(gen[1878])
		); 

/******************* CELL 1879 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1879 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1818]),
			.N(gen[1819]),
			.NE(gen[1820]),

			.O(gen[1878]),
			.E(gen[1880]),

			.SO(gen[1938]),
			.S(gen[1939]),
			.SE(gen[1940]),

			.SELF(gen[1879]),
			.cell_state(gen[1879])
		); 

/******************* CELL 1880 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1880 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1819]),
			.N(gen[1820]),
			.NE(gen[1821]),

			.O(gen[1879]),
			.E(gen[1881]),

			.SO(gen[1939]),
			.S(gen[1940]),
			.SE(gen[1941]),

			.SELF(gen[1880]),
			.cell_state(gen[1880])
		); 

/******************* CELL 1881 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1881 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1820]),
			.N(gen[1821]),
			.NE(gen[1822]),

			.O(gen[1880]),
			.E(gen[1882]),

			.SO(gen[1940]),
			.S(gen[1941]),
			.SE(gen[1942]),

			.SELF(gen[1881]),
			.cell_state(gen[1881])
		); 

/******************* CELL 1882 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1882 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1821]),
			.N(gen[1822]),
			.NE(gen[1823]),

			.O(gen[1881]),
			.E(gen[1883]),

			.SO(gen[1941]),
			.S(gen[1942]),
			.SE(gen[1943]),

			.SELF(gen[1882]),
			.cell_state(gen[1882])
		); 

/******************* CELL 1883 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1883 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1822]),
			.N(gen[1823]),
			.NE(gen[1824]),

			.O(gen[1882]),
			.E(gen[1884]),

			.SO(gen[1942]),
			.S(gen[1943]),
			.SE(gen[1944]),

			.SELF(gen[1883]),
			.cell_state(gen[1883])
		); 

/******************* CELL 1884 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1884 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1823]),
			.N(gen[1824]),
			.NE(gen[1825]),

			.O(gen[1883]),
			.E(gen[1885]),

			.SO(gen[1943]),
			.S(gen[1944]),
			.SE(gen[1945]),

			.SELF(gen[1884]),
			.cell_state(gen[1884])
		); 

/******************* CELL 1885 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1885 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1824]),
			.N(gen[1825]),
			.NE(gen[1826]),

			.O(gen[1884]),
			.E(gen[1886]),

			.SO(gen[1944]),
			.S(gen[1945]),
			.SE(gen[1946]),

			.SELF(gen[1885]),
			.cell_state(gen[1885])
		); 

/******************* CELL 1886 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1886 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1825]),
			.N(gen[1826]),
			.NE(gen[1827]),

			.O(gen[1885]),
			.E(gen[1887]),

			.SO(gen[1945]),
			.S(gen[1946]),
			.SE(gen[1947]),

			.SELF(gen[1886]),
			.cell_state(gen[1886])
		); 

/******************* CELL 1887 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1887 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1826]),
			.N(gen[1827]),
			.NE(gen[1828]),

			.O(gen[1886]),
			.E(gen[1888]),

			.SO(gen[1946]),
			.S(gen[1947]),
			.SE(gen[1948]),

			.SELF(gen[1887]),
			.cell_state(gen[1887])
		); 

/******************* CELL 1888 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1888 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1827]),
			.N(gen[1828]),
			.NE(gen[1829]),

			.O(gen[1887]),
			.E(gen[1889]),

			.SO(gen[1947]),
			.S(gen[1948]),
			.SE(gen[1949]),

			.SELF(gen[1888]),
			.cell_state(gen[1888])
		); 

/******************* CELL 1889 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1889 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1828]),
			.N(gen[1829]),
			.NE(gen[1830]),

			.O(gen[1888]),
			.E(gen[1890]),

			.SO(gen[1948]),
			.S(gen[1949]),
			.SE(gen[1950]),

			.SELF(gen[1889]),
			.cell_state(gen[1889])
		); 

/******************* CELL 1890 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1890 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1829]),
			.N(gen[1830]),
			.NE(gen[1831]),

			.O(gen[1889]),
			.E(gen[1891]),

			.SO(gen[1949]),
			.S(gen[1950]),
			.SE(gen[1951]),

			.SELF(gen[1890]),
			.cell_state(gen[1890])
		); 

/******************* CELL 1891 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1891 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1830]),
			.N(gen[1831]),
			.NE(gen[1832]),

			.O(gen[1890]),
			.E(gen[1892]),

			.SO(gen[1950]),
			.S(gen[1951]),
			.SE(gen[1952]),

			.SELF(gen[1891]),
			.cell_state(gen[1891])
		); 

/******************* CELL 1892 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1892 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1831]),
			.N(gen[1832]),
			.NE(gen[1833]),

			.O(gen[1891]),
			.E(gen[1893]),

			.SO(gen[1951]),
			.S(gen[1952]),
			.SE(gen[1953]),

			.SELF(gen[1892]),
			.cell_state(gen[1892])
		); 

/******************* CELL 1893 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1893 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1832]),
			.N(gen[1833]),
			.NE(gen[1834]),

			.O(gen[1892]),
			.E(gen[1894]),

			.SO(gen[1952]),
			.S(gen[1953]),
			.SE(gen[1954]),

			.SELF(gen[1893]),
			.cell_state(gen[1893])
		); 

/******************* CELL 1894 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1894 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1833]),
			.N(gen[1834]),
			.NE(gen[1835]),

			.O(gen[1893]),
			.E(gen[1895]),

			.SO(gen[1953]),
			.S(gen[1954]),
			.SE(gen[1955]),

			.SELF(gen[1894]),
			.cell_state(gen[1894])
		); 

/******************* CELL 1895 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1895 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1834]),
			.N(gen[1835]),
			.NE(gen[1836]),

			.O(gen[1894]),
			.E(gen[1896]),

			.SO(gen[1954]),
			.S(gen[1955]),
			.SE(gen[1956]),

			.SELF(gen[1895]),
			.cell_state(gen[1895])
		); 

/******************* CELL 1896 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1896 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1835]),
			.N(gen[1836]),
			.NE(gen[1837]),

			.O(gen[1895]),
			.E(gen[1897]),

			.SO(gen[1955]),
			.S(gen[1956]),
			.SE(gen[1957]),

			.SELF(gen[1896]),
			.cell_state(gen[1896])
		); 

/******************* CELL 1897 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1897 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1836]),
			.N(gen[1837]),
			.NE(gen[1838]),

			.O(gen[1896]),
			.E(gen[1898]),

			.SO(gen[1956]),
			.S(gen[1957]),
			.SE(gen[1958]),

			.SELF(gen[1897]),
			.cell_state(gen[1897])
		); 

/******************* CELL 1898 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1898 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1837]),
			.N(gen[1838]),
			.NE(gen[1839]),

			.O(gen[1897]),
			.E(gen[1899]),

			.SO(gen[1957]),
			.S(gen[1958]),
			.SE(gen[1959]),

			.SELF(gen[1898]),
			.cell_state(gen[1898])
		); 

/******************* CELL 1899 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1899 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1838]),
			.N(gen[1839]),
			.NE(gen[1840]),

			.O(gen[1898]),
			.E(gen[1900]),

			.SO(gen[1958]),
			.S(gen[1959]),
			.SE(gen[1960]),

			.SELF(gen[1899]),
			.cell_state(gen[1899])
		); 

/******************* CELL 1900 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1900 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1839]),
			.N(gen[1840]),
			.NE(gen[1841]),

			.O(gen[1899]),
			.E(gen[1901]),

			.SO(gen[1959]),
			.S(gen[1960]),
			.SE(gen[1961]),

			.SELF(gen[1900]),
			.cell_state(gen[1900])
		); 

/******************* CELL 1901 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1901 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1840]),
			.N(gen[1841]),
			.NE(gen[1842]),

			.O(gen[1900]),
			.E(gen[1902]),

			.SO(gen[1960]),
			.S(gen[1961]),
			.SE(gen[1962]),

			.SELF(gen[1901]),
			.cell_state(gen[1901])
		); 

/******************* CELL 1902 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1902 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1841]),
			.N(gen[1842]),
			.NE(gen[1843]),

			.O(gen[1901]),
			.E(gen[1903]),

			.SO(gen[1961]),
			.S(gen[1962]),
			.SE(gen[1963]),

			.SELF(gen[1902]),
			.cell_state(gen[1902])
		); 

/******************* CELL 1903 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1903 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1842]),
			.N(gen[1843]),
			.NE(gen[1844]),

			.O(gen[1902]),
			.E(gen[1904]),

			.SO(gen[1962]),
			.S(gen[1963]),
			.SE(gen[1964]),

			.SELF(gen[1903]),
			.cell_state(gen[1903])
		); 

/******************* CELL 1904 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1904 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1843]),
			.N(gen[1844]),
			.NE(gen[1845]),

			.O(gen[1903]),
			.E(gen[1905]),

			.SO(gen[1963]),
			.S(gen[1964]),
			.SE(gen[1965]),

			.SELF(gen[1904]),
			.cell_state(gen[1904])
		); 

/******************* CELL 1905 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1905 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1844]),
			.N(gen[1845]),
			.NE(gen[1846]),

			.O(gen[1904]),
			.E(gen[1906]),

			.SO(gen[1964]),
			.S(gen[1965]),
			.SE(gen[1966]),

			.SELF(gen[1905]),
			.cell_state(gen[1905])
		); 

/******************* CELL 1906 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1906 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1845]),
			.N(gen[1846]),
			.NE(gen[1847]),

			.O(gen[1905]),
			.E(gen[1907]),

			.SO(gen[1965]),
			.S(gen[1966]),
			.SE(gen[1967]),

			.SELF(gen[1906]),
			.cell_state(gen[1906])
		); 

/******************* CELL 1907 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1907 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1846]),
			.N(gen[1847]),
			.NE(gen[1848]),

			.O(gen[1906]),
			.E(gen[1908]),

			.SO(gen[1966]),
			.S(gen[1967]),
			.SE(gen[1968]),

			.SELF(gen[1907]),
			.cell_state(gen[1907])
		); 

/******************* CELL 1908 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1908 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1847]),
			.N(gen[1848]),
			.NE(gen[1849]),

			.O(gen[1907]),
			.E(gen[1909]),

			.SO(gen[1967]),
			.S(gen[1968]),
			.SE(gen[1969]),

			.SELF(gen[1908]),
			.cell_state(gen[1908])
		); 

/******************* CELL 1909 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1909 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1848]),
			.N(gen[1849]),
			.NE(gen[1850]),

			.O(gen[1908]),
			.E(gen[1910]),

			.SO(gen[1968]),
			.S(gen[1969]),
			.SE(gen[1970]),

			.SELF(gen[1909]),
			.cell_state(gen[1909])
		); 

/******************* CELL 1910 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1910 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1849]),
			.N(gen[1850]),
			.NE(gen[1851]),

			.O(gen[1909]),
			.E(gen[1911]),

			.SO(gen[1969]),
			.S(gen[1970]),
			.SE(gen[1971]),

			.SELF(gen[1910]),
			.cell_state(gen[1910])
		); 

/******************* CELL 1911 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1911 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1850]),
			.N(gen[1851]),
			.NE(gen[1852]),

			.O(gen[1910]),
			.E(gen[1912]),

			.SO(gen[1970]),
			.S(gen[1971]),
			.SE(gen[1972]),

			.SELF(gen[1911]),
			.cell_state(gen[1911])
		); 

/******************* CELL 1912 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1912 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1851]),
			.N(gen[1852]),
			.NE(gen[1853]),

			.O(gen[1911]),
			.E(gen[1913]),

			.SO(gen[1971]),
			.S(gen[1972]),
			.SE(gen[1973]),

			.SELF(gen[1912]),
			.cell_state(gen[1912])
		); 

/******************* CELL 1913 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1913 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1852]),
			.N(gen[1853]),
			.NE(gen[1854]),

			.O(gen[1912]),
			.E(gen[1914]),

			.SO(gen[1972]),
			.S(gen[1973]),
			.SE(gen[1974]),

			.SELF(gen[1913]),
			.cell_state(gen[1913])
		); 

/******************* CELL 1914 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1914 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1853]),
			.N(gen[1854]),
			.NE(gen[1855]),

			.O(gen[1913]),
			.E(gen[1915]),

			.SO(gen[1973]),
			.S(gen[1974]),
			.SE(gen[1975]),

			.SELF(gen[1914]),
			.cell_state(gen[1914])
		); 

/******************* CELL 1915 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1915 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1854]),
			.N(gen[1855]),
			.NE(gen[1856]),

			.O(gen[1914]),
			.E(gen[1916]),

			.SO(gen[1974]),
			.S(gen[1975]),
			.SE(gen[1976]),

			.SELF(gen[1915]),
			.cell_state(gen[1915])
		); 

/******************* CELL 1916 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1916 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1855]),
			.N(gen[1856]),
			.NE(gen[1857]),

			.O(gen[1915]),
			.E(gen[1917]),

			.SO(gen[1975]),
			.S(gen[1976]),
			.SE(gen[1977]),

			.SELF(gen[1916]),
			.cell_state(gen[1916])
		); 

/******************* CELL 1917 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1917 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1856]),
			.N(gen[1857]),
			.NE(gen[1858]),

			.O(gen[1916]),
			.E(gen[1918]),

			.SO(gen[1976]),
			.S(gen[1977]),
			.SE(gen[1978]),

			.SELF(gen[1917]),
			.cell_state(gen[1917])
		); 

/******************* CELL 1918 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1918 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1857]),
			.N(gen[1858]),
			.NE(gen[1859]),

			.O(gen[1917]),
			.E(gen[1919]),

			.SO(gen[1977]),
			.S(gen[1978]),
			.SE(gen[1979]),

			.SELF(gen[1918]),
			.cell_state(gen[1918])
		); 

/******************* CELL 1919 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1919 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1858]),
			.N(gen[1859]),
			.NE(gen[1858]),

			.O(gen[1918]),
			.E(gen[1918]),

			.SO(gen[1978]),
			.S(gen[1979]),
			.SE(gen[1978]),

			.SELF(gen[1919]),
			.cell_state(gen[1919])
		); 

/******************* CELL 1920 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1920 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1861]),
			.N(gen[1860]),
			.NE(gen[1861]),

			.O(gen[1921]),
			.E(gen[1921]),

			.SO(gen[1981]),
			.S(gen[1980]),
			.SE(gen[1981]),

			.SELF(gen[1920]),
			.cell_state(gen[1920])
		); 

/******************* CELL 1921 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1921 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1860]),
			.N(gen[1861]),
			.NE(gen[1862]),

			.O(gen[1920]),
			.E(gen[1922]),

			.SO(gen[1980]),
			.S(gen[1981]),
			.SE(gen[1982]),

			.SELF(gen[1921]),
			.cell_state(gen[1921])
		); 

/******************* CELL 1922 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1922 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1861]),
			.N(gen[1862]),
			.NE(gen[1863]),

			.O(gen[1921]),
			.E(gen[1923]),

			.SO(gen[1981]),
			.S(gen[1982]),
			.SE(gen[1983]),

			.SELF(gen[1922]),
			.cell_state(gen[1922])
		); 

/******************* CELL 1923 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1923 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1862]),
			.N(gen[1863]),
			.NE(gen[1864]),

			.O(gen[1922]),
			.E(gen[1924]),

			.SO(gen[1982]),
			.S(gen[1983]),
			.SE(gen[1984]),

			.SELF(gen[1923]),
			.cell_state(gen[1923])
		); 

/******************* CELL 1924 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1924 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1863]),
			.N(gen[1864]),
			.NE(gen[1865]),

			.O(gen[1923]),
			.E(gen[1925]),

			.SO(gen[1983]),
			.S(gen[1984]),
			.SE(gen[1985]),

			.SELF(gen[1924]),
			.cell_state(gen[1924])
		); 

/******************* CELL 1925 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1925 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1864]),
			.N(gen[1865]),
			.NE(gen[1866]),

			.O(gen[1924]),
			.E(gen[1926]),

			.SO(gen[1984]),
			.S(gen[1985]),
			.SE(gen[1986]),

			.SELF(gen[1925]),
			.cell_state(gen[1925])
		); 

/******************* CELL 1926 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1926 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1865]),
			.N(gen[1866]),
			.NE(gen[1867]),

			.O(gen[1925]),
			.E(gen[1927]),

			.SO(gen[1985]),
			.S(gen[1986]),
			.SE(gen[1987]),

			.SELF(gen[1926]),
			.cell_state(gen[1926])
		); 

/******************* CELL 1927 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1927 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1866]),
			.N(gen[1867]),
			.NE(gen[1868]),

			.O(gen[1926]),
			.E(gen[1928]),

			.SO(gen[1986]),
			.S(gen[1987]),
			.SE(gen[1988]),

			.SELF(gen[1927]),
			.cell_state(gen[1927])
		); 

/******************* CELL 1928 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1928 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1867]),
			.N(gen[1868]),
			.NE(gen[1869]),

			.O(gen[1927]),
			.E(gen[1929]),

			.SO(gen[1987]),
			.S(gen[1988]),
			.SE(gen[1989]),

			.SELF(gen[1928]),
			.cell_state(gen[1928])
		); 

/******************* CELL 1929 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1929 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1868]),
			.N(gen[1869]),
			.NE(gen[1870]),

			.O(gen[1928]),
			.E(gen[1930]),

			.SO(gen[1988]),
			.S(gen[1989]),
			.SE(gen[1990]),

			.SELF(gen[1929]),
			.cell_state(gen[1929])
		); 

/******************* CELL 1930 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1930 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1869]),
			.N(gen[1870]),
			.NE(gen[1871]),

			.O(gen[1929]),
			.E(gen[1931]),

			.SO(gen[1989]),
			.S(gen[1990]),
			.SE(gen[1991]),

			.SELF(gen[1930]),
			.cell_state(gen[1930])
		); 

/******************* CELL 1931 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1931 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1870]),
			.N(gen[1871]),
			.NE(gen[1872]),

			.O(gen[1930]),
			.E(gen[1932]),

			.SO(gen[1990]),
			.S(gen[1991]),
			.SE(gen[1992]),

			.SELF(gen[1931]),
			.cell_state(gen[1931])
		); 

/******************* CELL 1932 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1932 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1871]),
			.N(gen[1872]),
			.NE(gen[1873]),

			.O(gen[1931]),
			.E(gen[1933]),

			.SO(gen[1991]),
			.S(gen[1992]),
			.SE(gen[1993]),

			.SELF(gen[1932]),
			.cell_state(gen[1932])
		); 

/******************* CELL 1933 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1933 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1872]),
			.N(gen[1873]),
			.NE(gen[1874]),

			.O(gen[1932]),
			.E(gen[1934]),

			.SO(gen[1992]),
			.S(gen[1993]),
			.SE(gen[1994]),

			.SELF(gen[1933]),
			.cell_state(gen[1933])
		); 

/******************* CELL 1934 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1934 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1873]),
			.N(gen[1874]),
			.NE(gen[1875]),

			.O(gen[1933]),
			.E(gen[1935]),

			.SO(gen[1993]),
			.S(gen[1994]),
			.SE(gen[1995]),

			.SELF(gen[1934]),
			.cell_state(gen[1934])
		); 

/******************* CELL 1935 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1935 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1874]),
			.N(gen[1875]),
			.NE(gen[1876]),

			.O(gen[1934]),
			.E(gen[1936]),

			.SO(gen[1994]),
			.S(gen[1995]),
			.SE(gen[1996]),

			.SELF(gen[1935]),
			.cell_state(gen[1935])
		); 

/******************* CELL 1936 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1936 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1875]),
			.N(gen[1876]),
			.NE(gen[1877]),

			.O(gen[1935]),
			.E(gen[1937]),

			.SO(gen[1995]),
			.S(gen[1996]),
			.SE(gen[1997]),

			.SELF(gen[1936]),
			.cell_state(gen[1936])
		); 

/******************* CELL 1937 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1937 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1876]),
			.N(gen[1877]),
			.NE(gen[1878]),

			.O(gen[1936]),
			.E(gen[1938]),

			.SO(gen[1996]),
			.S(gen[1997]),
			.SE(gen[1998]),

			.SELF(gen[1937]),
			.cell_state(gen[1937])
		); 

/******************* CELL 1938 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1938 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1877]),
			.N(gen[1878]),
			.NE(gen[1879]),

			.O(gen[1937]),
			.E(gen[1939]),

			.SO(gen[1997]),
			.S(gen[1998]),
			.SE(gen[1999]),

			.SELF(gen[1938]),
			.cell_state(gen[1938])
		); 

/******************* CELL 1939 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1939 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1878]),
			.N(gen[1879]),
			.NE(gen[1880]),

			.O(gen[1938]),
			.E(gen[1940]),

			.SO(gen[1998]),
			.S(gen[1999]),
			.SE(gen[2000]),

			.SELF(gen[1939]),
			.cell_state(gen[1939])
		); 

/******************* CELL 1940 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1940 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1879]),
			.N(gen[1880]),
			.NE(gen[1881]),

			.O(gen[1939]),
			.E(gen[1941]),

			.SO(gen[1999]),
			.S(gen[2000]),
			.SE(gen[2001]),

			.SELF(gen[1940]),
			.cell_state(gen[1940])
		); 

/******************* CELL 1941 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1941 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1880]),
			.N(gen[1881]),
			.NE(gen[1882]),

			.O(gen[1940]),
			.E(gen[1942]),

			.SO(gen[2000]),
			.S(gen[2001]),
			.SE(gen[2002]),

			.SELF(gen[1941]),
			.cell_state(gen[1941])
		); 

/******************* CELL 1942 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1942 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1881]),
			.N(gen[1882]),
			.NE(gen[1883]),

			.O(gen[1941]),
			.E(gen[1943]),

			.SO(gen[2001]),
			.S(gen[2002]),
			.SE(gen[2003]),

			.SELF(gen[1942]),
			.cell_state(gen[1942])
		); 

/******************* CELL 1943 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1943 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1882]),
			.N(gen[1883]),
			.NE(gen[1884]),

			.O(gen[1942]),
			.E(gen[1944]),

			.SO(gen[2002]),
			.S(gen[2003]),
			.SE(gen[2004]),

			.SELF(gen[1943]),
			.cell_state(gen[1943])
		); 

/******************* CELL 1944 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1944 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1883]),
			.N(gen[1884]),
			.NE(gen[1885]),

			.O(gen[1943]),
			.E(gen[1945]),

			.SO(gen[2003]),
			.S(gen[2004]),
			.SE(gen[2005]),

			.SELF(gen[1944]),
			.cell_state(gen[1944])
		); 

/******************* CELL 1945 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1945 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1884]),
			.N(gen[1885]),
			.NE(gen[1886]),

			.O(gen[1944]),
			.E(gen[1946]),

			.SO(gen[2004]),
			.S(gen[2005]),
			.SE(gen[2006]),

			.SELF(gen[1945]),
			.cell_state(gen[1945])
		); 

/******************* CELL 1946 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1946 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1885]),
			.N(gen[1886]),
			.NE(gen[1887]),

			.O(gen[1945]),
			.E(gen[1947]),

			.SO(gen[2005]),
			.S(gen[2006]),
			.SE(gen[2007]),

			.SELF(gen[1946]),
			.cell_state(gen[1946])
		); 

/******************* CELL 1947 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1947 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1886]),
			.N(gen[1887]),
			.NE(gen[1888]),

			.O(gen[1946]),
			.E(gen[1948]),

			.SO(gen[2006]),
			.S(gen[2007]),
			.SE(gen[2008]),

			.SELF(gen[1947]),
			.cell_state(gen[1947])
		); 

/******************* CELL 1948 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1948 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1887]),
			.N(gen[1888]),
			.NE(gen[1889]),

			.O(gen[1947]),
			.E(gen[1949]),

			.SO(gen[2007]),
			.S(gen[2008]),
			.SE(gen[2009]),

			.SELF(gen[1948]),
			.cell_state(gen[1948])
		); 

/******************* CELL 1949 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1949 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1888]),
			.N(gen[1889]),
			.NE(gen[1890]),

			.O(gen[1948]),
			.E(gen[1950]),

			.SO(gen[2008]),
			.S(gen[2009]),
			.SE(gen[2010]),

			.SELF(gen[1949]),
			.cell_state(gen[1949])
		); 

/******************* CELL 1950 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1950 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1889]),
			.N(gen[1890]),
			.NE(gen[1891]),

			.O(gen[1949]),
			.E(gen[1951]),

			.SO(gen[2009]),
			.S(gen[2010]),
			.SE(gen[2011]),

			.SELF(gen[1950]),
			.cell_state(gen[1950])
		); 

/******************* CELL 1951 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1951 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1890]),
			.N(gen[1891]),
			.NE(gen[1892]),

			.O(gen[1950]),
			.E(gen[1952]),

			.SO(gen[2010]),
			.S(gen[2011]),
			.SE(gen[2012]),

			.SELF(gen[1951]),
			.cell_state(gen[1951])
		); 

/******************* CELL 1952 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1952 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1891]),
			.N(gen[1892]),
			.NE(gen[1893]),

			.O(gen[1951]),
			.E(gen[1953]),

			.SO(gen[2011]),
			.S(gen[2012]),
			.SE(gen[2013]),

			.SELF(gen[1952]),
			.cell_state(gen[1952])
		); 

/******************* CELL 1953 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1953 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1892]),
			.N(gen[1893]),
			.NE(gen[1894]),

			.O(gen[1952]),
			.E(gen[1954]),

			.SO(gen[2012]),
			.S(gen[2013]),
			.SE(gen[2014]),

			.SELF(gen[1953]),
			.cell_state(gen[1953])
		); 

/******************* CELL 1954 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1954 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1893]),
			.N(gen[1894]),
			.NE(gen[1895]),

			.O(gen[1953]),
			.E(gen[1955]),

			.SO(gen[2013]),
			.S(gen[2014]),
			.SE(gen[2015]),

			.SELF(gen[1954]),
			.cell_state(gen[1954])
		); 

/******************* CELL 1955 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1955 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1894]),
			.N(gen[1895]),
			.NE(gen[1896]),

			.O(gen[1954]),
			.E(gen[1956]),

			.SO(gen[2014]),
			.S(gen[2015]),
			.SE(gen[2016]),

			.SELF(gen[1955]),
			.cell_state(gen[1955])
		); 

/******************* CELL 1956 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1956 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1895]),
			.N(gen[1896]),
			.NE(gen[1897]),

			.O(gen[1955]),
			.E(gen[1957]),

			.SO(gen[2015]),
			.S(gen[2016]),
			.SE(gen[2017]),

			.SELF(gen[1956]),
			.cell_state(gen[1956])
		); 

/******************* CELL 1957 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1957 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1896]),
			.N(gen[1897]),
			.NE(gen[1898]),

			.O(gen[1956]),
			.E(gen[1958]),

			.SO(gen[2016]),
			.S(gen[2017]),
			.SE(gen[2018]),

			.SELF(gen[1957]),
			.cell_state(gen[1957])
		); 

/******************* CELL 1958 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1958 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1897]),
			.N(gen[1898]),
			.NE(gen[1899]),

			.O(gen[1957]),
			.E(gen[1959]),

			.SO(gen[2017]),
			.S(gen[2018]),
			.SE(gen[2019]),

			.SELF(gen[1958]),
			.cell_state(gen[1958])
		); 

/******************* CELL 1959 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1959 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1898]),
			.N(gen[1899]),
			.NE(gen[1900]),

			.O(gen[1958]),
			.E(gen[1960]),

			.SO(gen[2018]),
			.S(gen[2019]),
			.SE(gen[2020]),

			.SELF(gen[1959]),
			.cell_state(gen[1959])
		); 

/******************* CELL 1960 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1960 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1899]),
			.N(gen[1900]),
			.NE(gen[1901]),

			.O(gen[1959]),
			.E(gen[1961]),

			.SO(gen[2019]),
			.S(gen[2020]),
			.SE(gen[2021]),

			.SELF(gen[1960]),
			.cell_state(gen[1960])
		); 

/******************* CELL 1961 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1961 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1900]),
			.N(gen[1901]),
			.NE(gen[1902]),

			.O(gen[1960]),
			.E(gen[1962]),

			.SO(gen[2020]),
			.S(gen[2021]),
			.SE(gen[2022]),

			.SELF(gen[1961]),
			.cell_state(gen[1961])
		); 

/******************* CELL 1962 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1962 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1901]),
			.N(gen[1902]),
			.NE(gen[1903]),

			.O(gen[1961]),
			.E(gen[1963]),

			.SO(gen[2021]),
			.S(gen[2022]),
			.SE(gen[2023]),

			.SELF(gen[1962]),
			.cell_state(gen[1962])
		); 

/******************* CELL 1963 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1963 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1902]),
			.N(gen[1903]),
			.NE(gen[1904]),

			.O(gen[1962]),
			.E(gen[1964]),

			.SO(gen[2022]),
			.S(gen[2023]),
			.SE(gen[2024]),

			.SELF(gen[1963]),
			.cell_state(gen[1963])
		); 

/******************* CELL 1964 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1964 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1903]),
			.N(gen[1904]),
			.NE(gen[1905]),

			.O(gen[1963]),
			.E(gen[1965]),

			.SO(gen[2023]),
			.S(gen[2024]),
			.SE(gen[2025]),

			.SELF(gen[1964]),
			.cell_state(gen[1964])
		); 

/******************* CELL 1965 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1965 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1904]),
			.N(gen[1905]),
			.NE(gen[1906]),

			.O(gen[1964]),
			.E(gen[1966]),

			.SO(gen[2024]),
			.S(gen[2025]),
			.SE(gen[2026]),

			.SELF(gen[1965]),
			.cell_state(gen[1965])
		); 

/******************* CELL 1966 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1966 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1905]),
			.N(gen[1906]),
			.NE(gen[1907]),

			.O(gen[1965]),
			.E(gen[1967]),

			.SO(gen[2025]),
			.S(gen[2026]),
			.SE(gen[2027]),

			.SELF(gen[1966]),
			.cell_state(gen[1966])
		); 

/******************* CELL 1967 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1967 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1906]),
			.N(gen[1907]),
			.NE(gen[1908]),

			.O(gen[1966]),
			.E(gen[1968]),

			.SO(gen[2026]),
			.S(gen[2027]),
			.SE(gen[2028]),

			.SELF(gen[1967]),
			.cell_state(gen[1967])
		); 

/******************* CELL 1968 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1968 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1907]),
			.N(gen[1908]),
			.NE(gen[1909]),

			.O(gen[1967]),
			.E(gen[1969]),

			.SO(gen[2027]),
			.S(gen[2028]),
			.SE(gen[2029]),

			.SELF(gen[1968]),
			.cell_state(gen[1968])
		); 

/******************* CELL 1969 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1969 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1908]),
			.N(gen[1909]),
			.NE(gen[1910]),

			.O(gen[1968]),
			.E(gen[1970]),

			.SO(gen[2028]),
			.S(gen[2029]),
			.SE(gen[2030]),

			.SELF(gen[1969]),
			.cell_state(gen[1969])
		); 

/******************* CELL 1970 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1970 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1909]),
			.N(gen[1910]),
			.NE(gen[1911]),

			.O(gen[1969]),
			.E(gen[1971]),

			.SO(gen[2029]),
			.S(gen[2030]),
			.SE(gen[2031]),

			.SELF(gen[1970]),
			.cell_state(gen[1970])
		); 

/******************* CELL 1971 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1971 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1910]),
			.N(gen[1911]),
			.NE(gen[1912]),

			.O(gen[1970]),
			.E(gen[1972]),

			.SO(gen[2030]),
			.S(gen[2031]),
			.SE(gen[2032]),

			.SELF(gen[1971]),
			.cell_state(gen[1971])
		); 

/******************* CELL 1972 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1972 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1911]),
			.N(gen[1912]),
			.NE(gen[1913]),

			.O(gen[1971]),
			.E(gen[1973]),

			.SO(gen[2031]),
			.S(gen[2032]),
			.SE(gen[2033]),

			.SELF(gen[1972]),
			.cell_state(gen[1972])
		); 

/******************* CELL 1973 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1973 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1912]),
			.N(gen[1913]),
			.NE(gen[1914]),

			.O(gen[1972]),
			.E(gen[1974]),

			.SO(gen[2032]),
			.S(gen[2033]),
			.SE(gen[2034]),

			.SELF(gen[1973]),
			.cell_state(gen[1973])
		); 

/******************* CELL 1974 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1974 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1913]),
			.N(gen[1914]),
			.NE(gen[1915]),

			.O(gen[1973]),
			.E(gen[1975]),

			.SO(gen[2033]),
			.S(gen[2034]),
			.SE(gen[2035]),

			.SELF(gen[1974]),
			.cell_state(gen[1974])
		); 

/******************* CELL 1975 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1975 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1914]),
			.N(gen[1915]),
			.NE(gen[1916]),

			.O(gen[1974]),
			.E(gen[1976]),

			.SO(gen[2034]),
			.S(gen[2035]),
			.SE(gen[2036]),

			.SELF(gen[1975]),
			.cell_state(gen[1975])
		); 

/******************* CELL 1976 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1976 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1915]),
			.N(gen[1916]),
			.NE(gen[1917]),

			.O(gen[1975]),
			.E(gen[1977]),

			.SO(gen[2035]),
			.S(gen[2036]),
			.SE(gen[2037]),

			.SELF(gen[1976]),
			.cell_state(gen[1976])
		); 

/******************* CELL 1977 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1977 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1916]),
			.N(gen[1917]),
			.NE(gen[1918]),

			.O(gen[1976]),
			.E(gen[1978]),

			.SO(gen[2036]),
			.S(gen[2037]),
			.SE(gen[2038]),

			.SELF(gen[1977]),
			.cell_state(gen[1977])
		); 

/******************* CELL 1978 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1978 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1917]),
			.N(gen[1918]),
			.NE(gen[1919]),

			.O(gen[1977]),
			.E(gen[1979]),

			.SO(gen[2037]),
			.S(gen[2038]),
			.SE(gen[2039]),

			.SELF(gen[1978]),
			.cell_state(gen[1978])
		); 

/******************* CELL 1979 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1979 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1918]),
			.N(gen[1919]),
			.NE(gen[1918]),

			.O(gen[1978]),
			.E(gen[1978]),

			.SO(gen[2038]),
			.S(gen[2039]),
			.SE(gen[2038]),

			.SELF(gen[1979]),
			.cell_state(gen[1979])
		); 

/******************* CELL 1980 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1980 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1921]),
			.N(gen[1920]),
			.NE(gen[1921]),

			.O(gen[1981]),
			.E(gen[1981]),

			.SO(gen[2041]),
			.S(gen[2040]),
			.SE(gen[2041]),

			.SELF(gen[1980]),
			.cell_state(gen[1980])
		); 

/******************* CELL 1981 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1981 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1920]),
			.N(gen[1921]),
			.NE(gen[1922]),

			.O(gen[1980]),
			.E(gen[1982]),

			.SO(gen[2040]),
			.S(gen[2041]),
			.SE(gen[2042]),

			.SELF(gen[1981]),
			.cell_state(gen[1981])
		); 

/******************* CELL 1982 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1982 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1921]),
			.N(gen[1922]),
			.NE(gen[1923]),

			.O(gen[1981]),
			.E(gen[1983]),

			.SO(gen[2041]),
			.S(gen[2042]),
			.SE(gen[2043]),

			.SELF(gen[1982]),
			.cell_state(gen[1982])
		); 

/******************* CELL 1983 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1983 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1922]),
			.N(gen[1923]),
			.NE(gen[1924]),

			.O(gen[1982]),
			.E(gen[1984]),

			.SO(gen[2042]),
			.S(gen[2043]),
			.SE(gen[2044]),

			.SELF(gen[1983]),
			.cell_state(gen[1983])
		); 

/******************* CELL 1984 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1984 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1923]),
			.N(gen[1924]),
			.NE(gen[1925]),

			.O(gen[1983]),
			.E(gen[1985]),

			.SO(gen[2043]),
			.S(gen[2044]),
			.SE(gen[2045]),

			.SELF(gen[1984]),
			.cell_state(gen[1984])
		); 

/******************* CELL 1985 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1985 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1924]),
			.N(gen[1925]),
			.NE(gen[1926]),

			.O(gen[1984]),
			.E(gen[1986]),

			.SO(gen[2044]),
			.S(gen[2045]),
			.SE(gen[2046]),

			.SELF(gen[1985]),
			.cell_state(gen[1985])
		); 

/******************* CELL 1986 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1986 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1925]),
			.N(gen[1926]),
			.NE(gen[1927]),

			.O(gen[1985]),
			.E(gen[1987]),

			.SO(gen[2045]),
			.S(gen[2046]),
			.SE(gen[2047]),

			.SELF(gen[1986]),
			.cell_state(gen[1986])
		); 

/******************* CELL 1987 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1987 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1926]),
			.N(gen[1927]),
			.NE(gen[1928]),

			.O(gen[1986]),
			.E(gen[1988]),

			.SO(gen[2046]),
			.S(gen[2047]),
			.SE(gen[2048]),

			.SELF(gen[1987]),
			.cell_state(gen[1987])
		); 

/******************* CELL 1988 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1988 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1927]),
			.N(gen[1928]),
			.NE(gen[1929]),

			.O(gen[1987]),
			.E(gen[1989]),

			.SO(gen[2047]),
			.S(gen[2048]),
			.SE(gen[2049]),

			.SELF(gen[1988]),
			.cell_state(gen[1988])
		); 

/******************* CELL 1989 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1989 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1928]),
			.N(gen[1929]),
			.NE(gen[1930]),

			.O(gen[1988]),
			.E(gen[1990]),

			.SO(gen[2048]),
			.S(gen[2049]),
			.SE(gen[2050]),

			.SELF(gen[1989]),
			.cell_state(gen[1989])
		); 

/******************* CELL 1990 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1990 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1929]),
			.N(gen[1930]),
			.NE(gen[1931]),

			.O(gen[1989]),
			.E(gen[1991]),

			.SO(gen[2049]),
			.S(gen[2050]),
			.SE(gen[2051]),

			.SELF(gen[1990]),
			.cell_state(gen[1990])
		); 

/******************* CELL 1991 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1991 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1930]),
			.N(gen[1931]),
			.NE(gen[1932]),

			.O(gen[1990]),
			.E(gen[1992]),

			.SO(gen[2050]),
			.S(gen[2051]),
			.SE(gen[2052]),

			.SELF(gen[1991]),
			.cell_state(gen[1991])
		); 

/******************* CELL 1992 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1992 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1931]),
			.N(gen[1932]),
			.NE(gen[1933]),

			.O(gen[1991]),
			.E(gen[1993]),

			.SO(gen[2051]),
			.S(gen[2052]),
			.SE(gen[2053]),

			.SELF(gen[1992]),
			.cell_state(gen[1992])
		); 

/******************* CELL 1993 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1993 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1932]),
			.N(gen[1933]),
			.NE(gen[1934]),

			.O(gen[1992]),
			.E(gen[1994]),

			.SO(gen[2052]),
			.S(gen[2053]),
			.SE(gen[2054]),

			.SELF(gen[1993]),
			.cell_state(gen[1993])
		); 

/******************* CELL 1994 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1994 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1933]),
			.N(gen[1934]),
			.NE(gen[1935]),

			.O(gen[1993]),
			.E(gen[1995]),

			.SO(gen[2053]),
			.S(gen[2054]),
			.SE(gen[2055]),

			.SELF(gen[1994]),
			.cell_state(gen[1994])
		); 

/******************* CELL 1995 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1995 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1934]),
			.N(gen[1935]),
			.NE(gen[1936]),

			.O(gen[1994]),
			.E(gen[1996]),

			.SO(gen[2054]),
			.S(gen[2055]),
			.SE(gen[2056]),

			.SELF(gen[1995]),
			.cell_state(gen[1995])
		); 

/******************* CELL 1996 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1996 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1935]),
			.N(gen[1936]),
			.NE(gen[1937]),

			.O(gen[1995]),
			.E(gen[1997]),

			.SO(gen[2055]),
			.S(gen[2056]),
			.SE(gen[2057]),

			.SELF(gen[1996]),
			.cell_state(gen[1996])
		); 

/******************* CELL 1997 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1997 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1936]),
			.N(gen[1937]),
			.NE(gen[1938]),

			.O(gen[1996]),
			.E(gen[1998]),

			.SO(gen[2056]),
			.S(gen[2057]),
			.SE(gen[2058]),

			.SELF(gen[1997]),
			.cell_state(gen[1997])
		); 

/******************* CELL 1998 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1998 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1937]),
			.N(gen[1938]),
			.NE(gen[1939]),

			.O(gen[1997]),
			.E(gen[1999]),

			.SO(gen[2057]),
			.S(gen[2058]),
			.SE(gen[2059]),

			.SELF(gen[1998]),
			.cell_state(gen[1998])
		); 

/******************* CELL 1999 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell1999 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1938]),
			.N(gen[1939]),
			.NE(gen[1940]),

			.O(gen[1998]),
			.E(gen[2000]),

			.SO(gen[2058]),
			.S(gen[2059]),
			.SE(gen[2060]),

			.SELF(gen[1999]),
			.cell_state(gen[1999])
		); 

/******************* CELL 2000 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2000 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1939]),
			.N(gen[1940]),
			.NE(gen[1941]),

			.O(gen[1999]),
			.E(gen[2001]),

			.SO(gen[2059]),
			.S(gen[2060]),
			.SE(gen[2061]),

			.SELF(gen[2000]),
			.cell_state(gen[2000])
		); 

/******************* CELL 2001 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2001 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1940]),
			.N(gen[1941]),
			.NE(gen[1942]),

			.O(gen[2000]),
			.E(gen[2002]),

			.SO(gen[2060]),
			.S(gen[2061]),
			.SE(gen[2062]),

			.SELF(gen[2001]),
			.cell_state(gen[2001])
		); 

/******************* CELL 2002 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2002 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1941]),
			.N(gen[1942]),
			.NE(gen[1943]),

			.O(gen[2001]),
			.E(gen[2003]),

			.SO(gen[2061]),
			.S(gen[2062]),
			.SE(gen[2063]),

			.SELF(gen[2002]),
			.cell_state(gen[2002])
		); 

/******************* CELL 2003 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2003 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1942]),
			.N(gen[1943]),
			.NE(gen[1944]),

			.O(gen[2002]),
			.E(gen[2004]),

			.SO(gen[2062]),
			.S(gen[2063]),
			.SE(gen[2064]),

			.SELF(gen[2003]),
			.cell_state(gen[2003])
		); 

/******************* CELL 2004 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2004 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1943]),
			.N(gen[1944]),
			.NE(gen[1945]),

			.O(gen[2003]),
			.E(gen[2005]),

			.SO(gen[2063]),
			.S(gen[2064]),
			.SE(gen[2065]),

			.SELF(gen[2004]),
			.cell_state(gen[2004])
		); 

/******************* CELL 2005 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2005 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1944]),
			.N(gen[1945]),
			.NE(gen[1946]),

			.O(gen[2004]),
			.E(gen[2006]),

			.SO(gen[2064]),
			.S(gen[2065]),
			.SE(gen[2066]),

			.SELF(gen[2005]),
			.cell_state(gen[2005])
		); 

/******************* CELL 2006 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2006 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1945]),
			.N(gen[1946]),
			.NE(gen[1947]),

			.O(gen[2005]),
			.E(gen[2007]),

			.SO(gen[2065]),
			.S(gen[2066]),
			.SE(gen[2067]),

			.SELF(gen[2006]),
			.cell_state(gen[2006])
		); 

/******************* CELL 2007 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2007 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1946]),
			.N(gen[1947]),
			.NE(gen[1948]),

			.O(gen[2006]),
			.E(gen[2008]),

			.SO(gen[2066]),
			.S(gen[2067]),
			.SE(gen[2068]),

			.SELF(gen[2007]),
			.cell_state(gen[2007])
		); 

/******************* CELL 2008 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2008 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1947]),
			.N(gen[1948]),
			.NE(gen[1949]),

			.O(gen[2007]),
			.E(gen[2009]),

			.SO(gen[2067]),
			.S(gen[2068]),
			.SE(gen[2069]),

			.SELF(gen[2008]),
			.cell_state(gen[2008])
		); 

/******************* CELL 2009 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2009 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1948]),
			.N(gen[1949]),
			.NE(gen[1950]),

			.O(gen[2008]),
			.E(gen[2010]),

			.SO(gen[2068]),
			.S(gen[2069]),
			.SE(gen[2070]),

			.SELF(gen[2009]),
			.cell_state(gen[2009])
		); 

/******************* CELL 2010 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2010 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1949]),
			.N(gen[1950]),
			.NE(gen[1951]),

			.O(gen[2009]),
			.E(gen[2011]),

			.SO(gen[2069]),
			.S(gen[2070]),
			.SE(gen[2071]),

			.SELF(gen[2010]),
			.cell_state(gen[2010])
		); 

/******************* CELL 2011 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2011 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1950]),
			.N(gen[1951]),
			.NE(gen[1952]),

			.O(gen[2010]),
			.E(gen[2012]),

			.SO(gen[2070]),
			.S(gen[2071]),
			.SE(gen[2072]),

			.SELF(gen[2011]),
			.cell_state(gen[2011])
		); 

/******************* CELL 2012 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2012 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1951]),
			.N(gen[1952]),
			.NE(gen[1953]),

			.O(gen[2011]),
			.E(gen[2013]),

			.SO(gen[2071]),
			.S(gen[2072]),
			.SE(gen[2073]),

			.SELF(gen[2012]),
			.cell_state(gen[2012])
		); 

/******************* CELL 2013 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2013 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1952]),
			.N(gen[1953]),
			.NE(gen[1954]),

			.O(gen[2012]),
			.E(gen[2014]),

			.SO(gen[2072]),
			.S(gen[2073]),
			.SE(gen[2074]),

			.SELF(gen[2013]),
			.cell_state(gen[2013])
		); 

/******************* CELL 2014 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2014 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1953]),
			.N(gen[1954]),
			.NE(gen[1955]),

			.O(gen[2013]),
			.E(gen[2015]),

			.SO(gen[2073]),
			.S(gen[2074]),
			.SE(gen[2075]),

			.SELF(gen[2014]),
			.cell_state(gen[2014])
		); 

/******************* CELL 2015 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2015 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1954]),
			.N(gen[1955]),
			.NE(gen[1956]),

			.O(gen[2014]),
			.E(gen[2016]),

			.SO(gen[2074]),
			.S(gen[2075]),
			.SE(gen[2076]),

			.SELF(gen[2015]),
			.cell_state(gen[2015])
		); 

/******************* CELL 2016 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2016 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1955]),
			.N(gen[1956]),
			.NE(gen[1957]),

			.O(gen[2015]),
			.E(gen[2017]),

			.SO(gen[2075]),
			.S(gen[2076]),
			.SE(gen[2077]),

			.SELF(gen[2016]),
			.cell_state(gen[2016])
		); 

/******************* CELL 2017 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2017 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1956]),
			.N(gen[1957]),
			.NE(gen[1958]),

			.O(gen[2016]),
			.E(gen[2018]),

			.SO(gen[2076]),
			.S(gen[2077]),
			.SE(gen[2078]),

			.SELF(gen[2017]),
			.cell_state(gen[2017])
		); 

/******************* CELL 2018 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2018 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1957]),
			.N(gen[1958]),
			.NE(gen[1959]),

			.O(gen[2017]),
			.E(gen[2019]),

			.SO(gen[2077]),
			.S(gen[2078]),
			.SE(gen[2079]),

			.SELF(gen[2018]),
			.cell_state(gen[2018])
		); 

/******************* CELL 2019 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2019 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1958]),
			.N(gen[1959]),
			.NE(gen[1960]),

			.O(gen[2018]),
			.E(gen[2020]),

			.SO(gen[2078]),
			.S(gen[2079]),
			.SE(gen[2080]),

			.SELF(gen[2019]),
			.cell_state(gen[2019])
		); 

/******************* CELL 2020 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2020 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1959]),
			.N(gen[1960]),
			.NE(gen[1961]),

			.O(gen[2019]),
			.E(gen[2021]),

			.SO(gen[2079]),
			.S(gen[2080]),
			.SE(gen[2081]),

			.SELF(gen[2020]),
			.cell_state(gen[2020])
		); 

/******************* CELL 2021 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2021 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1960]),
			.N(gen[1961]),
			.NE(gen[1962]),

			.O(gen[2020]),
			.E(gen[2022]),

			.SO(gen[2080]),
			.S(gen[2081]),
			.SE(gen[2082]),

			.SELF(gen[2021]),
			.cell_state(gen[2021])
		); 

/******************* CELL 2022 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2022 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1961]),
			.N(gen[1962]),
			.NE(gen[1963]),

			.O(gen[2021]),
			.E(gen[2023]),

			.SO(gen[2081]),
			.S(gen[2082]),
			.SE(gen[2083]),

			.SELF(gen[2022]),
			.cell_state(gen[2022])
		); 

/******************* CELL 2023 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2023 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1962]),
			.N(gen[1963]),
			.NE(gen[1964]),

			.O(gen[2022]),
			.E(gen[2024]),

			.SO(gen[2082]),
			.S(gen[2083]),
			.SE(gen[2084]),

			.SELF(gen[2023]),
			.cell_state(gen[2023])
		); 

/******************* CELL 2024 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2024 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1963]),
			.N(gen[1964]),
			.NE(gen[1965]),

			.O(gen[2023]),
			.E(gen[2025]),

			.SO(gen[2083]),
			.S(gen[2084]),
			.SE(gen[2085]),

			.SELF(gen[2024]),
			.cell_state(gen[2024])
		); 

/******************* CELL 2025 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2025 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1964]),
			.N(gen[1965]),
			.NE(gen[1966]),

			.O(gen[2024]),
			.E(gen[2026]),

			.SO(gen[2084]),
			.S(gen[2085]),
			.SE(gen[2086]),

			.SELF(gen[2025]),
			.cell_state(gen[2025])
		); 

/******************* CELL 2026 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2026 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1965]),
			.N(gen[1966]),
			.NE(gen[1967]),

			.O(gen[2025]),
			.E(gen[2027]),

			.SO(gen[2085]),
			.S(gen[2086]),
			.SE(gen[2087]),

			.SELF(gen[2026]),
			.cell_state(gen[2026])
		); 

/******************* CELL 2027 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2027 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1966]),
			.N(gen[1967]),
			.NE(gen[1968]),

			.O(gen[2026]),
			.E(gen[2028]),

			.SO(gen[2086]),
			.S(gen[2087]),
			.SE(gen[2088]),

			.SELF(gen[2027]),
			.cell_state(gen[2027])
		); 

/******************* CELL 2028 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2028 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1967]),
			.N(gen[1968]),
			.NE(gen[1969]),

			.O(gen[2027]),
			.E(gen[2029]),

			.SO(gen[2087]),
			.S(gen[2088]),
			.SE(gen[2089]),

			.SELF(gen[2028]),
			.cell_state(gen[2028])
		); 

/******************* CELL 2029 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2029 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1968]),
			.N(gen[1969]),
			.NE(gen[1970]),

			.O(gen[2028]),
			.E(gen[2030]),

			.SO(gen[2088]),
			.S(gen[2089]),
			.SE(gen[2090]),

			.SELF(gen[2029]),
			.cell_state(gen[2029])
		); 

/******************* CELL 2030 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2030 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1969]),
			.N(gen[1970]),
			.NE(gen[1971]),

			.O(gen[2029]),
			.E(gen[2031]),

			.SO(gen[2089]),
			.S(gen[2090]),
			.SE(gen[2091]),

			.SELF(gen[2030]),
			.cell_state(gen[2030])
		); 

/******************* CELL 2031 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2031 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1970]),
			.N(gen[1971]),
			.NE(gen[1972]),

			.O(gen[2030]),
			.E(gen[2032]),

			.SO(gen[2090]),
			.S(gen[2091]),
			.SE(gen[2092]),

			.SELF(gen[2031]),
			.cell_state(gen[2031])
		); 

/******************* CELL 2032 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2032 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1971]),
			.N(gen[1972]),
			.NE(gen[1973]),

			.O(gen[2031]),
			.E(gen[2033]),

			.SO(gen[2091]),
			.S(gen[2092]),
			.SE(gen[2093]),

			.SELF(gen[2032]),
			.cell_state(gen[2032])
		); 

/******************* CELL 2033 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2033 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1972]),
			.N(gen[1973]),
			.NE(gen[1974]),

			.O(gen[2032]),
			.E(gen[2034]),

			.SO(gen[2092]),
			.S(gen[2093]),
			.SE(gen[2094]),

			.SELF(gen[2033]),
			.cell_state(gen[2033])
		); 

/******************* CELL 2034 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2034 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1973]),
			.N(gen[1974]),
			.NE(gen[1975]),

			.O(gen[2033]),
			.E(gen[2035]),

			.SO(gen[2093]),
			.S(gen[2094]),
			.SE(gen[2095]),

			.SELF(gen[2034]),
			.cell_state(gen[2034])
		); 

/******************* CELL 2035 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2035 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1974]),
			.N(gen[1975]),
			.NE(gen[1976]),

			.O(gen[2034]),
			.E(gen[2036]),

			.SO(gen[2094]),
			.S(gen[2095]),
			.SE(gen[2096]),

			.SELF(gen[2035]),
			.cell_state(gen[2035])
		); 

/******************* CELL 2036 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2036 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1975]),
			.N(gen[1976]),
			.NE(gen[1977]),

			.O(gen[2035]),
			.E(gen[2037]),

			.SO(gen[2095]),
			.S(gen[2096]),
			.SE(gen[2097]),

			.SELF(gen[2036]),
			.cell_state(gen[2036])
		); 

/******************* CELL 2037 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2037 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1976]),
			.N(gen[1977]),
			.NE(gen[1978]),

			.O(gen[2036]),
			.E(gen[2038]),

			.SO(gen[2096]),
			.S(gen[2097]),
			.SE(gen[2098]),

			.SELF(gen[2037]),
			.cell_state(gen[2037])
		); 

/******************* CELL 2038 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2038 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1977]),
			.N(gen[1978]),
			.NE(gen[1979]),

			.O(gen[2037]),
			.E(gen[2039]),

			.SO(gen[2097]),
			.S(gen[2098]),
			.SE(gen[2099]),

			.SELF(gen[2038]),
			.cell_state(gen[2038])
		); 

/******************* CELL 2039 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2039 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1978]),
			.N(gen[1979]),
			.NE(gen[1978]),

			.O(gen[2038]),
			.E(gen[2038]),

			.SO(gen[2098]),
			.S(gen[2099]),
			.SE(gen[2098]),

			.SELF(gen[2039]),
			.cell_state(gen[2039])
		); 

/******************* CELL 2040 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2040 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1981]),
			.N(gen[1980]),
			.NE(gen[1981]),

			.O(gen[2041]),
			.E(gen[2041]),

			.SO(gen[2101]),
			.S(gen[2100]),
			.SE(gen[2101]),

			.SELF(gen[2040]),
			.cell_state(gen[2040])
		); 

/******************* CELL 2041 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2041 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1980]),
			.N(gen[1981]),
			.NE(gen[1982]),

			.O(gen[2040]),
			.E(gen[2042]),

			.SO(gen[2100]),
			.S(gen[2101]),
			.SE(gen[2102]),

			.SELF(gen[2041]),
			.cell_state(gen[2041])
		); 

/******************* CELL 2042 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2042 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1981]),
			.N(gen[1982]),
			.NE(gen[1983]),

			.O(gen[2041]),
			.E(gen[2043]),

			.SO(gen[2101]),
			.S(gen[2102]),
			.SE(gen[2103]),

			.SELF(gen[2042]),
			.cell_state(gen[2042])
		); 

/******************* CELL 2043 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2043 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1982]),
			.N(gen[1983]),
			.NE(gen[1984]),

			.O(gen[2042]),
			.E(gen[2044]),

			.SO(gen[2102]),
			.S(gen[2103]),
			.SE(gen[2104]),

			.SELF(gen[2043]),
			.cell_state(gen[2043])
		); 

/******************* CELL 2044 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2044 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1983]),
			.N(gen[1984]),
			.NE(gen[1985]),

			.O(gen[2043]),
			.E(gen[2045]),

			.SO(gen[2103]),
			.S(gen[2104]),
			.SE(gen[2105]),

			.SELF(gen[2044]),
			.cell_state(gen[2044])
		); 

/******************* CELL 2045 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2045 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1984]),
			.N(gen[1985]),
			.NE(gen[1986]),

			.O(gen[2044]),
			.E(gen[2046]),

			.SO(gen[2104]),
			.S(gen[2105]),
			.SE(gen[2106]),

			.SELF(gen[2045]),
			.cell_state(gen[2045])
		); 

/******************* CELL 2046 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2046 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1985]),
			.N(gen[1986]),
			.NE(gen[1987]),

			.O(gen[2045]),
			.E(gen[2047]),

			.SO(gen[2105]),
			.S(gen[2106]),
			.SE(gen[2107]),

			.SELF(gen[2046]),
			.cell_state(gen[2046])
		); 

/******************* CELL 2047 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2047 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1986]),
			.N(gen[1987]),
			.NE(gen[1988]),

			.O(gen[2046]),
			.E(gen[2048]),

			.SO(gen[2106]),
			.S(gen[2107]),
			.SE(gen[2108]),

			.SELF(gen[2047]),
			.cell_state(gen[2047])
		); 

/******************* CELL 2048 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2048 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1987]),
			.N(gen[1988]),
			.NE(gen[1989]),

			.O(gen[2047]),
			.E(gen[2049]),

			.SO(gen[2107]),
			.S(gen[2108]),
			.SE(gen[2109]),

			.SELF(gen[2048]),
			.cell_state(gen[2048])
		); 

/******************* CELL 2049 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2049 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1988]),
			.N(gen[1989]),
			.NE(gen[1990]),

			.O(gen[2048]),
			.E(gen[2050]),

			.SO(gen[2108]),
			.S(gen[2109]),
			.SE(gen[2110]),

			.SELF(gen[2049]),
			.cell_state(gen[2049])
		); 

/******************* CELL 2050 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2050 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1989]),
			.N(gen[1990]),
			.NE(gen[1991]),

			.O(gen[2049]),
			.E(gen[2051]),

			.SO(gen[2109]),
			.S(gen[2110]),
			.SE(gen[2111]),

			.SELF(gen[2050]),
			.cell_state(gen[2050])
		); 

/******************* CELL 2051 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2051 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1990]),
			.N(gen[1991]),
			.NE(gen[1992]),

			.O(gen[2050]),
			.E(gen[2052]),

			.SO(gen[2110]),
			.S(gen[2111]),
			.SE(gen[2112]),

			.SELF(gen[2051]),
			.cell_state(gen[2051])
		); 

/******************* CELL 2052 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2052 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1991]),
			.N(gen[1992]),
			.NE(gen[1993]),

			.O(gen[2051]),
			.E(gen[2053]),

			.SO(gen[2111]),
			.S(gen[2112]),
			.SE(gen[2113]),

			.SELF(gen[2052]),
			.cell_state(gen[2052])
		); 

/******************* CELL 2053 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2053 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1992]),
			.N(gen[1993]),
			.NE(gen[1994]),

			.O(gen[2052]),
			.E(gen[2054]),

			.SO(gen[2112]),
			.S(gen[2113]),
			.SE(gen[2114]),

			.SELF(gen[2053]),
			.cell_state(gen[2053])
		); 

/******************* CELL 2054 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2054 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1993]),
			.N(gen[1994]),
			.NE(gen[1995]),

			.O(gen[2053]),
			.E(gen[2055]),

			.SO(gen[2113]),
			.S(gen[2114]),
			.SE(gen[2115]),

			.SELF(gen[2054]),
			.cell_state(gen[2054])
		); 

/******************* CELL 2055 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2055 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1994]),
			.N(gen[1995]),
			.NE(gen[1996]),

			.O(gen[2054]),
			.E(gen[2056]),

			.SO(gen[2114]),
			.S(gen[2115]),
			.SE(gen[2116]),

			.SELF(gen[2055]),
			.cell_state(gen[2055])
		); 

/******************* CELL 2056 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2056 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1995]),
			.N(gen[1996]),
			.NE(gen[1997]),

			.O(gen[2055]),
			.E(gen[2057]),

			.SO(gen[2115]),
			.S(gen[2116]),
			.SE(gen[2117]),

			.SELF(gen[2056]),
			.cell_state(gen[2056])
		); 

/******************* CELL 2057 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2057 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1996]),
			.N(gen[1997]),
			.NE(gen[1998]),

			.O(gen[2056]),
			.E(gen[2058]),

			.SO(gen[2116]),
			.S(gen[2117]),
			.SE(gen[2118]),

			.SELF(gen[2057]),
			.cell_state(gen[2057])
		); 

/******************* CELL 2058 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2058 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1997]),
			.N(gen[1998]),
			.NE(gen[1999]),

			.O(gen[2057]),
			.E(gen[2059]),

			.SO(gen[2117]),
			.S(gen[2118]),
			.SE(gen[2119]),

			.SELF(gen[2058]),
			.cell_state(gen[2058])
		); 

/******************* CELL 2059 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2059 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1998]),
			.N(gen[1999]),
			.NE(gen[2000]),

			.O(gen[2058]),
			.E(gen[2060]),

			.SO(gen[2118]),
			.S(gen[2119]),
			.SE(gen[2120]),

			.SELF(gen[2059]),
			.cell_state(gen[2059])
		); 

/******************* CELL 2060 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2060 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[1999]),
			.N(gen[2000]),
			.NE(gen[2001]),

			.O(gen[2059]),
			.E(gen[2061]),

			.SO(gen[2119]),
			.S(gen[2120]),
			.SE(gen[2121]),

			.SELF(gen[2060]),
			.cell_state(gen[2060])
		); 

/******************* CELL 2061 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2061 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2000]),
			.N(gen[2001]),
			.NE(gen[2002]),

			.O(gen[2060]),
			.E(gen[2062]),

			.SO(gen[2120]),
			.S(gen[2121]),
			.SE(gen[2122]),

			.SELF(gen[2061]),
			.cell_state(gen[2061])
		); 

/******************* CELL 2062 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2062 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2001]),
			.N(gen[2002]),
			.NE(gen[2003]),

			.O(gen[2061]),
			.E(gen[2063]),

			.SO(gen[2121]),
			.S(gen[2122]),
			.SE(gen[2123]),

			.SELF(gen[2062]),
			.cell_state(gen[2062])
		); 

/******************* CELL 2063 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2063 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2002]),
			.N(gen[2003]),
			.NE(gen[2004]),

			.O(gen[2062]),
			.E(gen[2064]),

			.SO(gen[2122]),
			.S(gen[2123]),
			.SE(gen[2124]),

			.SELF(gen[2063]),
			.cell_state(gen[2063])
		); 

/******************* CELL 2064 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2064 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2003]),
			.N(gen[2004]),
			.NE(gen[2005]),

			.O(gen[2063]),
			.E(gen[2065]),

			.SO(gen[2123]),
			.S(gen[2124]),
			.SE(gen[2125]),

			.SELF(gen[2064]),
			.cell_state(gen[2064])
		); 

/******************* CELL 2065 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2065 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2004]),
			.N(gen[2005]),
			.NE(gen[2006]),

			.O(gen[2064]),
			.E(gen[2066]),

			.SO(gen[2124]),
			.S(gen[2125]),
			.SE(gen[2126]),

			.SELF(gen[2065]),
			.cell_state(gen[2065])
		); 

/******************* CELL 2066 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2066 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2005]),
			.N(gen[2006]),
			.NE(gen[2007]),

			.O(gen[2065]),
			.E(gen[2067]),

			.SO(gen[2125]),
			.S(gen[2126]),
			.SE(gen[2127]),

			.SELF(gen[2066]),
			.cell_state(gen[2066])
		); 

/******************* CELL 2067 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2067 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2006]),
			.N(gen[2007]),
			.NE(gen[2008]),

			.O(gen[2066]),
			.E(gen[2068]),

			.SO(gen[2126]),
			.S(gen[2127]),
			.SE(gen[2128]),

			.SELF(gen[2067]),
			.cell_state(gen[2067])
		); 

/******************* CELL 2068 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2068 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2007]),
			.N(gen[2008]),
			.NE(gen[2009]),

			.O(gen[2067]),
			.E(gen[2069]),

			.SO(gen[2127]),
			.S(gen[2128]),
			.SE(gen[2129]),

			.SELF(gen[2068]),
			.cell_state(gen[2068])
		); 

/******************* CELL 2069 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2069 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2008]),
			.N(gen[2009]),
			.NE(gen[2010]),

			.O(gen[2068]),
			.E(gen[2070]),

			.SO(gen[2128]),
			.S(gen[2129]),
			.SE(gen[2130]),

			.SELF(gen[2069]),
			.cell_state(gen[2069])
		); 

/******************* CELL 2070 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2070 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2009]),
			.N(gen[2010]),
			.NE(gen[2011]),

			.O(gen[2069]),
			.E(gen[2071]),

			.SO(gen[2129]),
			.S(gen[2130]),
			.SE(gen[2131]),

			.SELF(gen[2070]),
			.cell_state(gen[2070])
		); 

/******************* CELL 2071 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2071 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2010]),
			.N(gen[2011]),
			.NE(gen[2012]),

			.O(gen[2070]),
			.E(gen[2072]),

			.SO(gen[2130]),
			.S(gen[2131]),
			.SE(gen[2132]),

			.SELF(gen[2071]),
			.cell_state(gen[2071])
		); 

/******************* CELL 2072 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2072 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2011]),
			.N(gen[2012]),
			.NE(gen[2013]),

			.O(gen[2071]),
			.E(gen[2073]),

			.SO(gen[2131]),
			.S(gen[2132]),
			.SE(gen[2133]),

			.SELF(gen[2072]),
			.cell_state(gen[2072])
		); 

/******************* CELL 2073 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2073 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2012]),
			.N(gen[2013]),
			.NE(gen[2014]),

			.O(gen[2072]),
			.E(gen[2074]),

			.SO(gen[2132]),
			.S(gen[2133]),
			.SE(gen[2134]),

			.SELF(gen[2073]),
			.cell_state(gen[2073])
		); 

/******************* CELL 2074 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2074 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2013]),
			.N(gen[2014]),
			.NE(gen[2015]),

			.O(gen[2073]),
			.E(gen[2075]),

			.SO(gen[2133]),
			.S(gen[2134]),
			.SE(gen[2135]),

			.SELF(gen[2074]),
			.cell_state(gen[2074])
		); 

/******************* CELL 2075 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2075 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2014]),
			.N(gen[2015]),
			.NE(gen[2016]),

			.O(gen[2074]),
			.E(gen[2076]),

			.SO(gen[2134]),
			.S(gen[2135]),
			.SE(gen[2136]),

			.SELF(gen[2075]),
			.cell_state(gen[2075])
		); 

/******************* CELL 2076 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2076 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2015]),
			.N(gen[2016]),
			.NE(gen[2017]),

			.O(gen[2075]),
			.E(gen[2077]),

			.SO(gen[2135]),
			.S(gen[2136]),
			.SE(gen[2137]),

			.SELF(gen[2076]),
			.cell_state(gen[2076])
		); 

/******************* CELL 2077 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2077 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2016]),
			.N(gen[2017]),
			.NE(gen[2018]),

			.O(gen[2076]),
			.E(gen[2078]),

			.SO(gen[2136]),
			.S(gen[2137]),
			.SE(gen[2138]),

			.SELF(gen[2077]),
			.cell_state(gen[2077])
		); 

/******************* CELL 2078 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2078 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2017]),
			.N(gen[2018]),
			.NE(gen[2019]),

			.O(gen[2077]),
			.E(gen[2079]),

			.SO(gen[2137]),
			.S(gen[2138]),
			.SE(gen[2139]),

			.SELF(gen[2078]),
			.cell_state(gen[2078])
		); 

/******************* CELL 2079 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2079 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2018]),
			.N(gen[2019]),
			.NE(gen[2020]),

			.O(gen[2078]),
			.E(gen[2080]),

			.SO(gen[2138]),
			.S(gen[2139]),
			.SE(gen[2140]),

			.SELF(gen[2079]),
			.cell_state(gen[2079])
		); 

/******************* CELL 2080 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2080 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2019]),
			.N(gen[2020]),
			.NE(gen[2021]),

			.O(gen[2079]),
			.E(gen[2081]),

			.SO(gen[2139]),
			.S(gen[2140]),
			.SE(gen[2141]),

			.SELF(gen[2080]),
			.cell_state(gen[2080])
		); 

/******************* CELL 2081 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2081 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2020]),
			.N(gen[2021]),
			.NE(gen[2022]),

			.O(gen[2080]),
			.E(gen[2082]),

			.SO(gen[2140]),
			.S(gen[2141]),
			.SE(gen[2142]),

			.SELF(gen[2081]),
			.cell_state(gen[2081])
		); 

/******************* CELL 2082 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2082 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2021]),
			.N(gen[2022]),
			.NE(gen[2023]),

			.O(gen[2081]),
			.E(gen[2083]),

			.SO(gen[2141]),
			.S(gen[2142]),
			.SE(gen[2143]),

			.SELF(gen[2082]),
			.cell_state(gen[2082])
		); 

/******************* CELL 2083 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2083 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2022]),
			.N(gen[2023]),
			.NE(gen[2024]),

			.O(gen[2082]),
			.E(gen[2084]),

			.SO(gen[2142]),
			.S(gen[2143]),
			.SE(gen[2144]),

			.SELF(gen[2083]),
			.cell_state(gen[2083])
		); 

/******************* CELL 2084 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2084 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2023]),
			.N(gen[2024]),
			.NE(gen[2025]),

			.O(gen[2083]),
			.E(gen[2085]),

			.SO(gen[2143]),
			.S(gen[2144]),
			.SE(gen[2145]),

			.SELF(gen[2084]),
			.cell_state(gen[2084])
		); 

/******************* CELL 2085 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2085 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2024]),
			.N(gen[2025]),
			.NE(gen[2026]),

			.O(gen[2084]),
			.E(gen[2086]),

			.SO(gen[2144]),
			.S(gen[2145]),
			.SE(gen[2146]),

			.SELF(gen[2085]),
			.cell_state(gen[2085])
		); 

/******************* CELL 2086 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2086 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2025]),
			.N(gen[2026]),
			.NE(gen[2027]),

			.O(gen[2085]),
			.E(gen[2087]),

			.SO(gen[2145]),
			.S(gen[2146]),
			.SE(gen[2147]),

			.SELF(gen[2086]),
			.cell_state(gen[2086])
		); 

/******************* CELL 2087 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2087 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2026]),
			.N(gen[2027]),
			.NE(gen[2028]),

			.O(gen[2086]),
			.E(gen[2088]),

			.SO(gen[2146]),
			.S(gen[2147]),
			.SE(gen[2148]),

			.SELF(gen[2087]),
			.cell_state(gen[2087])
		); 

/******************* CELL 2088 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2088 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2027]),
			.N(gen[2028]),
			.NE(gen[2029]),

			.O(gen[2087]),
			.E(gen[2089]),

			.SO(gen[2147]),
			.S(gen[2148]),
			.SE(gen[2149]),

			.SELF(gen[2088]),
			.cell_state(gen[2088])
		); 

/******************* CELL 2089 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2089 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2028]),
			.N(gen[2029]),
			.NE(gen[2030]),

			.O(gen[2088]),
			.E(gen[2090]),

			.SO(gen[2148]),
			.S(gen[2149]),
			.SE(gen[2150]),

			.SELF(gen[2089]),
			.cell_state(gen[2089])
		); 

/******************* CELL 2090 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2090 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2029]),
			.N(gen[2030]),
			.NE(gen[2031]),

			.O(gen[2089]),
			.E(gen[2091]),

			.SO(gen[2149]),
			.S(gen[2150]),
			.SE(gen[2151]),

			.SELF(gen[2090]),
			.cell_state(gen[2090])
		); 

/******************* CELL 2091 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2091 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2030]),
			.N(gen[2031]),
			.NE(gen[2032]),

			.O(gen[2090]),
			.E(gen[2092]),

			.SO(gen[2150]),
			.S(gen[2151]),
			.SE(gen[2152]),

			.SELF(gen[2091]),
			.cell_state(gen[2091])
		); 

/******************* CELL 2092 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2092 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2031]),
			.N(gen[2032]),
			.NE(gen[2033]),

			.O(gen[2091]),
			.E(gen[2093]),

			.SO(gen[2151]),
			.S(gen[2152]),
			.SE(gen[2153]),

			.SELF(gen[2092]),
			.cell_state(gen[2092])
		); 

/******************* CELL 2093 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2093 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2032]),
			.N(gen[2033]),
			.NE(gen[2034]),

			.O(gen[2092]),
			.E(gen[2094]),

			.SO(gen[2152]),
			.S(gen[2153]),
			.SE(gen[2154]),

			.SELF(gen[2093]),
			.cell_state(gen[2093])
		); 

/******************* CELL 2094 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2094 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2033]),
			.N(gen[2034]),
			.NE(gen[2035]),

			.O(gen[2093]),
			.E(gen[2095]),

			.SO(gen[2153]),
			.S(gen[2154]),
			.SE(gen[2155]),

			.SELF(gen[2094]),
			.cell_state(gen[2094])
		); 

/******************* CELL 2095 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2095 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2034]),
			.N(gen[2035]),
			.NE(gen[2036]),

			.O(gen[2094]),
			.E(gen[2096]),

			.SO(gen[2154]),
			.S(gen[2155]),
			.SE(gen[2156]),

			.SELF(gen[2095]),
			.cell_state(gen[2095])
		); 

/******************* CELL 2096 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2096 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2035]),
			.N(gen[2036]),
			.NE(gen[2037]),

			.O(gen[2095]),
			.E(gen[2097]),

			.SO(gen[2155]),
			.S(gen[2156]),
			.SE(gen[2157]),

			.SELF(gen[2096]),
			.cell_state(gen[2096])
		); 

/******************* CELL 2097 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2097 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2036]),
			.N(gen[2037]),
			.NE(gen[2038]),

			.O(gen[2096]),
			.E(gen[2098]),

			.SO(gen[2156]),
			.S(gen[2157]),
			.SE(gen[2158]),

			.SELF(gen[2097]),
			.cell_state(gen[2097])
		); 

/******************* CELL 2098 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2098 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2037]),
			.N(gen[2038]),
			.NE(gen[2039]),

			.O(gen[2097]),
			.E(gen[2099]),

			.SO(gen[2157]),
			.S(gen[2158]),
			.SE(gen[2159]),

			.SELF(gen[2098]),
			.cell_state(gen[2098])
		); 

/******************* CELL 2099 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2099 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2038]),
			.N(gen[2039]),
			.NE(gen[2038]),

			.O(gen[2098]),
			.E(gen[2098]),

			.SO(gen[2158]),
			.S(gen[2159]),
			.SE(gen[2158]),

			.SELF(gen[2099]),
			.cell_state(gen[2099])
		); 

/******************* CELL 2100 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2100 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2041]),
			.N(gen[2040]),
			.NE(gen[2041]),

			.O(gen[2101]),
			.E(gen[2101]),

			.SO(gen[2161]),
			.S(gen[2160]),
			.SE(gen[2161]),

			.SELF(gen[2100]),
			.cell_state(gen[2100])
		); 

/******************* CELL 2101 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2101 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2040]),
			.N(gen[2041]),
			.NE(gen[2042]),

			.O(gen[2100]),
			.E(gen[2102]),

			.SO(gen[2160]),
			.S(gen[2161]),
			.SE(gen[2162]),

			.SELF(gen[2101]),
			.cell_state(gen[2101])
		); 

/******************* CELL 2102 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2102 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2041]),
			.N(gen[2042]),
			.NE(gen[2043]),

			.O(gen[2101]),
			.E(gen[2103]),

			.SO(gen[2161]),
			.S(gen[2162]),
			.SE(gen[2163]),

			.SELF(gen[2102]),
			.cell_state(gen[2102])
		); 

/******************* CELL 2103 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2103 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2042]),
			.N(gen[2043]),
			.NE(gen[2044]),

			.O(gen[2102]),
			.E(gen[2104]),

			.SO(gen[2162]),
			.S(gen[2163]),
			.SE(gen[2164]),

			.SELF(gen[2103]),
			.cell_state(gen[2103])
		); 

/******************* CELL 2104 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2104 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2043]),
			.N(gen[2044]),
			.NE(gen[2045]),

			.O(gen[2103]),
			.E(gen[2105]),

			.SO(gen[2163]),
			.S(gen[2164]),
			.SE(gen[2165]),

			.SELF(gen[2104]),
			.cell_state(gen[2104])
		); 

/******************* CELL 2105 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2105 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2044]),
			.N(gen[2045]),
			.NE(gen[2046]),

			.O(gen[2104]),
			.E(gen[2106]),

			.SO(gen[2164]),
			.S(gen[2165]),
			.SE(gen[2166]),

			.SELF(gen[2105]),
			.cell_state(gen[2105])
		); 

/******************* CELL 2106 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2106 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2045]),
			.N(gen[2046]),
			.NE(gen[2047]),

			.O(gen[2105]),
			.E(gen[2107]),

			.SO(gen[2165]),
			.S(gen[2166]),
			.SE(gen[2167]),

			.SELF(gen[2106]),
			.cell_state(gen[2106])
		); 

/******************* CELL 2107 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2107 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2046]),
			.N(gen[2047]),
			.NE(gen[2048]),

			.O(gen[2106]),
			.E(gen[2108]),

			.SO(gen[2166]),
			.S(gen[2167]),
			.SE(gen[2168]),

			.SELF(gen[2107]),
			.cell_state(gen[2107])
		); 

/******************* CELL 2108 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2108 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2047]),
			.N(gen[2048]),
			.NE(gen[2049]),

			.O(gen[2107]),
			.E(gen[2109]),

			.SO(gen[2167]),
			.S(gen[2168]),
			.SE(gen[2169]),

			.SELF(gen[2108]),
			.cell_state(gen[2108])
		); 

/******************* CELL 2109 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2109 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2048]),
			.N(gen[2049]),
			.NE(gen[2050]),

			.O(gen[2108]),
			.E(gen[2110]),

			.SO(gen[2168]),
			.S(gen[2169]),
			.SE(gen[2170]),

			.SELF(gen[2109]),
			.cell_state(gen[2109])
		); 

/******************* CELL 2110 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2110 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2049]),
			.N(gen[2050]),
			.NE(gen[2051]),

			.O(gen[2109]),
			.E(gen[2111]),

			.SO(gen[2169]),
			.S(gen[2170]),
			.SE(gen[2171]),

			.SELF(gen[2110]),
			.cell_state(gen[2110])
		); 

/******************* CELL 2111 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2111 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2050]),
			.N(gen[2051]),
			.NE(gen[2052]),

			.O(gen[2110]),
			.E(gen[2112]),

			.SO(gen[2170]),
			.S(gen[2171]),
			.SE(gen[2172]),

			.SELF(gen[2111]),
			.cell_state(gen[2111])
		); 

/******************* CELL 2112 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2112 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2051]),
			.N(gen[2052]),
			.NE(gen[2053]),

			.O(gen[2111]),
			.E(gen[2113]),

			.SO(gen[2171]),
			.S(gen[2172]),
			.SE(gen[2173]),

			.SELF(gen[2112]),
			.cell_state(gen[2112])
		); 

/******************* CELL 2113 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2113 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2052]),
			.N(gen[2053]),
			.NE(gen[2054]),

			.O(gen[2112]),
			.E(gen[2114]),

			.SO(gen[2172]),
			.S(gen[2173]),
			.SE(gen[2174]),

			.SELF(gen[2113]),
			.cell_state(gen[2113])
		); 

/******************* CELL 2114 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2114 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2053]),
			.N(gen[2054]),
			.NE(gen[2055]),

			.O(gen[2113]),
			.E(gen[2115]),

			.SO(gen[2173]),
			.S(gen[2174]),
			.SE(gen[2175]),

			.SELF(gen[2114]),
			.cell_state(gen[2114])
		); 

/******************* CELL 2115 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2115 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2054]),
			.N(gen[2055]),
			.NE(gen[2056]),

			.O(gen[2114]),
			.E(gen[2116]),

			.SO(gen[2174]),
			.S(gen[2175]),
			.SE(gen[2176]),

			.SELF(gen[2115]),
			.cell_state(gen[2115])
		); 

/******************* CELL 2116 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2116 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2055]),
			.N(gen[2056]),
			.NE(gen[2057]),

			.O(gen[2115]),
			.E(gen[2117]),

			.SO(gen[2175]),
			.S(gen[2176]),
			.SE(gen[2177]),

			.SELF(gen[2116]),
			.cell_state(gen[2116])
		); 

/******************* CELL 2117 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2117 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2056]),
			.N(gen[2057]),
			.NE(gen[2058]),

			.O(gen[2116]),
			.E(gen[2118]),

			.SO(gen[2176]),
			.S(gen[2177]),
			.SE(gen[2178]),

			.SELF(gen[2117]),
			.cell_state(gen[2117])
		); 

/******************* CELL 2118 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2118 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2057]),
			.N(gen[2058]),
			.NE(gen[2059]),

			.O(gen[2117]),
			.E(gen[2119]),

			.SO(gen[2177]),
			.S(gen[2178]),
			.SE(gen[2179]),

			.SELF(gen[2118]),
			.cell_state(gen[2118])
		); 

/******************* CELL 2119 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2119 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2058]),
			.N(gen[2059]),
			.NE(gen[2060]),

			.O(gen[2118]),
			.E(gen[2120]),

			.SO(gen[2178]),
			.S(gen[2179]),
			.SE(gen[2180]),

			.SELF(gen[2119]),
			.cell_state(gen[2119])
		); 

/******************* CELL 2120 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2120 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2059]),
			.N(gen[2060]),
			.NE(gen[2061]),

			.O(gen[2119]),
			.E(gen[2121]),

			.SO(gen[2179]),
			.S(gen[2180]),
			.SE(gen[2181]),

			.SELF(gen[2120]),
			.cell_state(gen[2120])
		); 

/******************* CELL 2121 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2121 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2060]),
			.N(gen[2061]),
			.NE(gen[2062]),

			.O(gen[2120]),
			.E(gen[2122]),

			.SO(gen[2180]),
			.S(gen[2181]),
			.SE(gen[2182]),

			.SELF(gen[2121]),
			.cell_state(gen[2121])
		); 

/******************* CELL 2122 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2122 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2061]),
			.N(gen[2062]),
			.NE(gen[2063]),

			.O(gen[2121]),
			.E(gen[2123]),

			.SO(gen[2181]),
			.S(gen[2182]),
			.SE(gen[2183]),

			.SELF(gen[2122]),
			.cell_state(gen[2122])
		); 

/******************* CELL 2123 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2123 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2062]),
			.N(gen[2063]),
			.NE(gen[2064]),

			.O(gen[2122]),
			.E(gen[2124]),

			.SO(gen[2182]),
			.S(gen[2183]),
			.SE(gen[2184]),

			.SELF(gen[2123]),
			.cell_state(gen[2123])
		); 

/******************* CELL 2124 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2124 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2063]),
			.N(gen[2064]),
			.NE(gen[2065]),

			.O(gen[2123]),
			.E(gen[2125]),

			.SO(gen[2183]),
			.S(gen[2184]),
			.SE(gen[2185]),

			.SELF(gen[2124]),
			.cell_state(gen[2124])
		); 

/******************* CELL 2125 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2125 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2064]),
			.N(gen[2065]),
			.NE(gen[2066]),

			.O(gen[2124]),
			.E(gen[2126]),

			.SO(gen[2184]),
			.S(gen[2185]),
			.SE(gen[2186]),

			.SELF(gen[2125]),
			.cell_state(gen[2125])
		); 

/******************* CELL 2126 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2126 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2065]),
			.N(gen[2066]),
			.NE(gen[2067]),

			.O(gen[2125]),
			.E(gen[2127]),

			.SO(gen[2185]),
			.S(gen[2186]),
			.SE(gen[2187]),

			.SELF(gen[2126]),
			.cell_state(gen[2126])
		); 

/******************* CELL 2127 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2127 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2066]),
			.N(gen[2067]),
			.NE(gen[2068]),

			.O(gen[2126]),
			.E(gen[2128]),

			.SO(gen[2186]),
			.S(gen[2187]),
			.SE(gen[2188]),

			.SELF(gen[2127]),
			.cell_state(gen[2127])
		); 

/******************* CELL 2128 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2128 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2067]),
			.N(gen[2068]),
			.NE(gen[2069]),

			.O(gen[2127]),
			.E(gen[2129]),

			.SO(gen[2187]),
			.S(gen[2188]),
			.SE(gen[2189]),

			.SELF(gen[2128]),
			.cell_state(gen[2128])
		); 

/******************* CELL 2129 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2129 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2068]),
			.N(gen[2069]),
			.NE(gen[2070]),

			.O(gen[2128]),
			.E(gen[2130]),

			.SO(gen[2188]),
			.S(gen[2189]),
			.SE(gen[2190]),

			.SELF(gen[2129]),
			.cell_state(gen[2129])
		); 

/******************* CELL 2130 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2130 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2069]),
			.N(gen[2070]),
			.NE(gen[2071]),

			.O(gen[2129]),
			.E(gen[2131]),

			.SO(gen[2189]),
			.S(gen[2190]),
			.SE(gen[2191]),

			.SELF(gen[2130]),
			.cell_state(gen[2130])
		); 

/******************* CELL 2131 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2131 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2070]),
			.N(gen[2071]),
			.NE(gen[2072]),

			.O(gen[2130]),
			.E(gen[2132]),

			.SO(gen[2190]),
			.S(gen[2191]),
			.SE(gen[2192]),

			.SELF(gen[2131]),
			.cell_state(gen[2131])
		); 

/******************* CELL 2132 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2132 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2071]),
			.N(gen[2072]),
			.NE(gen[2073]),

			.O(gen[2131]),
			.E(gen[2133]),

			.SO(gen[2191]),
			.S(gen[2192]),
			.SE(gen[2193]),

			.SELF(gen[2132]),
			.cell_state(gen[2132])
		); 

/******************* CELL 2133 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2133 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2072]),
			.N(gen[2073]),
			.NE(gen[2074]),

			.O(gen[2132]),
			.E(gen[2134]),

			.SO(gen[2192]),
			.S(gen[2193]),
			.SE(gen[2194]),

			.SELF(gen[2133]),
			.cell_state(gen[2133])
		); 

/******************* CELL 2134 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2134 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2073]),
			.N(gen[2074]),
			.NE(gen[2075]),

			.O(gen[2133]),
			.E(gen[2135]),

			.SO(gen[2193]),
			.S(gen[2194]),
			.SE(gen[2195]),

			.SELF(gen[2134]),
			.cell_state(gen[2134])
		); 

/******************* CELL 2135 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2135 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2074]),
			.N(gen[2075]),
			.NE(gen[2076]),

			.O(gen[2134]),
			.E(gen[2136]),

			.SO(gen[2194]),
			.S(gen[2195]),
			.SE(gen[2196]),

			.SELF(gen[2135]),
			.cell_state(gen[2135])
		); 

/******************* CELL 2136 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2136 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2075]),
			.N(gen[2076]),
			.NE(gen[2077]),

			.O(gen[2135]),
			.E(gen[2137]),

			.SO(gen[2195]),
			.S(gen[2196]),
			.SE(gen[2197]),

			.SELF(gen[2136]),
			.cell_state(gen[2136])
		); 

/******************* CELL 2137 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2137 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2076]),
			.N(gen[2077]),
			.NE(gen[2078]),

			.O(gen[2136]),
			.E(gen[2138]),

			.SO(gen[2196]),
			.S(gen[2197]),
			.SE(gen[2198]),

			.SELF(gen[2137]),
			.cell_state(gen[2137])
		); 

/******************* CELL 2138 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2138 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2077]),
			.N(gen[2078]),
			.NE(gen[2079]),

			.O(gen[2137]),
			.E(gen[2139]),

			.SO(gen[2197]),
			.S(gen[2198]),
			.SE(gen[2199]),

			.SELF(gen[2138]),
			.cell_state(gen[2138])
		); 

/******************* CELL 2139 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2139 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2078]),
			.N(gen[2079]),
			.NE(gen[2080]),

			.O(gen[2138]),
			.E(gen[2140]),

			.SO(gen[2198]),
			.S(gen[2199]),
			.SE(gen[2200]),

			.SELF(gen[2139]),
			.cell_state(gen[2139])
		); 

/******************* CELL 2140 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2140 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2079]),
			.N(gen[2080]),
			.NE(gen[2081]),

			.O(gen[2139]),
			.E(gen[2141]),

			.SO(gen[2199]),
			.S(gen[2200]),
			.SE(gen[2201]),

			.SELF(gen[2140]),
			.cell_state(gen[2140])
		); 

/******************* CELL 2141 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2141 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2080]),
			.N(gen[2081]),
			.NE(gen[2082]),

			.O(gen[2140]),
			.E(gen[2142]),

			.SO(gen[2200]),
			.S(gen[2201]),
			.SE(gen[2202]),

			.SELF(gen[2141]),
			.cell_state(gen[2141])
		); 

/******************* CELL 2142 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2142 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2081]),
			.N(gen[2082]),
			.NE(gen[2083]),

			.O(gen[2141]),
			.E(gen[2143]),

			.SO(gen[2201]),
			.S(gen[2202]),
			.SE(gen[2203]),

			.SELF(gen[2142]),
			.cell_state(gen[2142])
		); 

/******************* CELL 2143 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2143 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2082]),
			.N(gen[2083]),
			.NE(gen[2084]),

			.O(gen[2142]),
			.E(gen[2144]),

			.SO(gen[2202]),
			.S(gen[2203]),
			.SE(gen[2204]),

			.SELF(gen[2143]),
			.cell_state(gen[2143])
		); 

/******************* CELL 2144 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2144 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2083]),
			.N(gen[2084]),
			.NE(gen[2085]),

			.O(gen[2143]),
			.E(gen[2145]),

			.SO(gen[2203]),
			.S(gen[2204]),
			.SE(gen[2205]),

			.SELF(gen[2144]),
			.cell_state(gen[2144])
		); 

/******************* CELL 2145 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2145 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2084]),
			.N(gen[2085]),
			.NE(gen[2086]),

			.O(gen[2144]),
			.E(gen[2146]),

			.SO(gen[2204]),
			.S(gen[2205]),
			.SE(gen[2206]),

			.SELF(gen[2145]),
			.cell_state(gen[2145])
		); 

/******************* CELL 2146 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2146 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2085]),
			.N(gen[2086]),
			.NE(gen[2087]),

			.O(gen[2145]),
			.E(gen[2147]),

			.SO(gen[2205]),
			.S(gen[2206]),
			.SE(gen[2207]),

			.SELF(gen[2146]),
			.cell_state(gen[2146])
		); 

/******************* CELL 2147 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2147 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2086]),
			.N(gen[2087]),
			.NE(gen[2088]),

			.O(gen[2146]),
			.E(gen[2148]),

			.SO(gen[2206]),
			.S(gen[2207]),
			.SE(gen[2208]),

			.SELF(gen[2147]),
			.cell_state(gen[2147])
		); 

/******************* CELL 2148 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2148 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2087]),
			.N(gen[2088]),
			.NE(gen[2089]),

			.O(gen[2147]),
			.E(gen[2149]),

			.SO(gen[2207]),
			.S(gen[2208]),
			.SE(gen[2209]),

			.SELF(gen[2148]),
			.cell_state(gen[2148])
		); 

/******************* CELL 2149 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2149 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2088]),
			.N(gen[2089]),
			.NE(gen[2090]),

			.O(gen[2148]),
			.E(gen[2150]),

			.SO(gen[2208]),
			.S(gen[2209]),
			.SE(gen[2210]),

			.SELF(gen[2149]),
			.cell_state(gen[2149])
		); 

/******************* CELL 2150 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2150 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2089]),
			.N(gen[2090]),
			.NE(gen[2091]),

			.O(gen[2149]),
			.E(gen[2151]),

			.SO(gen[2209]),
			.S(gen[2210]),
			.SE(gen[2211]),

			.SELF(gen[2150]),
			.cell_state(gen[2150])
		); 

/******************* CELL 2151 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2151 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2090]),
			.N(gen[2091]),
			.NE(gen[2092]),

			.O(gen[2150]),
			.E(gen[2152]),

			.SO(gen[2210]),
			.S(gen[2211]),
			.SE(gen[2212]),

			.SELF(gen[2151]),
			.cell_state(gen[2151])
		); 

/******************* CELL 2152 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2152 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2091]),
			.N(gen[2092]),
			.NE(gen[2093]),

			.O(gen[2151]),
			.E(gen[2153]),

			.SO(gen[2211]),
			.S(gen[2212]),
			.SE(gen[2213]),

			.SELF(gen[2152]),
			.cell_state(gen[2152])
		); 

/******************* CELL 2153 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2153 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2092]),
			.N(gen[2093]),
			.NE(gen[2094]),

			.O(gen[2152]),
			.E(gen[2154]),

			.SO(gen[2212]),
			.S(gen[2213]),
			.SE(gen[2214]),

			.SELF(gen[2153]),
			.cell_state(gen[2153])
		); 

/******************* CELL 2154 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2154 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2093]),
			.N(gen[2094]),
			.NE(gen[2095]),

			.O(gen[2153]),
			.E(gen[2155]),

			.SO(gen[2213]),
			.S(gen[2214]),
			.SE(gen[2215]),

			.SELF(gen[2154]),
			.cell_state(gen[2154])
		); 

/******************* CELL 2155 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2155 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2094]),
			.N(gen[2095]),
			.NE(gen[2096]),

			.O(gen[2154]),
			.E(gen[2156]),

			.SO(gen[2214]),
			.S(gen[2215]),
			.SE(gen[2216]),

			.SELF(gen[2155]),
			.cell_state(gen[2155])
		); 

/******************* CELL 2156 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2156 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2095]),
			.N(gen[2096]),
			.NE(gen[2097]),

			.O(gen[2155]),
			.E(gen[2157]),

			.SO(gen[2215]),
			.S(gen[2216]),
			.SE(gen[2217]),

			.SELF(gen[2156]),
			.cell_state(gen[2156])
		); 

/******************* CELL 2157 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2157 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2096]),
			.N(gen[2097]),
			.NE(gen[2098]),

			.O(gen[2156]),
			.E(gen[2158]),

			.SO(gen[2216]),
			.S(gen[2217]),
			.SE(gen[2218]),

			.SELF(gen[2157]),
			.cell_state(gen[2157])
		); 

/******************* CELL 2158 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2158 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2097]),
			.N(gen[2098]),
			.NE(gen[2099]),

			.O(gen[2157]),
			.E(gen[2159]),

			.SO(gen[2217]),
			.S(gen[2218]),
			.SE(gen[2219]),

			.SELF(gen[2158]),
			.cell_state(gen[2158])
		); 

/******************* CELL 2159 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2159 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2098]),
			.N(gen[2099]),
			.NE(gen[2098]),

			.O(gen[2158]),
			.E(gen[2158]),

			.SO(gen[2218]),
			.S(gen[2219]),
			.SE(gen[2218]),

			.SELF(gen[2159]),
			.cell_state(gen[2159])
		); 

/******************* CELL 2160 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2160 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2101]),
			.N(gen[2100]),
			.NE(gen[2101]),

			.O(gen[2161]),
			.E(gen[2161]),

			.SO(gen[2221]),
			.S(gen[2220]),
			.SE(gen[2221]),

			.SELF(gen[2160]),
			.cell_state(gen[2160])
		); 

/******************* CELL 2161 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2161 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2100]),
			.N(gen[2101]),
			.NE(gen[2102]),

			.O(gen[2160]),
			.E(gen[2162]),

			.SO(gen[2220]),
			.S(gen[2221]),
			.SE(gen[2222]),

			.SELF(gen[2161]),
			.cell_state(gen[2161])
		); 

/******************* CELL 2162 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2162 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2101]),
			.N(gen[2102]),
			.NE(gen[2103]),

			.O(gen[2161]),
			.E(gen[2163]),

			.SO(gen[2221]),
			.S(gen[2222]),
			.SE(gen[2223]),

			.SELF(gen[2162]),
			.cell_state(gen[2162])
		); 

/******************* CELL 2163 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2163 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2102]),
			.N(gen[2103]),
			.NE(gen[2104]),

			.O(gen[2162]),
			.E(gen[2164]),

			.SO(gen[2222]),
			.S(gen[2223]),
			.SE(gen[2224]),

			.SELF(gen[2163]),
			.cell_state(gen[2163])
		); 

/******************* CELL 2164 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2164 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2103]),
			.N(gen[2104]),
			.NE(gen[2105]),

			.O(gen[2163]),
			.E(gen[2165]),

			.SO(gen[2223]),
			.S(gen[2224]),
			.SE(gen[2225]),

			.SELF(gen[2164]),
			.cell_state(gen[2164])
		); 

/******************* CELL 2165 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2165 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2104]),
			.N(gen[2105]),
			.NE(gen[2106]),

			.O(gen[2164]),
			.E(gen[2166]),

			.SO(gen[2224]),
			.S(gen[2225]),
			.SE(gen[2226]),

			.SELF(gen[2165]),
			.cell_state(gen[2165])
		); 

/******************* CELL 2166 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2166 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2105]),
			.N(gen[2106]),
			.NE(gen[2107]),

			.O(gen[2165]),
			.E(gen[2167]),

			.SO(gen[2225]),
			.S(gen[2226]),
			.SE(gen[2227]),

			.SELF(gen[2166]),
			.cell_state(gen[2166])
		); 

/******************* CELL 2167 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2167 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2106]),
			.N(gen[2107]),
			.NE(gen[2108]),

			.O(gen[2166]),
			.E(gen[2168]),

			.SO(gen[2226]),
			.S(gen[2227]),
			.SE(gen[2228]),

			.SELF(gen[2167]),
			.cell_state(gen[2167])
		); 

/******************* CELL 2168 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2168 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2107]),
			.N(gen[2108]),
			.NE(gen[2109]),

			.O(gen[2167]),
			.E(gen[2169]),

			.SO(gen[2227]),
			.S(gen[2228]),
			.SE(gen[2229]),

			.SELF(gen[2168]),
			.cell_state(gen[2168])
		); 

/******************* CELL 2169 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2169 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2108]),
			.N(gen[2109]),
			.NE(gen[2110]),

			.O(gen[2168]),
			.E(gen[2170]),

			.SO(gen[2228]),
			.S(gen[2229]),
			.SE(gen[2230]),

			.SELF(gen[2169]),
			.cell_state(gen[2169])
		); 

/******************* CELL 2170 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2170 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2109]),
			.N(gen[2110]),
			.NE(gen[2111]),

			.O(gen[2169]),
			.E(gen[2171]),

			.SO(gen[2229]),
			.S(gen[2230]),
			.SE(gen[2231]),

			.SELF(gen[2170]),
			.cell_state(gen[2170])
		); 

/******************* CELL 2171 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2171 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2110]),
			.N(gen[2111]),
			.NE(gen[2112]),

			.O(gen[2170]),
			.E(gen[2172]),

			.SO(gen[2230]),
			.S(gen[2231]),
			.SE(gen[2232]),

			.SELF(gen[2171]),
			.cell_state(gen[2171])
		); 

/******************* CELL 2172 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2172 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2111]),
			.N(gen[2112]),
			.NE(gen[2113]),

			.O(gen[2171]),
			.E(gen[2173]),

			.SO(gen[2231]),
			.S(gen[2232]),
			.SE(gen[2233]),

			.SELF(gen[2172]),
			.cell_state(gen[2172])
		); 

/******************* CELL 2173 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2173 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2112]),
			.N(gen[2113]),
			.NE(gen[2114]),

			.O(gen[2172]),
			.E(gen[2174]),

			.SO(gen[2232]),
			.S(gen[2233]),
			.SE(gen[2234]),

			.SELF(gen[2173]),
			.cell_state(gen[2173])
		); 

/******************* CELL 2174 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2174 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2113]),
			.N(gen[2114]),
			.NE(gen[2115]),

			.O(gen[2173]),
			.E(gen[2175]),

			.SO(gen[2233]),
			.S(gen[2234]),
			.SE(gen[2235]),

			.SELF(gen[2174]),
			.cell_state(gen[2174])
		); 

/******************* CELL 2175 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2175 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2114]),
			.N(gen[2115]),
			.NE(gen[2116]),

			.O(gen[2174]),
			.E(gen[2176]),

			.SO(gen[2234]),
			.S(gen[2235]),
			.SE(gen[2236]),

			.SELF(gen[2175]),
			.cell_state(gen[2175])
		); 

/******************* CELL 2176 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2176 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2115]),
			.N(gen[2116]),
			.NE(gen[2117]),

			.O(gen[2175]),
			.E(gen[2177]),

			.SO(gen[2235]),
			.S(gen[2236]),
			.SE(gen[2237]),

			.SELF(gen[2176]),
			.cell_state(gen[2176])
		); 

/******************* CELL 2177 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2177 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2116]),
			.N(gen[2117]),
			.NE(gen[2118]),

			.O(gen[2176]),
			.E(gen[2178]),

			.SO(gen[2236]),
			.S(gen[2237]),
			.SE(gen[2238]),

			.SELF(gen[2177]),
			.cell_state(gen[2177])
		); 

/******************* CELL 2178 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2178 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2117]),
			.N(gen[2118]),
			.NE(gen[2119]),

			.O(gen[2177]),
			.E(gen[2179]),

			.SO(gen[2237]),
			.S(gen[2238]),
			.SE(gen[2239]),

			.SELF(gen[2178]),
			.cell_state(gen[2178])
		); 

/******************* CELL 2179 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2179 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2118]),
			.N(gen[2119]),
			.NE(gen[2120]),

			.O(gen[2178]),
			.E(gen[2180]),

			.SO(gen[2238]),
			.S(gen[2239]),
			.SE(gen[2240]),

			.SELF(gen[2179]),
			.cell_state(gen[2179])
		); 

/******************* CELL 2180 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2180 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2119]),
			.N(gen[2120]),
			.NE(gen[2121]),

			.O(gen[2179]),
			.E(gen[2181]),

			.SO(gen[2239]),
			.S(gen[2240]),
			.SE(gen[2241]),

			.SELF(gen[2180]),
			.cell_state(gen[2180])
		); 

/******************* CELL 2181 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2181 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2120]),
			.N(gen[2121]),
			.NE(gen[2122]),

			.O(gen[2180]),
			.E(gen[2182]),

			.SO(gen[2240]),
			.S(gen[2241]),
			.SE(gen[2242]),

			.SELF(gen[2181]),
			.cell_state(gen[2181])
		); 

/******************* CELL 2182 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2182 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2121]),
			.N(gen[2122]),
			.NE(gen[2123]),

			.O(gen[2181]),
			.E(gen[2183]),

			.SO(gen[2241]),
			.S(gen[2242]),
			.SE(gen[2243]),

			.SELF(gen[2182]),
			.cell_state(gen[2182])
		); 

/******************* CELL 2183 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2183 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2122]),
			.N(gen[2123]),
			.NE(gen[2124]),

			.O(gen[2182]),
			.E(gen[2184]),

			.SO(gen[2242]),
			.S(gen[2243]),
			.SE(gen[2244]),

			.SELF(gen[2183]),
			.cell_state(gen[2183])
		); 

/******************* CELL 2184 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2184 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2123]),
			.N(gen[2124]),
			.NE(gen[2125]),

			.O(gen[2183]),
			.E(gen[2185]),

			.SO(gen[2243]),
			.S(gen[2244]),
			.SE(gen[2245]),

			.SELF(gen[2184]),
			.cell_state(gen[2184])
		); 

/******************* CELL 2185 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2185 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2124]),
			.N(gen[2125]),
			.NE(gen[2126]),

			.O(gen[2184]),
			.E(gen[2186]),

			.SO(gen[2244]),
			.S(gen[2245]),
			.SE(gen[2246]),

			.SELF(gen[2185]),
			.cell_state(gen[2185])
		); 

/******************* CELL 2186 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2186 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2125]),
			.N(gen[2126]),
			.NE(gen[2127]),

			.O(gen[2185]),
			.E(gen[2187]),

			.SO(gen[2245]),
			.S(gen[2246]),
			.SE(gen[2247]),

			.SELF(gen[2186]),
			.cell_state(gen[2186])
		); 

/******************* CELL 2187 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2187 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2126]),
			.N(gen[2127]),
			.NE(gen[2128]),

			.O(gen[2186]),
			.E(gen[2188]),

			.SO(gen[2246]),
			.S(gen[2247]),
			.SE(gen[2248]),

			.SELF(gen[2187]),
			.cell_state(gen[2187])
		); 

/******************* CELL 2188 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2188 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2127]),
			.N(gen[2128]),
			.NE(gen[2129]),

			.O(gen[2187]),
			.E(gen[2189]),

			.SO(gen[2247]),
			.S(gen[2248]),
			.SE(gen[2249]),

			.SELF(gen[2188]),
			.cell_state(gen[2188])
		); 

/******************* CELL 2189 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2189 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2128]),
			.N(gen[2129]),
			.NE(gen[2130]),

			.O(gen[2188]),
			.E(gen[2190]),

			.SO(gen[2248]),
			.S(gen[2249]),
			.SE(gen[2250]),

			.SELF(gen[2189]),
			.cell_state(gen[2189])
		); 

/******************* CELL 2190 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2190 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2129]),
			.N(gen[2130]),
			.NE(gen[2131]),

			.O(gen[2189]),
			.E(gen[2191]),

			.SO(gen[2249]),
			.S(gen[2250]),
			.SE(gen[2251]),

			.SELF(gen[2190]),
			.cell_state(gen[2190])
		); 

/******************* CELL 2191 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2191 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2130]),
			.N(gen[2131]),
			.NE(gen[2132]),

			.O(gen[2190]),
			.E(gen[2192]),

			.SO(gen[2250]),
			.S(gen[2251]),
			.SE(gen[2252]),

			.SELF(gen[2191]),
			.cell_state(gen[2191])
		); 

/******************* CELL 2192 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2192 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2131]),
			.N(gen[2132]),
			.NE(gen[2133]),

			.O(gen[2191]),
			.E(gen[2193]),

			.SO(gen[2251]),
			.S(gen[2252]),
			.SE(gen[2253]),

			.SELF(gen[2192]),
			.cell_state(gen[2192])
		); 

/******************* CELL 2193 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2193 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2132]),
			.N(gen[2133]),
			.NE(gen[2134]),

			.O(gen[2192]),
			.E(gen[2194]),

			.SO(gen[2252]),
			.S(gen[2253]),
			.SE(gen[2254]),

			.SELF(gen[2193]),
			.cell_state(gen[2193])
		); 

/******************* CELL 2194 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2194 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2133]),
			.N(gen[2134]),
			.NE(gen[2135]),

			.O(gen[2193]),
			.E(gen[2195]),

			.SO(gen[2253]),
			.S(gen[2254]),
			.SE(gen[2255]),

			.SELF(gen[2194]),
			.cell_state(gen[2194])
		); 

/******************* CELL 2195 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2195 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2134]),
			.N(gen[2135]),
			.NE(gen[2136]),

			.O(gen[2194]),
			.E(gen[2196]),

			.SO(gen[2254]),
			.S(gen[2255]),
			.SE(gen[2256]),

			.SELF(gen[2195]),
			.cell_state(gen[2195])
		); 

/******************* CELL 2196 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2196 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2135]),
			.N(gen[2136]),
			.NE(gen[2137]),

			.O(gen[2195]),
			.E(gen[2197]),

			.SO(gen[2255]),
			.S(gen[2256]),
			.SE(gen[2257]),

			.SELF(gen[2196]),
			.cell_state(gen[2196])
		); 

/******************* CELL 2197 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2197 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2136]),
			.N(gen[2137]),
			.NE(gen[2138]),

			.O(gen[2196]),
			.E(gen[2198]),

			.SO(gen[2256]),
			.S(gen[2257]),
			.SE(gen[2258]),

			.SELF(gen[2197]),
			.cell_state(gen[2197])
		); 

/******************* CELL 2198 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2198 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2137]),
			.N(gen[2138]),
			.NE(gen[2139]),

			.O(gen[2197]),
			.E(gen[2199]),

			.SO(gen[2257]),
			.S(gen[2258]),
			.SE(gen[2259]),

			.SELF(gen[2198]),
			.cell_state(gen[2198])
		); 

/******************* CELL 2199 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2199 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2138]),
			.N(gen[2139]),
			.NE(gen[2140]),

			.O(gen[2198]),
			.E(gen[2200]),

			.SO(gen[2258]),
			.S(gen[2259]),
			.SE(gen[2260]),

			.SELF(gen[2199]),
			.cell_state(gen[2199])
		); 

/******************* CELL 2200 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2200 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2139]),
			.N(gen[2140]),
			.NE(gen[2141]),

			.O(gen[2199]),
			.E(gen[2201]),

			.SO(gen[2259]),
			.S(gen[2260]),
			.SE(gen[2261]),

			.SELF(gen[2200]),
			.cell_state(gen[2200])
		); 

/******************* CELL 2201 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2201 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2140]),
			.N(gen[2141]),
			.NE(gen[2142]),

			.O(gen[2200]),
			.E(gen[2202]),

			.SO(gen[2260]),
			.S(gen[2261]),
			.SE(gen[2262]),

			.SELF(gen[2201]),
			.cell_state(gen[2201])
		); 

/******************* CELL 2202 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2202 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2141]),
			.N(gen[2142]),
			.NE(gen[2143]),

			.O(gen[2201]),
			.E(gen[2203]),

			.SO(gen[2261]),
			.S(gen[2262]),
			.SE(gen[2263]),

			.SELF(gen[2202]),
			.cell_state(gen[2202])
		); 

/******************* CELL 2203 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2203 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2142]),
			.N(gen[2143]),
			.NE(gen[2144]),

			.O(gen[2202]),
			.E(gen[2204]),

			.SO(gen[2262]),
			.S(gen[2263]),
			.SE(gen[2264]),

			.SELF(gen[2203]),
			.cell_state(gen[2203])
		); 

/******************* CELL 2204 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2204 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2143]),
			.N(gen[2144]),
			.NE(gen[2145]),

			.O(gen[2203]),
			.E(gen[2205]),

			.SO(gen[2263]),
			.S(gen[2264]),
			.SE(gen[2265]),

			.SELF(gen[2204]),
			.cell_state(gen[2204])
		); 

/******************* CELL 2205 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2205 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2144]),
			.N(gen[2145]),
			.NE(gen[2146]),

			.O(gen[2204]),
			.E(gen[2206]),

			.SO(gen[2264]),
			.S(gen[2265]),
			.SE(gen[2266]),

			.SELF(gen[2205]),
			.cell_state(gen[2205])
		); 

/******************* CELL 2206 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2206 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2145]),
			.N(gen[2146]),
			.NE(gen[2147]),

			.O(gen[2205]),
			.E(gen[2207]),

			.SO(gen[2265]),
			.S(gen[2266]),
			.SE(gen[2267]),

			.SELF(gen[2206]),
			.cell_state(gen[2206])
		); 

/******************* CELL 2207 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2207 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2146]),
			.N(gen[2147]),
			.NE(gen[2148]),

			.O(gen[2206]),
			.E(gen[2208]),

			.SO(gen[2266]),
			.S(gen[2267]),
			.SE(gen[2268]),

			.SELF(gen[2207]),
			.cell_state(gen[2207])
		); 

/******************* CELL 2208 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2208 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2147]),
			.N(gen[2148]),
			.NE(gen[2149]),

			.O(gen[2207]),
			.E(gen[2209]),

			.SO(gen[2267]),
			.S(gen[2268]),
			.SE(gen[2269]),

			.SELF(gen[2208]),
			.cell_state(gen[2208])
		); 

/******************* CELL 2209 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2209 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2148]),
			.N(gen[2149]),
			.NE(gen[2150]),

			.O(gen[2208]),
			.E(gen[2210]),

			.SO(gen[2268]),
			.S(gen[2269]),
			.SE(gen[2270]),

			.SELF(gen[2209]),
			.cell_state(gen[2209])
		); 

/******************* CELL 2210 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2210 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2149]),
			.N(gen[2150]),
			.NE(gen[2151]),

			.O(gen[2209]),
			.E(gen[2211]),

			.SO(gen[2269]),
			.S(gen[2270]),
			.SE(gen[2271]),

			.SELF(gen[2210]),
			.cell_state(gen[2210])
		); 

/******************* CELL 2211 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2211 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2150]),
			.N(gen[2151]),
			.NE(gen[2152]),

			.O(gen[2210]),
			.E(gen[2212]),

			.SO(gen[2270]),
			.S(gen[2271]),
			.SE(gen[2272]),

			.SELF(gen[2211]),
			.cell_state(gen[2211])
		); 

/******************* CELL 2212 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2212 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2151]),
			.N(gen[2152]),
			.NE(gen[2153]),

			.O(gen[2211]),
			.E(gen[2213]),

			.SO(gen[2271]),
			.S(gen[2272]),
			.SE(gen[2273]),

			.SELF(gen[2212]),
			.cell_state(gen[2212])
		); 

/******************* CELL 2213 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2213 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2152]),
			.N(gen[2153]),
			.NE(gen[2154]),

			.O(gen[2212]),
			.E(gen[2214]),

			.SO(gen[2272]),
			.S(gen[2273]),
			.SE(gen[2274]),

			.SELF(gen[2213]),
			.cell_state(gen[2213])
		); 

/******************* CELL 2214 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2214 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2153]),
			.N(gen[2154]),
			.NE(gen[2155]),

			.O(gen[2213]),
			.E(gen[2215]),

			.SO(gen[2273]),
			.S(gen[2274]),
			.SE(gen[2275]),

			.SELF(gen[2214]),
			.cell_state(gen[2214])
		); 

/******************* CELL 2215 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2215 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2154]),
			.N(gen[2155]),
			.NE(gen[2156]),

			.O(gen[2214]),
			.E(gen[2216]),

			.SO(gen[2274]),
			.S(gen[2275]),
			.SE(gen[2276]),

			.SELF(gen[2215]),
			.cell_state(gen[2215])
		); 

/******************* CELL 2216 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2216 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2155]),
			.N(gen[2156]),
			.NE(gen[2157]),

			.O(gen[2215]),
			.E(gen[2217]),

			.SO(gen[2275]),
			.S(gen[2276]),
			.SE(gen[2277]),

			.SELF(gen[2216]),
			.cell_state(gen[2216])
		); 

/******************* CELL 2217 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2217 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2156]),
			.N(gen[2157]),
			.NE(gen[2158]),

			.O(gen[2216]),
			.E(gen[2218]),

			.SO(gen[2276]),
			.S(gen[2277]),
			.SE(gen[2278]),

			.SELF(gen[2217]),
			.cell_state(gen[2217])
		); 

/******************* CELL 2218 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2218 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2157]),
			.N(gen[2158]),
			.NE(gen[2159]),

			.O(gen[2217]),
			.E(gen[2219]),

			.SO(gen[2277]),
			.S(gen[2278]),
			.SE(gen[2279]),

			.SELF(gen[2218]),
			.cell_state(gen[2218])
		); 

/******************* CELL 2219 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2219 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2158]),
			.N(gen[2159]),
			.NE(gen[2158]),

			.O(gen[2218]),
			.E(gen[2218]),

			.SO(gen[2278]),
			.S(gen[2279]),
			.SE(gen[2278]),

			.SELF(gen[2219]),
			.cell_state(gen[2219])
		); 

/******************* CELL 2220 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2220 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2161]),
			.N(gen[2160]),
			.NE(gen[2161]),

			.O(gen[2221]),
			.E(gen[2221]),

			.SO(gen[2281]),
			.S(gen[2280]),
			.SE(gen[2281]),

			.SELF(gen[2220]),
			.cell_state(gen[2220])
		); 

/******************* CELL 2221 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2221 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2160]),
			.N(gen[2161]),
			.NE(gen[2162]),

			.O(gen[2220]),
			.E(gen[2222]),

			.SO(gen[2280]),
			.S(gen[2281]),
			.SE(gen[2282]),

			.SELF(gen[2221]),
			.cell_state(gen[2221])
		); 

/******************* CELL 2222 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2222 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2161]),
			.N(gen[2162]),
			.NE(gen[2163]),

			.O(gen[2221]),
			.E(gen[2223]),

			.SO(gen[2281]),
			.S(gen[2282]),
			.SE(gen[2283]),

			.SELF(gen[2222]),
			.cell_state(gen[2222])
		); 

/******************* CELL 2223 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2223 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2162]),
			.N(gen[2163]),
			.NE(gen[2164]),

			.O(gen[2222]),
			.E(gen[2224]),

			.SO(gen[2282]),
			.S(gen[2283]),
			.SE(gen[2284]),

			.SELF(gen[2223]),
			.cell_state(gen[2223])
		); 

/******************* CELL 2224 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2224 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2163]),
			.N(gen[2164]),
			.NE(gen[2165]),

			.O(gen[2223]),
			.E(gen[2225]),

			.SO(gen[2283]),
			.S(gen[2284]),
			.SE(gen[2285]),

			.SELF(gen[2224]),
			.cell_state(gen[2224])
		); 

/******************* CELL 2225 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2225 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2164]),
			.N(gen[2165]),
			.NE(gen[2166]),

			.O(gen[2224]),
			.E(gen[2226]),

			.SO(gen[2284]),
			.S(gen[2285]),
			.SE(gen[2286]),

			.SELF(gen[2225]),
			.cell_state(gen[2225])
		); 

/******************* CELL 2226 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2226 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2165]),
			.N(gen[2166]),
			.NE(gen[2167]),

			.O(gen[2225]),
			.E(gen[2227]),

			.SO(gen[2285]),
			.S(gen[2286]),
			.SE(gen[2287]),

			.SELF(gen[2226]),
			.cell_state(gen[2226])
		); 

/******************* CELL 2227 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2227 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2166]),
			.N(gen[2167]),
			.NE(gen[2168]),

			.O(gen[2226]),
			.E(gen[2228]),

			.SO(gen[2286]),
			.S(gen[2287]),
			.SE(gen[2288]),

			.SELF(gen[2227]),
			.cell_state(gen[2227])
		); 

/******************* CELL 2228 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2228 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2167]),
			.N(gen[2168]),
			.NE(gen[2169]),

			.O(gen[2227]),
			.E(gen[2229]),

			.SO(gen[2287]),
			.S(gen[2288]),
			.SE(gen[2289]),

			.SELF(gen[2228]),
			.cell_state(gen[2228])
		); 

/******************* CELL 2229 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2229 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2168]),
			.N(gen[2169]),
			.NE(gen[2170]),

			.O(gen[2228]),
			.E(gen[2230]),

			.SO(gen[2288]),
			.S(gen[2289]),
			.SE(gen[2290]),

			.SELF(gen[2229]),
			.cell_state(gen[2229])
		); 

/******************* CELL 2230 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2230 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2169]),
			.N(gen[2170]),
			.NE(gen[2171]),

			.O(gen[2229]),
			.E(gen[2231]),

			.SO(gen[2289]),
			.S(gen[2290]),
			.SE(gen[2291]),

			.SELF(gen[2230]),
			.cell_state(gen[2230])
		); 

/******************* CELL 2231 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2231 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2170]),
			.N(gen[2171]),
			.NE(gen[2172]),

			.O(gen[2230]),
			.E(gen[2232]),

			.SO(gen[2290]),
			.S(gen[2291]),
			.SE(gen[2292]),

			.SELF(gen[2231]),
			.cell_state(gen[2231])
		); 

/******************* CELL 2232 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2232 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2171]),
			.N(gen[2172]),
			.NE(gen[2173]),

			.O(gen[2231]),
			.E(gen[2233]),

			.SO(gen[2291]),
			.S(gen[2292]),
			.SE(gen[2293]),

			.SELF(gen[2232]),
			.cell_state(gen[2232])
		); 

/******************* CELL 2233 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2233 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2172]),
			.N(gen[2173]),
			.NE(gen[2174]),

			.O(gen[2232]),
			.E(gen[2234]),

			.SO(gen[2292]),
			.S(gen[2293]),
			.SE(gen[2294]),

			.SELF(gen[2233]),
			.cell_state(gen[2233])
		); 

/******************* CELL 2234 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2234 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2173]),
			.N(gen[2174]),
			.NE(gen[2175]),

			.O(gen[2233]),
			.E(gen[2235]),

			.SO(gen[2293]),
			.S(gen[2294]),
			.SE(gen[2295]),

			.SELF(gen[2234]),
			.cell_state(gen[2234])
		); 

/******************* CELL 2235 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2235 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2174]),
			.N(gen[2175]),
			.NE(gen[2176]),

			.O(gen[2234]),
			.E(gen[2236]),

			.SO(gen[2294]),
			.S(gen[2295]),
			.SE(gen[2296]),

			.SELF(gen[2235]),
			.cell_state(gen[2235])
		); 

/******************* CELL 2236 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2236 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2175]),
			.N(gen[2176]),
			.NE(gen[2177]),

			.O(gen[2235]),
			.E(gen[2237]),

			.SO(gen[2295]),
			.S(gen[2296]),
			.SE(gen[2297]),

			.SELF(gen[2236]),
			.cell_state(gen[2236])
		); 

/******************* CELL 2237 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2237 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2176]),
			.N(gen[2177]),
			.NE(gen[2178]),

			.O(gen[2236]),
			.E(gen[2238]),

			.SO(gen[2296]),
			.S(gen[2297]),
			.SE(gen[2298]),

			.SELF(gen[2237]),
			.cell_state(gen[2237])
		); 

/******************* CELL 2238 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2238 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2177]),
			.N(gen[2178]),
			.NE(gen[2179]),

			.O(gen[2237]),
			.E(gen[2239]),

			.SO(gen[2297]),
			.S(gen[2298]),
			.SE(gen[2299]),

			.SELF(gen[2238]),
			.cell_state(gen[2238])
		); 

/******************* CELL 2239 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2239 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2178]),
			.N(gen[2179]),
			.NE(gen[2180]),

			.O(gen[2238]),
			.E(gen[2240]),

			.SO(gen[2298]),
			.S(gen[2299]),
			.SE(gen[2300]),

			.SELF(gen[2239]),
			.cell_state(gen[2239])
		); 

/******************* CELL 2240 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2240 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2179]),
			.N(gen[2180]),
			.NE(gen[2181]),

			.O(gen[2239]),
			.E(gen[2241]),

			.SO(gen[2299]),
			.S(gen[2300]),
			.SE(gen[2301]),

			.SELF(gen[2240]),
			.cell_state(gen[2240])
		); 

/******************* CELL 2241 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2241 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2180]),
			.N(gen[2181]),
			.NE(gen[2182]),

			.O(gen[2240]),
			.E(gen[2242]),

			.SO(gen[2300]),
			.S(gen[2301]),
			.SE(gen[2302]),

			.SELF(gen[2241]),
			.cell_state(gen[2241])
		); 

/******************* CELL 2242 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2242 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2181]),
			.N(gen[2182]),
			.NE(gen[2183]),

			.O(gen[2241]),
			.E(gen[2243]),

			.SO(gen[2301]),
			.S(gen[2302]),
			.SE(gen[2303]),

			.SELF(gen[2242]),
			.cell_state(gen[2242])
		); 

/******************* CELL 2243 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2243 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2182]),
			.N(gen[2183]),
			.NE(gen[2184]),

			.O(gen[2242]),
			.E(gen[2244]),

			.SO(gen[2302]),
			.S(gen[2303]),
			.SE(gen[2304]),

			.SELF(gen[2243]),
			.cell_state(gen[2243])
		); 

/******************* CELL 2244 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2244 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2183]),
			.N(gen[2184]),
			.NE(gen[2185]),

			.O(gen[2243]),
			.E(gen[2245]),

			.SO(gen[2303]),
			.S(gen[2304]),
			.SE(gen[2305]),

			.SELF(gen[2244]),
			.cell_state(gen[2244])
		); 

/******************* CELL 2245 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2245 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2184]),
			.N(gen[2185]),
			.NE(gen[2186]),

			.O(gen[2244]),
			.E(gen[2246]),

			.SO(gen[2304]),
			.S(gen[2305]),
			.SE(gen[2306]),

			.SELF(gen[2245]),
			.cell_state(gen[2245])
		); 

/******************* CELL 2246 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2246 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2185]),
			.N(gen[2186]),
			.NE(gen[2187]),

			.O(gen[2245]),
			.E(gen[2247]),

			.SO(gen[2305]),
			.S(gen[2306]),
			.SE(gen[2307]),

			.SELF(gen[2246]),
			.cell_state(gen[2246])
		); 

/******************* CELL 2247 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2247 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2186]),
			.N(gen[2187]),
			.NE(gen[2188]),

			.O(gen[2246]),
			.E(gen[2248]),

			.SO(gen[2306]),
			.S(gen[2307]),
			.SE(gen[2308]),

			.SELF(gen[2247]),
			.cell_state(gen[2247])
		); 

/******************* CELL 2248 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2248 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2187]),
			.N(gen[2188]),
			.NE(gen[2189]),

			.O(gen[2247]),
			.E(gen[2249]),

			.SO(gen[2307]),
			.S(gen[2308]),
			.SE(gen[2309]),

			.SELF(gen[2248]),
			.cell_state(gen[2248])
		); 

/******************* CELL 2249 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2249 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2188]),
			.N(gen[2189]),
			.NE(gen[2190]),

			.O(gen[2248]),
			.E(gen[2250]),

			.SO(gen[2308]),
			.S(gen[2309]),
			.SE(gen[2310]),

			.SELF(gen[2249]),
			.cell_state(gen[2249])
		); 

/******************* CELL 2250 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2250 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2189]),
			.N(gen[2190]),
			.NE(gen[2191]),

			.O(gen[2249]),
			.E(gen[2251]),

			.SO(gen[2309]),
			.S(gen[2310]),
			.SE(gen[2311]),

			.SELF(gen[2250]),
			.cell_state(gen[2250])
		); 

/******************* CELL 2251 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2251 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2190]),
			.N(gen[2191]),
			.NE(gen[2192]),

			.O(gen[2250]),
			.E(gen[2252]),

			.SO(gen[2310]),
			.S(gen[2311]),
			.SE(gen[2312]),

			.SELF(gen[2251]),
			.cell_state(gen[2251])
		); 

/******************* CELL 2252 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2252 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2191]),
			.N(gen[2192]),
			.NE(gen[2193]),

			.O(gen[2251]),
			.E(gen[2253]),

			.SO(gen[2311]),
			.S(gen[2312]),
			.SE(gen[2313]),

			.SELF(gen[2252]),
			.cell_state(gen[2252])
		); 

/******************* CELL 2253 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2253 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2192]),
			.N(gen[2193]),
			.NE(gen[2194]),

			.O(gen[2252]),
			.E(gen[2254]),

			.SO(gen[2312]),
			.S(gen[2313]),
			.SE(gen[2314]),

			.SELF(gen[2253]),
			.cell_state(gen[2253])
		); 

/******************* CELL 2254 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2254 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2193]),
			.N(gen[2194]),
			.NE(gen[2195]),

			.O(gen[2253]),
			.E(gen[2255]),

			.SO(gen[2313]),
			.S(gen[2314]),
			.SE(gen[2315]),

			.SELF(gen[2254]),
			.cell_state(gen[2254])
		); 

/******************* CELL 2255 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2255 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2194]),
			.N(gen[2195]),
			.NE(gen[2196]),

			.O(gen[2254]),
			.E(gen[2256]),

			.SO(gen[2314]),
			.S(gen[2315]),
			.SE(gen[2316]),

			.SELF(gen[2255]),
			.cell_state(gen[2255])
		); 

/******************* CELL 2256 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2256 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2195]),
			.N(gen[2196]),
			.NE(gen[2197]),

			.O(gen[2255]),
			.E(gen[2257]),

			.SO(gen[2315]),
			.S(gen[2316]),
			.SE(gen[2317]),

			.SELF(gen[2256]),
			.cell_state(gen[2256])
		); 

/******************* CELL 2257 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2257 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2196]),
			.N(gen[2197]),
			.NE(gen[2198]),

			.O(gen[2256]),
			.E(gen[2258]),

			.SO(gen[2316]),
			.S(gen[2317]),
			.SE(gen[2318]),

			.SELF(gen[2257]),
			.cell_state(gen[2257])
		); 

/******************* CELL 2258 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2258 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2197]),
			.N(gen[2198]),
			.NE(gen[2199]),

			.O(gen[2257]),
			.E(gen[2259]),

			.SO(gen[2317]),
			.S(gen[2318]),
			.SE(gen[2319]),

			.SELF(gen[2258]),
			.cell_state(gen[2258])
		); 

/******************* CELL 2259 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2259 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2198]),
			.N(gen[2199]),
			.NE(gen[2200]),

			.O(gen[2258]),
			.E(gen[2260]),

			.SO(gen[2318]),
			.S(gen[2319]),
			.SE(gen[2320]),

			.SELF(gen[2259]),
			.cell_state(gen[2259])
		); 

/******************* CELL 2260 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2260 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2199]),
			.N(gen[2200]),
			.NE(gen[2201]),

			.O(gen[2259]),
			.E(gen[2261]),

			.SO(gen[2319]),
			.S(gen[2320]),
			.SE(gen[2321]),

			.SELF(gen[2260]),
			.cell_state(gen[2260])
		); 

/******************* CELL 2261 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2261 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2200]),
			.N(gen[2201]),
			.NE(gen[2202]),

			.O(gen[2260]),
			.E(gen[2262]),

			.SO(gen[2320]),
			.S(gen[2321]),
			.SE(gen[2322]),

			.SELF(gen[2261]),
			.cell_state(gen[2261])
		); 

/******************* CELL 2262 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2262 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2201]),
			.N(gen[2202]),
			.NE(gen[2203]),

			.O(gen[2261]),
			.E(gen[2263]),

			.SO(gen[2321]),
			.S(gen[2322]),
			.SE(gen[2323]),

			.SELF(gen[2262]),
			.cell_state(gen[2262])
		); 

/******************* CELL 2263 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2263 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2202]),
			.N(gen[2203]),
			.NE(gen[2204]),

			.O(gen[2262]),
			.E(gen[2264]),

			.SO(gen[2322]),
			.S(gen[2323]),
			.SE(gen[2324]),

			.SELF(gen[2263]),
			.cell_state(gen[2263])
		); 

/******************* CELL 2264 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2264 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2203]),
			.N(gen[2204]),
			.NE(gen[2205]),

			.O(gen[2263]),
			.E(gen[2265]),

			.SO(gen[2323]),
			.S(gen[2324]),
			.SE(gen[2325]),

			.SELF(gen[2264]),
			.cell_state(gen[2264])
		); 

/******************* CELL 2265 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2265 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2204]),
			.N(gen[2205]),
			.NE(gen[2206]),

			.O(gen[2264]),
			.E(gen[2266]),

			.SO(gen[2324]),
			.S(gen[2325]),
			.SE(gen[2326]),

			.SELF(gen[2265]),
			.cell_state(gen[2265])
		); 

/******************* CELL 2266 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2266 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2205]),
			.N(gen[2206]),
			.NE(gen[2207]),

			.O(gen[2265]),
			.E(gen[2267]),

			.SO(gen[2325]),
			.S(gen[2326]),
			.SE(gen[2327]),

			.SELF(gen[2266]),
			.cell_state(gen[2266])
		); 

/******************* CELL 2267 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2267 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2206]),
			.N(gen[2207]),
			.NE(gen[2208]),

			.O(gen[2266]),
			.E(gen[2268]),

			.SO(gen[2326]),
			.S(gen[2327]),
			.SE(gen[2328]),

			.SELF(gen[2267]),
			.cell_state(gen[2267])
		); 

/******************* CELL 2268 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2268 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2207]),
			.N(gen[2208]),
			.NE(gen[2209]),

			.O(gen[2267]),
			.E(gen[2269]),

			.SO(gen[2327]),
			.S(gen[2328]),
			.SE(gen[2329]),

			.SELF(gen[2268]),
			.cell_state(gen[2268])
		); 

/******************* CELL 2269 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2269 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2208]),
			.N(gen[2209]),
			.NE(gen[2210]),

			.O(gen[2268]),
			.E(gen[2270]),

			.SO(gen[2328]),
			.S(gen[2329]),
			.SE(gen[2330]),

			.SELF(gen[2269]),
			.cell_state(gen[2269])
		); 

/******************* CELL 2270 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2270 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2209]),
			.N(gen[2210]),
			.NE(gen[2211]),

			.O(gen[2269]),
			.E(gen[2271]),

			.SO(gen[2329]),
			.S(gen[2330]),
			.SE(gen[2331]),

			.SELF(gen[2270]),
			.cell_state(gen[2270])
		); 

/******************* CELL 2271 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2271 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2210]),
			.N(gen[2211]),
			.NE(gen[2212]),

			.O(gen[2270]),
			.E(gen[2272]),

			.SO(gen[2330]),
			.S(gen[2331]),
			.SE(gen[2332]),

			.SELF(gen[2271]),
			.cell_state(gen[2271])
		); 

/******************* CELL 2272 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2272 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2211]),
			.N(gen[2212]),
			.NE(gen[2213]),

			.O(gen[2271]),
			.E(gen[2273]),

			.SO(gen[2331]),
			.S(gen[2332]),
			.SE(gen[2333]),

			.SELF(gen[2272]),
			.cell_state(gen[2272])
		); 

/******************* CELL 2273 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2273 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2212]),
			.N(gen[2213]),
			.NE(gen[2214]),

			.O(gen[2272]),
			.E(gen[2274]),

			.SO(gen[2332]),
			.S(gen[2333]),
			.SE(gen[2334]),

			.SELF(gen[2273]),
			.cell_state(gen[2273])
		); 

/******************* CELL 2274 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2274 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2213]),
			.N(gen[2214]),
			.NE(gen[2215]),

			.O(gen[2273]),
			.E(gen[2275]),

			.SO(gen[2333]),
			.S(gen[2334]),
			.SE(gen[2335]),

			.SELF(gen[2274]),
			.cell_state(gen[2274])
		); 

/******************* CELL 2275 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2275 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2214]),
			.N(gen[2215]),
			.NE(gen[2216]),

			.O(gen[2274]),
			.E(gen[2276]),

			.SO(gen[2334]),
			.S(gen[2335]),
			.SE(gen[2336]),

			.SELF(gen[2275]),
			.cell_state(gen[2275])
		); 

/******************* CELL 2276 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2276 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2215]),
			.N(gen[2216]),
			.NE(gen[2217]),

			.O(gen[2275]),
			.E(gen[2277]),

			.SO(gen[2335]),
			.S(gen[2336]),
			.SE(gen[2337]),

			.SELF(gen[2276]),
			.cell_state(gen[2276])
		); 

/******************* CELL 2277 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2277 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2216]),
			.N(gen[2217]),
			.NE(gen[2218]),

			.O(gen[2276]),
			.E(gen[2278]),

			.SO(gen[2336]),
			.S(gen[2337]),
			.SE(gen[2338]),

			.SELF(gen[2277]),
			.cell_state(gen[2277])
		); 

/******************* CELL 2278 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2278 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2217]),
			.N(gen[2218]),
			.NE(gen[2219]),

			.O(gen[2277]),
			.E(gen[2279]),

			.SO(gen[2337]),
			.S(gen[2338]),
			.SE(gen[2339]),

			.SELF(gen[2278]),
			.cell_state(gen[2278])
		); 

/******************* CELL 2279 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2279 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2218]),
			.N(gen[2219]),
			.NE(gen[2218]),

			.O(gen[2278]),
			.E(gen[2278]),

			.SO(gen[2338]),
			.S(gen[2339]),
			.SE(gen[2338]),

			.SELF(gen[2279]),
			.cell_state(gen[2279])
		); 

/******************* CELL 2280 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2280 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2221]),
			.N(gen[2220]),
			.NE(gen[2221]),

			.O(gen[2281]),
			.E(gen[2281]),

			.SO(gen[2341]),
			.S(gen[2340]),
			.SE(gen[2341]),

			.SELF(gen[2280]),
			.cell_state(gen[2280])
		); 

/******************* CELL 2281 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2281 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2220]),
			.N(gen[2221]),
			.NE(gen[2222]),

			.O(gen[2280]),
			.E(gen[2282]),

			.SO(gen[2340]),
			.S(gen[2341]),
			.SE(gen[2342]),

			.SELF(gen[2281]),
			.cell_state(gen[2281])
		); 

/******************* CELL 2282 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2282 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2221]),
			.N(gen[2222]),
			.NE(gen[2223]),

			.O(gen[2281]),
			.E(gen[2283]),

			.SO(gen[2341]),
			.S(gen[2342]),
			.SE(gen[2343]),

			.SELF(gen[2282]),
			.cell_state(gen[2282])
		); 

/******************* CELL 2283 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2283 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2222]),
			.N(gen[2223]),
			.NE(gen[2224]),

			.O(gen[2282]),
			.E(gen[2284]),

			.SO(gen[2342]),
			.S(gen[2343]),
			.SE(gen[2344]),

			.SELF(gen[2283]),
			.cell_state(gen[2283])
		); 

/******************* CELL 2284 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2284 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2223]),
			.N(gen[2224]),
			.NE(gen[2225]),

			.O(gen[2283]),
			.E(gen[2285]),

			.SO(gen[2343]),
			.S(gen[2344]),
			.SE(gen[2345]),

			.SELF(gen[2284]),
			.cell_state(gen[2284])
		); 

/******************* CELL 2285 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2285 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2224]),
			.N(gen[2225]),
			.NE(gen[2226]),

			.O(gen[2284]),
			.E(gen[2286]),

			.SO(gen[2344]),
			.S(gen[2345]),
			.SE(gen[2346]),

			.SELF(gen[2285]),
			.cell_state(gen[2285])
		); 

/******************* CELL 2286 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2286 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2225]),
			.N(gen[2226]),
			.NE(gen[2227]),

			.O(gen[2285]),
			.E(gen[2287]),

			.SO(gen[2345]),
			.S(gen[2346]),
			.SE(gen[2347]),

			.SELF(gen[2286]),
			.cell_state(gen[2286])
		); 

/******************* CELL 2287 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2287 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2226]),
			.N(gen[2227]),
			.NE(gen[2228]),

			.O(gen[2286]),
			.E(gen[2288]),

			.SO(gen[2346]),
			.S(gen[2347]),
			.SE(gen[2348]),

			.SELF(gen[2287]),
			.cell_state(gen[2287])
		); 

/******************* CELL 2288 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2288 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2227]),
			.N(gen[2228]),
			.NE(gen[2229]),

			.O(gen[2287]),
			.E(gen[2289]),

			.SO(gen[2347]),
			.S(gen[2348]),
			.SE(gen[2349]),

			.SELF(gen[2288]),
			.cell_state(gen[2288])
		); 

/******************* CELL 2289 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2289 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2228]),
			.N(gen[2229]),
			.NE(gen[2230]),

			.O(gen[2288]),
			.E(gen[2290]),

			.SO(gen[2348]),
			.S(gen[2349]),
			.SE(gen[2350]),

			.SELF(gen[2289]),
			.cell_state(gen[2289])
		); 

/******************* CELL 2290 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2290 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2229]),
			.N(gen[2230]),
			.NE(gen[2231]),

			.O(gen[2289]),
			.E(gen[2291]),

			.SO(gen[2349]),
			.S(gen[2350]),
			.SE(gen[2351]),

			.SELF(gen[2290]),
			.cell_state(gen[2290])
		); 

/******************* CELL 2291 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2291 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2230]),
			.N(gen[2231]),
			.NE(gen[2232]),

			.O(gen[2290]),
			.E(gen[2292]),

			.SO(gen[2350]),
			.S(gen[2351]),
			.SE(gen[2352]),

			.SELF(gen[2291]),
			.cell_state(gen[2291])
		); 

/******************* CELL 2292 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2292 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2231]),
			.N(gen[2232]),
			.NE(gen[2233]),

			.O(gen[2291]),
			.E(gen[2293]),

			.SO(gen[2351]),
			.S(gen[2352]),
			.SE(gen[2353]),

			.SELF(gen[2292]),
			.cell_state(gen[2292])
		); 

/******************* CELL 2293 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2293 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2232]),
			.N(gen[2233]),
			.NE(gen[2234]),

			.O(gen[2292]),
			.E(gen[2294]),

			.SO(gen[2352]),
			.S(gen[2353]),
			.SE(gen[2354]),

			.SELF(gen[2293]),
			.cell_state(gen[2293])
		); 

/******************* CELL 2294 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2294 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2233]),
			.N(gen[2234]),
			.NE(gen[2235]),

			.O(gen[2293]),
			.E(gen[2295]),

			.SO(gen[2353]),
			.S(gen[2354]),
			.SE(gen[2355]),

			.SELF(gen[2294]),
			.cell_state(gen[2294])
		); 

/******************* CELL 2295 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2295 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2234]),
			.N(gen[2235]),
			.NE(gen[2236]),

			.O(gen[2294]),
			.E(gen[2296]),

			.SO(gen[2354]),
			.S(gen[2355]),
			.SE(gen[2356]),

			.SELF(gen[2295]),
			.cell_state(gen[2295])
		); 

/******************* CELL 2296 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2296 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2235]),
			.N(gen[2236]),
			.NE(gen[2237]),

			.O(gen[2295]),
			.E(gen[2297]),

			.SO(gen[2355]),
			.S(gen[2356]),
			.SE(gen[2357]),

			.SELF(gen[2296]),
			.cell_state(gen[2296])
		); 

/******************* CELL 2297 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2297 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2236]),
			.N(gen[2237]),
			.NE(gen[2238]),

			.O(gen[2296]),
			.E(gen[2298]),

			.SO(gen[2356]),
			.S(gen[2357]),
			.SE(gen[2358]),

			.SELF(gen[2297]),
			.cell_state(gen[2297])
		); 

/******************* CELL 2298 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2298 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2237]),
			.N(gen[2238]),
			.NE(gen[2239]),

			.O(gen[2297]),
			.E(gen[2299]),

			.SO(gen[2357]),
			.S(gen[2358]),
			.SE(gen[2359]),

			.SELF(gen[2298]),
			.cell_state(gen[2298])
		); 

/******************* CELL 2299 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2299 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2238]),
			.N(gen[2239]),
			.NE(gen[2240]),

			.O(gen[2298]),
			.E(gen[2300]),

			.SO(gen[2358]),
			.S(gen[2359]),
			.SE(gen[2360]),

			.SELF(gen[2299]),
			.cell_state(gen[2299])
		); 

/******************* CELL 2300 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2300 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2239]),
			.N(gen[2240]),
			.NE(gen[2241]),

			.O(gen[2299]),
			.E(gen[2301]),

			.SO(gen[2359]),
			.S(gen[2360]),
			.SE(gen[2361]),

			.SELF(gen[2300]),
			.cell_state(gen[2300])
		); 

/******************* CELL 2301 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2301 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2240]),
			.N(gen[2241]),
			.NE(gen[2242]),

			.O(gen[2300]),
			.E(gen[2302]),

			.SO(gen[2360]),
			.S(gen[2361]),
			.SE(gen[2362]),

			.SELF(gen[2301]),
			.cell_state(gen[2301])
		); 

/******************* CELL 2302 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2302 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2241]),
			.N(gen[2242]),
			.NE(gen[2243]),

			.O(gen[2301]),
			.E(gen[2303]),

			.SO(gen[2361]),
			.S(gen[2362]),
			.SE(gen[2363]),

			.SELF(gen[2302]),
			.cell_state(gen[2302])
		); 

/******************* CELL 2303 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2303 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2242]),
			.N(gen[2243]),
			.NE(gen[2244]),

			.O(gen[2302]),
			.E(gen[2304]),

			.SO(gen[2362]),
			.S(gen[2363]),
			.SE(gen[2364]),

			.SELF(gen[2303]),
			.cell_state(gen[2303])
		); 

/******************* CELL 2304 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2304 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2243]),
			.N(gen[2244]),
			.NE(gen[2245]),

			.O(gen[2303]),
			.E(gen[2305]),

			.SO(gen[2363]),
			.S(gen[2364]),
			.SE(gen[2365]),

			.SELF(gen[2304]),
			.cell_state(gen[2304])
		); 

/******************* CELL 2305 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2305 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2244]),
			.N(gen[2245]),
			.NE(gen[2246]),

			.O(gen[2304]),
			.E(gen[2306]),

			.SO(gen[2364]),
			.S(gen[2365]),
			.SE(gen[2366]),

			.SELF(gen[2305]),
			.cell_state(gen[2305])
		); 

/******************* CELL 2306 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2306 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2245]),
			.N(gen[2246]),
			.NE(gen[2247]),

			.O(gen[2305]),
			.E(gen[2307]),

			.SO(gen[2365]),
			.S(gen[2366]),
			.SE(gen[2367]),

			.SELF(gen[2306]),
			.cell_state(gen[2306])
		); 

/******************* CELL 2307 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2307 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2246]),
			.N(gen[2247]),
			.NE(gen[2248]),

			.O(gen[2306]),
			.E(gen[2308]),

			.SO(gen[2366]),
			.S(gen[2367]),
			.SE(gen[2368]),

			.SELF(gen[2307]),
			.cell_state(gen[2307])
		); 

/******************* CELL 2308 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2308 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2247]),
			.N(gen[2248]),
			.NE(gen[2249]),

			.O(gen[2307]),
			.E(gen[2309]),

			.SO(gen[2367]),
			.S(gen[2368]),
			.SE(gen[2369]),

			.SELF(gen[2308]),
			.cell_state(gen[2308])
		); 

/******************* CELL 2309 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2309 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2248]),
			.N(gen[2249]),
			.NE(gen[2250]),

			.O(gen[2308]),
			.E(gen[2310]),

			.SO(gen[2368]),
			.S(gen[2369]),
			.SE(gen[2370]),

			.SELF(gen[2309]),
			.cell_state(gen[2309])
		); 

/******************* CELL 2310 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2310 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2249]),
			.N(gen[2250]),
			.NE(gen[2251]),

			.O(gen[2309]),
			.E(gen[2311]),

			.SO(gen[2369]),
			.S(gen[2370]),
			.SE(gen[2371]),

			.SELF(gen[2310]),
			.cell_state(gen[2310])
		); 

/******************* CELL 2311 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2311 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2250]),
			.N(gen[2251]),
			.NE(gen[2252]),

			.O(gen[2310]),
			.E(gen[2312]),

			.SO(gen[2370]),
			.S(gen[2371]),
			.SE(gen[2372]),

			.SELF(gen[2311]),
			.cell_state(gen[2311])
		); 

/******************* CELL 2312 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2312 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2251]),
			.N(gen[2252]),
			.NE(gen[2253]),

			.O(gen[2311]),
			.E(gen[2313]),

			.SO(gen[2371]),
			.S(gen[2372]),
			.SE(gen[2373]),

			.SELF(gen[2312]),
			.cell_state(gen[2312])
		); 

/******************* CELL 2313 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2313 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2252]),
			.N(gen[2253]),
			.NE(gen[2254]),

			.O(gen[2312]),
			.E(gen[2314]),

			.SO(gen[2372]),
			.S(gen[2373]),
			.SE(gen[2374]),

			.SELF(gen[2313]),
			.cell_state(gen[2313])
		); 

/******************* CELL 2314 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2314 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2253]),
			.N(gen[2254]),
			.NE(gen[2255]),

			.O(gen[2313]),
			.E(gen[2315]),

			.SO(gen[2373]),
			.S(gen[2374]),
			.SE(gen[2375]),

			.SELF(gen[2314]),
			.cell_state(gen[2314])
		); 

/******************* CELL 2315 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2315 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2254]),
			.N(gen[2255]),
			.NE(gen[2256]),

			.O(gen[2314]),
			.E(gen[2316]),

			.SO(gen[2374]),
			.S(gen[2375]),
			.SE(gen[2376]),

			.SELF(gen[2315]),
			.cell_state(gen[2315])
		); 

/******************* CELL 2316 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2316 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2255]),
			.N(gen[2256]),
			.NE(gen[2257]),

			.O(gen[2315]),
			.E(gen[2317]),

			.SO(gen[2375]),
			.S(gen[2376]),
			.SE(gen[2377]),

			.SELF(gen[2316]),
			.cell_state(gen[2316])
		); 

/******************* CELL 2317 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2317 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2256]),
			.N(gen[2257]),
			.NE(gen[2258]),

			.O(gen[2316]),
			.E(gen[2318]),

			.SO(gen[2376]),
			.S(gen[2377]),
			.SE(gen[2378]),

			.SELF(gen[2317]),
			.cell_state(gen[2317])
		); 

/******************* CELL 2318 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2318 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2257]),
			.N(gen[2258]),
			.NE(gen[2259]),

			.O(gen[2317]),
			.E(gen[2319]),

			.SO(gen[2377]),
			.S(gen[2378]),
			.SE(gen[2379]),

			.SELF(gen[2318]),
			.cell_state(gen[2318])
		); 

/******************* CELL 2319 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2319 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2258]),
			.N(gen[2259]),
			.NE(gen[2260]),

			.O(gen[2318]),
			.E(gen[2320]),

			.SO(gen[2378]),
			.S(gen[2379]),
			.SE(gen[2380]),

			.SELF(gen[2319]),
			.cell_state(gen[2319])
		); 

/******************* CELL 2320 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2320 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2259]),
			.N(gen[2260]),
			.NE(gen[2261]),

			.O(gen[2319]),
			.E(gen[2321]),

			.SO(gen[2379]),
			.S(gen[2380]),
			.SE(gen[2381]),

			.SELF(gen[2320]),
			.cell_state(gen[2320])
		); 

/******************* CELL 2321 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2321 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2260]),
			.N(gen[2261]),
			.NE(gen[2262]),

			.O(gen[2320]),
			.E(gen[2322]),

			.SO(gen[2380]),
			.S(gen[2381]),
			.SE(gen[2382]),

			.SELF(gen[2321]),
			.cell_state(gen[2321])
		); 

/******************* CELL 2322 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2322 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2261]),
			.N(gen[2262]),
			.NE(gen[2263]),

			.O(gen[2321]),
			.E(gen[2323]),

			.SO(gen[2381]),
			.S(gen[2382]),
			.SE(gen[2383]),

			.SELF(gen[2322]),
			.cell_state(gen[2322])
		); 

/******************* CELL 2323 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2323 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2262]),
			.N(gen[2263]),
			.NE(gen[2264]),

			.O(gen[2322]),
			.E(gen[2324]),

			.SO(gen[2382]),
			.S(gen[2383]),
			.SE(gen[2384]),

			.SELF(gen[2323]),
			.cell_state(gen[2323])
		); 

/******************* CELL 2324 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2324 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2263]),
			.N(gen[2264]),
			.NE(gen[2265]),

			.O(gen[2323]),
			.E(gen[2325]),

			.SO(gen[2383]),
			.S(gen[2384]),
			.SE(gen[2385]),

			.SELF(gen[2324]),
			.cell_state(gen[2324])
		); 

/******************* CELL 2325 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2325 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2264]),
			.N(gen[2265]),
			.NE(gen[2266]),

			.O(gen[2324]),
			.E(gen[2326]),

			.SO(gen[2384]),
			.S(gen[2385]),
			.SE(gen[2386]),

			.SELF(gen[2325]),
			.cell_state(gen[2325])
		); 

/******************* CELL 2326 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2326 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2265]),
			.N(gen[2266]),
			.NE(gen[2267]),

			.O(gen[2325]),
			.E(gen[2327]),

			.SO(gen[2385]),
			.S(gen[2386]),
			.SE(gen[2387]),

			.SELF(gen[2326]),
			.cell_state(gen[2326])
		); 

/******************* CELL 2327 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2327 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2266]),
			.N(gen[2267]),
			.NE(gen[2268]),

			.O(gen[2326]),
			.E(gen[2328]),

			.SO(gen[2386]),
			.S(gen[2387]),
			.SE(gen[2388]),

			.SELF(gen[2327]),
			.cell_state(gen[2327])
		); 

/******************* CELL 2328 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2328 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2267]),
			.N(gen[2268]),
			.NE(gen[2269]),

			.O(gen[2327]),
			.E(gen[2329]),

			.SO(gen[2387]),
			.S(gen[2388]),
			.SE(gen[2389]),

			.SELF(gen[2328]),
			.cell_state(gen[2328])
		); 

/******************* CELL 2329 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2329 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2268]),
			.N(gen[2269]),
			.NE(gen[2270]),

			.O(gen[2328]),
			.E(gen[2330]),

			.SO(gen[2388]),
			.S(gen[2389]),
			.SE(gen[2390]),

			.SELF(gen[2329]),
			.cell_state(gen[2329])
		); 

/******************* CELL 2330 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2330 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2269]),
			.N(gen[2270]),
			.NE(gen[2271]),

			.O(gen[2329]),
			.E(gen[2331]),

			.SO(gen[2389]),
			.S(gen[2390]),
			.SE(gen[2391]),

			.SELF(gen[2330]),
			.cell_state(gen[2330])
		); 

/******************* CELL 2331 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2331 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2270]),
			.N(gen[2271]),
			.NE(gen[2272]),

			.O(gen[2330]),
			.E(gen[2332]),

			.SO(gen[2390]),
			.S(gen[2391]),
			.SE(gen[2392]),

			.SELF(gen[2331]),
			.cell_state(gen[2331])
		); 

/******************* CELL 2332 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2332 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2271]),
			.N(gen[2272]),
			.NE(gen[2273]),

			.O(gen[2331]),
			.E(gen[2333]),

			.SO(gen[2391]),
			.S(gen[2392]),
			.SE(gen[2393]),

			.SELF(gen[2332]),
			.cell_state(gen[2332])
		); 

/******************* CELL 2333 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2333 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2272]),
			.N(gen[2273]),
			.NE(gen[2274]),

			.O(gen[2332]),
			.E(gen[2334]),

			.SO(gen[2392]),
			.S(gen[2393]),
			.SE(gen[2394]),

			.SELF(gen[2333]),
			.cell_state(gen[2333])
		); 

/******************* CELL 2334 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2334 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2273]),
			.N(gen[2274]),
			.NE(gen[2275]),

			.O(gen[2333]),
			.E(gen[2335]),

			.SO(gen[2393]),
			.S(gen[2394]),
			.SE(gen[2395]),

			.SELF(gen[2334]),
			.cell_state(gen[2334])
		); 

/******************* CELL 2335 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2335 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2274]),
			.N(gen[2275]),
			.NE(gen[2276]),

			.O(gen[2334]),
			.E(gen[2336]),

			.SO(gen[2394]),
			.S(gen[2395]),
			.SE(gen[2396]),

			.SELF(gen[2335]),
			.cell_state(gen[2335])
		); 

/******************* CELL 2336 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2336 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2275]),
			.N(gen[2276]),
			.NE(gen[2277]),

			.O(gen[2335]),
			.E(gen[2337]),

			.SO(gen[2395]),
			.S(gen[2396]),
			.SE(gen[2397]),

			.SELF(gen[2336]),
			.cell_state(gen[2336])
		); 

/******************* CELL 2337 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2337 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2276]),
			.N(gen[2277]),
			.NE(gen[2278]),

			.O(gen[2336]),
			.E(gen[2338]),

			.SO(gen[2396]),
			.S(gen[2397]),
			.SE(gen[2398]),

			.SELF(gen[2337]),
			.cell_state(gen[2337])
		); 

/******************* CELL 2338 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2338 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2277]),
			.N(gen[2278]),
			.NE(gen[2279]),

			.O(gen[2337]),
			.E(gen[2339]),

			.SO(gen[2397]),
			.S(gen[2398]),
			.SE(gen[2399]),

			.SELF(gen[2338]),
			.cell_state(gen[2338])
		); 

/******************* CELL 2339 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2339 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2278]),
			.N(gen[2279]),
			.NE(gen[2278]),

			.O(gen[2338]),
			.E(gen[2338]),

			.SO(gen[2398]),
			.S(gen[2399]),
			.SE(gen[2398]),

			.SELF(gen[2339]),
			.cell_state(gen[2339])
		); 

/******************* CELL 2340 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2340 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2281]),
			.N(gen[2280]),
			.NE(gen[2281]),

			.O(gen[2341]),
			.E(gen[2341]),

			.SO(gen[2401]),
			.S(gen[2400]),
			.SE(gen[2401]),

			.SELF(gen[2340]),
			.cell_state(gen[2340])
		); 

/******************* CELL 2341 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2341 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2280]),
			.N(gen[2281]),
			.NE(gen[2282]),

			.O(gen[2340]),
			.E(gen[2342]),

			.SO(gen[2400]),
			.S(gen[2401]),
			.SE(gen[2402]),

			.SELF(gen[2341]),
			.cell_state(gen[2341])
		); 

/******************* CELL 2342 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2342 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2281]),
			.N(gen[2282]),
			.NE(gen[2283]),

			.O(gen[2341]),
			.E(gen[2343]),

			.SO(gen[2401]),
			.S(gen[2402]),
			.SE(gen[2403]),

			.SELF(gen[2342]),
			.cell_state(gen[2342])
		); 

/******************* CELL 2343 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2343 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2282]),
			.N(gen[2283]),
			.NE(gen[2284]),

			.O(gen[2342]),
			.E(gen[2344]),

			.SO(gen[2402]),
			.S(gen[2403]),
			.SE(gen[2404]),

			.SELF(gen[2343]),
			.cell_state(gen[2343])
		); 

/******************* CELL 2344 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2344 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2283]),
			.N(gen[2284]),
			.NE(gen[2285]),

			.O(gen[2343]),
			.E(gen[2345]),

			.SO(gen[2403]),
			.S(gen[2404]),
			.SE(gen[2405]),

			.SELF(gen[2344]),
			.cell_state(gen[2344])
		); 

/******************* CELL 2345 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2345 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2284]),
			.N(gen[2285]),
			.NE(gen[2286]),

			.O(gen[2344]),
			.E(gen[2346]),

			.SO(gen[2404]),
			.S(gen[2405]),
			.SE(gen[2406]),

			.SELF(gen[2345]),
			.cell_state(gen[2345])
		); 

/******************* CELL 2346 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2346 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2285]),
			.N(gen[2286]),
			.NE(gen[2287]),

			.O(gen[2345]),
			.E(gen[2347]),

			.SO(gen[2405]),
			.S(gen[2406]),
			.SE(gen[2407]),

			.SELF(gen[2346]),
			.cell_state(gen[2346])
		); 

/******************* CELL 2347 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2347 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2286]),
			.N(gen[2287]),
			.NE(gen[2288]),

			.O(gen[2346]),
			.E(gen[2348]),

			.SO(gen[2406]),
			.S(gen[2407]),
			.SE(gen[2408]),

			.SELF(gen[2347]),
			.cell_state(gen[2347])
		); 

/******************* CELL 2348 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2348 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2287]),
			.N(gen[2288]),
			.NE(gen[2289]),

			.O(gen[2347]),
			.E(gen[2349]),

			.SO(gen[2407]),
			.S(gen[2408]),
			.SE(gen[2409]),

			.SELF(gen[2348]),
			.cell_state(gen[2348])
		); 

/******************* CELL 2349 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2349 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2288]),
			.N(gen[2289]),
			.NE(gen[2290]),

			.O(gen[2348]),
			.E(gen[2350]),

			.SO(gen[2408]),
			.S(gen[2409]),
			.SE(gen[2410]),

			.SELF(gen[2349]),
			.cell_state(gen[2349])
		); 

/******************* CELL 2350 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2350 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2289]),
			.N(gen[2290]),
			.NE(gen[2291]),

			.O(gen[2349]),
			.E(gen[2351]),

			.SO(gen[2409]),
			.S(gen[2410]),
			.SE(gen[2411]),

			.SELF(gen[2350]),
			.cell_state(gen[2350])
		); 

/******************* CELL 2351 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2351 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2290]),
			.N(gen[2291]),
			.NE(gen[2292]),

			.O(gen[2350]),
			.E(gen[2352]),

			.SO(gen[2410]),
			.S(gen[2411]),
			.SE(gen[2412]),

			.SELF(gen[2351]),
			.cell_state(gen[2351])
		); 

/******************* CELL 2352 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2352 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2291]),
			.N(gen[2292]),
			.NE(gen[2293]),

			.O(gen[2351]),
			.E(gen[2353]),

			.SO(gen[2411]),
			.S(gen[2412]),
			.SE(gen[2413]),

			.SELF(gen[2352]),
			.cell_state(gen[2352])
		); 

/******************* CELL 2353 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2353 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2292]),
			.N(gen[2293]),
			.NE(gen[2294]),

			.O(gen[2352]),
			.E(gen[2354]),

			.SO(gen[2412]),
			.S(gen[2413]),
			.SE(gen[2414]),

			.SELF(gen[2353]),
			.cell_state(gen[2353])
		); 

/******************* CELL 2354 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2354 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2293]),
			.N(gen[2294]),
			.NE(gen[2295]),

			.O(gen[2353]),
			.E(gen[2355]),

			.SO(gen[2413]),
			.S(gen[2414]),
			.SE(gen[2415]),

			.SELF(gen[2354]),
			.cell_state(gen[2354])
		); 

/******************* CELL 2355 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2355 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2294]),
			.N(gen[2295]),
			.NE(gen[2296]),

			.O(gen[2354]),
			.E(gen[2356]),

			.SO(gen[2414]),
			.S(gen[2415]),
			.SE(gen[2416]),

			.SELF(gen[2355]),
			.cell_state(gen[2355])
		); 

/******************* CELL 2356 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2356 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2295]),
			.N(gen[2296]),
			.NE(gen[2297]),

			.O(gen[2355]),
			.E(gen[2357]),

			.SO(gen[2415]),
			.S(gen[2416]),
			.SE(gen[2417]),

			.SELF(gen[2356]),
			.cell_state(gen[2356])
		); 

/******************* CELL 2357 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2357 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2296]),
			.N(gen[2297]),
			.NE(gen[2298]),

			.O(gen[2356]),
			.E(gen[2358]),

			.SO(gen[2416]),
			.S(gen[2417]),
			.SE(gen[2418]),

			.SELF(gen[2357]),
			.cell_state(gen[2357])
		); 

/******************* CELL 2358 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2358 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2297]),
			.N(gen[2298]),
			.NE(gen[2299]),

			.O(gen[2357]),
			.E(gen[2359]),

			.SO(gen[2417]),
			.S(gen[2418]),
			.SE(gen[2419]),

			.SELF(gen[2358]),
			.cell_state(gen[2358])
		); 

/******************* CELL 2359 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2359 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2298]),
			.N(gen[2299]),
			.NE(gen[2300]),

			.O(gen[2358]),
			.E(gen[2360]),

			.SO(gen[2418]),
			.S(gen[2419]),
			.SE(gen[2420]),

			.SELF(gen[2359]),
			.cell_state(gen[2359])
		); 

/******************* CELL 2360 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2360 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2299]),
			.N(gen[2300]),
			.NE(gen[2301]),

			.O(gen[2359]),
			.E(gen[2361]),

			.SO(gen[2419]),
			.S(gen[2420]),
			.SE(gen[2421]),

			.SELF(gen[2360]),
			.cell_state(gen[2360])
		); 

/******************* CELL 2361 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2361 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2300]),
			.N(gen[2301]),
			.NE(gen[2302]),

			.O(gen[2360]),
			.E(gen[2362]),

			.SO(gen[2420]),
			.S(gen[2421]),
			.SE(gen[2422]),

			.SELF(gen[2361]),
			.cell_state(gen[2361])
		); 

/******************* CELL 2362 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2362 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2301]),
			.N(gen[2302]),
			.NE(gen[2303]),

			.O(gen[2361]),
			.E(gen[2363]),

			.SO(gen[2421]),
			.S(gen[2422]),
			.SE(gen[2423]),

			.SELF(gen[2362]),
			.cell_state(gen[2362])
		); 

/******************* CELL 2363 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2363 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2302]),
			.N(gen[2303]),
			.NE(gen[2304]),

			.O(gen[2362]),
			.E(gen[2364]),

			.SO(gen[2422]),
			.S(gen[2423]),
			.SE(gen[2424]),

			.SELF(gen[2363]),
			.cell_state(gen[2363])
		); 

/******************* CELL 2364 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2364 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2303]),
			.N(gen[2304]),
			.NE(gen[2305]),

			.O(gen[2363]),
			.E(gen[2365]),

			.SO(gen[2423]),
			.S(gen[2424]),
			.SE(gen[2425]),

			.SELF(gen[2364]),
			.cell_state(gen[2364])
		); 

/******************* CELL 2365 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2365 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2304]),
			.N(gen[2305]),
			.NE(gen[2306]),

			.O(gen[2364]),
			.E(gen[2366]),

			.SO(gen[2424]),
			.S(gen[2425]),
			.SE(gen[2426]),

			.SELF(gen[2365]),
			.cell_state(gen[2365])
		); 

/******************* CELL 2366 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2366 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2305]),
			.N(gen[2306]),
			.NE(gen[2307]),

			.O(gen[2365]),
			.E(gen[2367]),

			.SO(gen[2425]),
			.S(gen[2426]),
			.SE(gen[2427]),

			.SELF(gen[2366]),
			.cell_state(gen[2366])
		); 

/******************* CELL 2367 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2367 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2306]),
			.N(gen[2307]),
			.NE(gen[2308]),

			.O(gen[2366]),
			.E(gen[2368]),

			.SO(gen[2426]),
			.S(gen[2427]),
			.SE(gen[2428]),

			.SELF(gen[2367]),
			.cell_state(gen[2367])
		); 

/******************* CELL 2368 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2368 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2307]),
			.N(gen[2308]),
			.NE(gen[2309]),

			.O(gen[2367]),
			.E(gen[2369]),

			.SO(gen[2427]),
			.S(gen[2428]),
			.SE(gen[2429]),

			.SELF(gen[2368]),
			.cell_state(gen[2368])
		); 

/******************* CELL 2369 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2369 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2308]),
			.N(gen[2309]),
			.NE(gen[2310]),

			.O(gen[2368]),
			.E(gen[2370]),

			.SO(gen[2428]),
			.S(gen[2429]),
			.SE(gen[2430]),

			.SELF(gen[2369]),
			.cell_state(gen[2369])
		); 

/******************* CELL 2370 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2370 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2309]),
			.N(gen[2310]),
			.NE(gen[2311]),

			.O(gen[2369]),
			.E(gen[2371]),

			.SO(gen[2429]),
			.S(gen[2430]),
			.SE(gen[2431]),

			.SELF(gen[2370]),
			.cell_state(gen[2370])
		); 

/******************* CELL 2371 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2371 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2310]),
			.N(gen[2311]),
			.NE(gen[2312]),

			.O(gen[2370]),
			.E(gen[2372]),

			.SO(gen[2430]),
			.S(gen[2431]),
			.SE(gen[2432]),

			.SELF(gen[2371]),
			.cell_state(gen[2371])
		); 

/******************* CELL 2372 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2372 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2311]),
			.N(gen[2312]),
			.NE(gen[2313]),

			.O(gen[2371]),
			.E(gen[2373]),

			.SO(gen[2431]),
			.S(gen[2432]),
			.SE(gen[2433]),

			.SELF(gen[2372]),
			.cell_state(gen[2372])
		); 

/******************* CELL 2373 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2373 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2312]),
			.N(gen[2313]),
			.NE(gen[2314]),

			.O(gen[2372]),
			.E(gen[2374]),

			.SO(gen[2432]),
			.S(gen[2433]),
			.SE(gen[2434]),

			.SELF(gen[2373]),
			.cell_state(gen[2373])
		); 

/******************* CELL 2374 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2374 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2313]),
			.N(gen[2314]),
			.NE(gen[2315]),

			.O(gen[2373]),
			.E(gen[2375]),

			.SO(gen[2433]),
			.S(gen[2434]),
			.SE(gen[2435]),

			.SELF(gen[2374]),
			.cell_state(gen[2374])
		); 

/******************* CELL 2375 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2375 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2314]),
			.N(gen[2315]),
			.NE(gen[2316]),

			.O(gen[2374]),
			.E(gen[2376]),

			.SO(gen[2434]),
			.S(gen[2435]),
			.SE(gen[2436]),

			.SELF(gen[2375]),
			.cell_state(gen[2375])
		); 

/******************* CELL 2376 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2376 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2315]),
			.N(gen[2316]),
			.NE(gen[2317]),

			.O(gen[2375]),
			.E(gen[2377]),

			.SO(gen[2435]),
			.S(gen[2436]),
			.SE(gen[2437]),

			.SELF(gen[2376]),
			.cell_state(gen[2376])
		); 

/******************* CELL 2377 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2377 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2316]),
			.N(gen[2317]),
			.NE(gen[2318]),

			.O(gen[2376]),
			.E(gen[2378]),

			.SO(gen[2436]),
			.S(gen[2437]),
			.SE(gen[2438]),

			.SELF(gen[2377]),
			.cell_state(gen[2377])
		); 

/******************* CELL 2378 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2378 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2317]),
			.N(gen[2318]),
			.NE(gen[2319]),

			.O(gen[2377]),
			.E(gen[2379]),

			.SO(gen[2437]),
			.S(gen[2438]),
			.SE(gen[2439]),

			.SELF(gen[2378]),
			.cell_state(gen[2378])
		); 

/******************* CELL 2379 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2379 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2318]),
			.N(gen[2319]),
			.NE(gen[2320]),

			.O(gen[2378]),
			.E(gen[2380]),

			.SO(gen[2438]),
			.S(gen[2439]),
			.SE(gen[2440]),

			.SELF(gen[2379]),
			.cell_state(gen[2379])
		); 

/******************* CELL 2380 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2380 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2319]),
			.N(gen[2320]),
			.NE(gen[2321]),

			.O(gen[2379]),
			.E(gen[2381]),

			.SO(gen[2439]),
			.S(gen[2440]),
			.SE(gen[2441]),

			.SELF(gen[2380]),
			.cell_state(gen[2380])
		); 

/******************* CELL 2381 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2381 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2320]),
			.N(gen[2321]),
			.NE(gen[2322]),

			.O(gen[2380]),
			.E(gen[2382]),

			.SO(gen[2440]),
			.S(gen[2441]),
			.SE(gen[2442]),

			.SELF(gen[2381]),
			.cell_state(gen[2381])
		); 

/******************* CELL 2382 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2382 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2321]),
			.N(gen[2322]),
			.NE(gen[2323]),

			.O(gen[2381]),
			.E(gen[2383]),

			.SO(gen[2441]),
			.S(gen[2442]),
			.SE(gen[2443]),

			.SELF(gen[2382]),
			.cell_state(gen[2382])
		); 

/******************* CELL 2383 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2383 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2322]),
			.N(gen[2323]),
			.NE(gen[2324]),

			.O(gen[2382]),
			.E(gen[2384]),

			.SO(gen[2442]),
			.S(gen[2443]),
			.SE(gen[2444]),

			.SELF(gen[2383]),
			.cell_state(gen[2383])
		); 

/******************* CELL 2384 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2384 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2323]),
			.N(gen[2324]),
			.NE(gen[2325]),

			.O(gen[2383]),
			.E(gen[2385]),

			.SO(gen[2443]),
			.S(gen[2444]),
			.SE(gen[2445]),

			.SELF(gen[2384]),
			.cell_state(gen[2384])
		); 

/******************* CELL 2385 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2385 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2324]),
			.N(gen[2325]),
			.NE(gen[2326]),

			.O(gen[2384]),
			.E(gen[2386]),

			.SO(gen[2444]),
			.S(gen[2445]),
			.SE(gen[2446]),

			.SELF(gen[2385]),
			.cell_state(gen[2385])
		); 

/******************* CELL 2386 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2386 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2325]),
			.N(gen[2326]),
			.NE(gen[2327]),

			.O(gen[2385]),
			.E(gen[2387]),

			.SO(gen[2445]),
			.S(gen[2446]),
			.SE(gen[2447]),

			.SELF(gen[2386]),
			.cell_state(gen[2386])
		); 

/******************* CELL 2387 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2387 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2326]),
			.N(gen[2327]),
			.NE(gen[2328]),

			.O(gen[2386]),
			.E(gen[2388]),

			.SO(gen[2446]),
			.S(gen[2447]),
			.SE(gen[2448]),

			.SELF(gen[2387]),
			.cell_state(gen[2387])
		); 

/******************* CELL 2388 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2388 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2327]),
			.N(gen[2328]),
			.NE(gen[2329]),

			.O(gen[2387]),
			.E(gen[2389]),

			.SO(gen[2447]),
			.S(gen[2448]),
			.SE(gen[2449]),

			.SELF(gen[2388]),
			.cell_state(gen[2388])
		); 

/******************* CELL 2389 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2389 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2328]),
			.N(gen[2329]),
			.NE(gen[2330]),

			.O(gen[2388]),
			.E(gen[2390]),

			.SO(gen[2448]),
			.S(gen[2449]),
			.SE(gen[2450]),

			.SELF(gen[2389]),
			.cell_state(gen[2389])
		); 

/******************* CELL 2390 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2390 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2329]),
			.N(gen[2330]),
			.NE(gen[2331]),

			.O(gen[2389]),
			.E(gen[2391]),

			.SO(gen[2449]),
			.S(gen[2450]),
			.SE(gen[2451]),

			.SELF(gen[2390]),
			.cell_state(gen[2390])
		); 

/******************* CELL 2391 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2391 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2330]),
			.N(gen[2331]),
			.NE(gen[2332]),

			.O(gen[2390]),
			.E(gen[2392]),

			.SO(gen[2450]),
			.S(gen[2451]),
			.SE(gen[2452]),

			.SELF(gen[2391]),
			.cell_state(gen[2391])
		); 

/******************* CELL 2392 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2392 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2331]),
			.N(gen[2332]),
			.NE(gen[2333]),

			.O(gen[2391]),
			.E(gen[2393]),

			.SO(gen[2451]),
			.S(gen[2452]),
			.SE(gen[2453]),

			.SELF(gen[2392]),
			.cell_state(gen[2392])
		); 

/******************* CELL 2393 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2393 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2332]),
			.N(gen[2333]),
			.NE(gen[2334]),

			.O(gen[2392]),
			.E(gen[2394]),

			.SO(gen[2452]),
			.S(gen[2453]),
			.SE(gen[2454]),

			.SELF(gen[2393]),
			.cell_state(gen[2393])
		); 

/******************* CELL 2394 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2394 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2333]),
			.N(gen[2334]),
			.NE(gen[2335]),

			.O(gen[2393]),
			.E(gen[2395]),

			.SO(gen[2453]),
			.S(gen[2454]),
			.SE(gen[2455]),

			.SELF(gen[2394]),
			.cell_state(gen[2394])
		); 

/******************* CELL 2395 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2395 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2334]),
			.N(gen[2335]),
			.NE(gen[2336]),

			.O(gen[2394]),
			.E(gen[2396]),

			.SO(gen[2454]),
			.S(gen[2455]),
			.SE(gen[2456]),

			.SELF(gen[2395]),
			.cell_state(gen[2395])
		); 

/******************* CELL 2396 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2396 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2335]),
			.N(gen[2336]),
			.NE(gen[2337]),

			.O(gen[2395]),
			.E(gen[2397]),

			.SO(gen[2455]),
			.S(gen[2456]),
			.SE(gen[2457]),

			.SELF(gen[2396]),
			.cell_state(gen[2396])
		); 

/******************* CELL 2397 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2397 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2336]),
			.N(gen[2337]),
			.NE(gen[2338]),

			.O(gen[2396]),
			.E(gen[2398]),

			.SO(gen[2456]),
			.S(gen[2457]),
			.SE(gen[2458]),

			.SELF(gen[2397]),
			.cell_state(gen[2397])
		); 

/******************* CELL 2398 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2398 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2337]),
			.N(gen[2338]),
			.NE(gen[2339]),

			.O(gen[2397]),
			.E(gen[2399]),

			.SO(gen[2457]),
			.S(gen[2458]),
			.SE(gen[2459]),

			.SELF(gen[2398]),
			.cell_state(gen[2398])
		); 

/******************* CELL 2399 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2399 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2338]),
			.N(gen[2339]),
			.NE(gen[2338]),

			.O(gen[2398]),
			.E(gen[2398]),

			.SO(gen[2458]),
			.S(gen[2459]),
			.SE(gen[2458]),

			.SELF(gen[2399]),
			.cell_state(gen[2399])
		); 

/******************* CELL 2400 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2400 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2341]),
			.N(gen[2340]),
			.NE(gen[2341]),

			.O(gen[2401]),
			.E(gen[2401]),

			.SO(gen[2461]),
			.S(gen[2460]),
			.SE(gen[2461]),

			.SELF(gen[2400]),
			.cell_state(gen[2400])
		); 

/******************* CELL 2401 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2401 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2340]),
			.N(gen[2341]),
			.NE(gen[2342]),

			.O(gen[2400]),
			.E(gen[2402]),

			.SO(gen[2460]),
			.S(gen[2461]),
			.SE(gen[2462]),

			.SELF(gen[2401]),
			.cell_state(gen[2401])
		); 

/******************* CELL 2402 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2402 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2341]),
			.N(gen[2342]),
			.NE(gen[2343]),

			.O(gen[2401]),
			.E(gen[2403]),

			.SO(gen[2461]),
			.S(gen[2462]),
			.SE(gen[2463]),

			.SELF(gen[2402]),
			.cell_state(gen[2402])
		); 

/******************* CELL 2403 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2403 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2342]),
			.N(gen[2343]),
			.NE(gen[2344]),

			.O(gen[2402]),
			.E(gen[2404]),

			.SO(gen[2462]),
			.S(gen[2463]),
			.SE(gen[2464]),

			.SELF(gen[2403]),
			.cell_state(gen[2403])
		); 

/******************* CELL 2404 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2404 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2343]),
			.N(gen[2344]),
			.NE(gen[2345]),

			.O(gen[2403]),
			.E(gen[2405]),

			.SO(gen[2463]),
			.S(gen[2464]),
			.SE(gen[2465]),

			.SELF(gen[2404]),
			.cell_state(gen[2404])
		); 

/******************* CELL 2405 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2405 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2344]),
			.N(gen[2345]),
			.NE(gen[2346]),

			.O(gen[2404]),
			.E(gen[2406]),

			.SO(gen[2464]),
			.S(gen[2465]),
			.SE(gen[2466]),

			.SELF(gen[2405]),
			.cell_state(gen[2405])
		); 

/******************* CELL 2406 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2406 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2345]),
			.N(gen[2346]),
			.NE(gen[2347]),

			.O(gen[2405]),
			.E(gen[2407]),

			.SO(gen[2465]),
			.S(gen[2466]),
			.SE(gen[2467]),

			.SELF(gen[2406]),
			.cell_state(gen[2406])
		); 

/******************* CELL 2407 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2407 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2346]),
			.N(gen[2347]),
			.NE(gen[2348]),

			.O(gen[2406]),
			.E(gen[2408]),

			.SO(gen[2466]),
			.S(gen[2467]),
			.SE(gen[2468]),

			.SELF(gen[2407]),
			.cell_state(gen[2407])
		); 

/******************* CELL 2408 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2408 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2347]),
			.N(gen[2348]),
			.NE(gen[2349]),

			.O(gen[2407]),
			.E(gen[2409]),

			.SO(gen[2467]),
			.S(gen[2468]),
			.SE(gen[2469]),

			.SELF(gen[2408]),
			.cell_state(gen[2408])
		); 

/******************* CELL 2409 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2409 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2348]),
			.N(gen[2349]),
			.NE(gen[2350]),

			.O(gen[2408]),
			.E(gen[2410]),

			.SO(gen[2468]),
			.S(gen[2469]),
			.SE(gen[2470]),

			.SELF(gen[2409]),
			.cell_state(gen[2409])
		); 

/******************* CELL 2410 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2410 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2349]),
			.N(gen[2350]),
			.NE(gen[2351]),

			.O(gen[2409]),
			.E(gen[2411]),

			.SO(gen[2469]),
			.S(gen[2470]),
			.SE(gen[2471]),

			.SELF(gen[2410]),
			.cell_state(gen[2410])
		); 

/******************* CELL 2411 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2411 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2350]),
			.N(gen[2351]),
			.NE(gen[2352]),

			.O(gen[2410]),
			.E(gen[2412]),

			.SO(gen[2470]),
			.S(gen[2471]),
			.SE(gen[2472]),

			.SELF(gen[2411]),
			.cell_state(gen[2411])
		); 

/******************* CELL 2412 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2412 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2351]),
			.N(gen[2352]),
			.NE(gen[2353]),

			.O(gen[2411]),
			.E(gen[2413]),

			.SO(gen[2471]),
			.S(gen[2472]),
			.SE(gen[2473]),

			.SELF(gen[2412]),
			.cell_state(gen[2412])
		); 

/******************* CELL 2413 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2413 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2352]),
			.N(gen[2353]),
			.NE(gen[2354]),

			.O(gen[2412]),
			.E(gen[2414]),

			.SO(gen[2472]),
			.S(gen[2473]),
			.SE(gen[2474]),

			.SELF(gen[2413]),
			.cell_state(gen[2413])
		); 

/******************* CELL 2414 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2414 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2353]),
			.N(gen[2354]),
			.NE(gen[2355]),

			.O(gen[2413]),
			.E(gen[2415]),

			.SO(gen[2473]),
			.S(gen[2474]),
			.SE(gen[2475]),

			.SELF(gen[2414]),
			.cell_state(gen[2414])
		); 

/******************* CELL 2415 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2415 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2354]),
			.N(gen[2355]),
			.NE(gen[2356]),

			.O(gen[2414]),
			.E(gen[2416]),

			.SO(gen[2474]),
			.S(gen[2475]),
			.SE(gen[2476]),

			.SELF(gen[2415]),
			.cell_state(gen[2415])
		); 

/******************* CELL 2416 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2416 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2355]),
			.N(gen[2356]),
			.NE(gen[2357]),

			.O(gen[2415]),
			.E(gen[2417]),

			.SO(gen[2475]),
			.S(gen[2476]),
			.SE(gen[2477]),

			.SELF(gen[2416]),
			.cell_state(gen[2416])
		); 

/******************* CELL 2417 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2417 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2356]),
			.N(gen[2357]),
			.NE(gen[2358]),

			.O(gen[2416]),
			.E(gen[2418]),

			.SO(gen[2476]),
			.S(gen[2477]),
			.SE(gen[2478]),

			.SELF(gen[2417]),
			.cell_state(gen[2417])
		); 

/******************* CELL 2418 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2418 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2357]),
			.N(gen[2358]),
			.NE(gen[2359]),

			.O(gen[2417]),
			.E(gen[2419]),

			.SO(gen[2477]),
			.S(gen[2478]),
			.SE(gen[2479]),

			.SELF(gen[2418]),
			.cell_state(gen[2418])
		); 

/******************* CELL 2419 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2419 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2358]),
			.N(gen[2359]),
			.NE(gen[2360]),

			.O(gen[2418]),
			.E(gen[2420]),

			.SO(gen[2478]),
			.S(gen[2479]),
			.SE(gen[2480]),

			.SELF(gen[2419]),
			.cell_state(gen[2419])
		); 

/******************* CELL 2420 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2420 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2359]),
			.N(gen[2360]),
			.NE(gen[2361]),

			.O(gen[2419]),
			.E(gen[2421]),

			.SO(gen[2479]),
			.S(gen[2480]),
			.SE(gen[2481]),

			.SELF(gen[2420]),
			.cell_state(gen[2420])
		); 

/******************* CELL 2421 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2421 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2360]),
			.N(gen[2361]),
			.NE(gen[2362]),

			.O(gen[2420]),
			.E(gen[2422]),

			.SO(gen[2480]),
			.S(gen[2481]),
			.SE(gen[2482]),

			.SELF(gen[2421]),
			.cell_state(gen[2421])
		); 

/******************* CELL 2422 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2422 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2361]),
			.N(gen[2362]),
			.NE(gen[2363]),

			.O(gen[2421]),
			.E(gen[2423]),

			.SO(gen[2481]),
			.S(gen[2482]),
			.SE(gen[2483]),

			.SELF(gen[2422]),
			.cell_state(gen[2422])
		); 

/******************* CELL 2423 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2423 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2362]),
			.N(gen[2363]),
			.NE(gen[2364]),

			.O(gen[2422]),
			.E(gen[2424]),

			.SO(gen[2482]),
			.S(gen[2483]),
			.SE(gen[2484]),

			.SELF(gen[2423]),
			.cell_state(gen[2423])
		); 

/******************* CELL 2424 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2424 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2363]),
			.N(gen[2364]),
			.NE(gen[2365]),

			.O(gen[2423]),
			.E(gen[2425]),

			.SO(gen[2483]),
			.S(gen[2484]),
			.SE(gen[2485]),

			.SELF(gen[2424]),
			.cell_state(gen[2424])
		); 

/******************* CELL 2425 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2425 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2364]),
			.N(gen[2365]),
			.NE(gen[2366]),

			.O(gen[2424]),
			.E(gen[2426]),

			.SO(gen[2484]),
			.S(gen[2485]),
			.SE(gen[2486]),

			.SELF(gen[2425]),
			.cell_state(gen[2425])
		); 

/******************* CELL 2426 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2426 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2365]),
			.N(gen[2366]),
			.NE(gen[2367]),

			.O(gen[2425]),
			.E(gen[2427]),

			.SO(gen[2485]),
			.S(gen[2486]),
			.SE(gen[2487]),

			.SELF(gen[2426]),
			.cell_state(gen[2426])
		); 

/******************* CELL 2427 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2427 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2366]),
			.N(gen[2367]),
			.NE(gen[2368]),

			.O(gen[2426]),
			.E(gen[2428]),

			.SO(gen[2486]),
			.S(gen[2487]),
			.SE(gen[2488]),

			.SELF(gen[2427]),
			.cell_state(gen[2427])
		); 

/******************* CELL 2428 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2428 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2367]),
			.N(gen[2368]),
			.NE(gen[2369]),

			.O(gen[2427]),
			.E(gen[2429]),

			.SO(gen[2487]),
			.S(gen[2488]),
			.SE(gen[2489]),

			.SELF(gen[2428]),
			.cell_state(gen[2428])
		); 

/******************* CELL 2429 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2429 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2368]),
			.N(gen[2369]),
			.NE(gen[2370]),

			.O(gen[2428]),
			.E(gen[2430]),

			.SO(gen[2488]),
			.S(gen[2489]),
			.SE(gen[2490]),

			.SELF(gen[2429]),
			.cell_state(gen[2429])
		); 

/******************* CELL 2430 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2430 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2369]),
			.N(gen[2370]),
			.NE(gen[2371]),

			.O(gen[2429]),
			.E(gen[2431]),

			.SO(gen[2489]),
			.S(gen[2490]),
			.SE(gen[2491]),

			.SELF(gen[2430]),
			.cell_state(gen[2430])
		); 

/******************* CELL 2431 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2431 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2370]),
			.N(gen[2371]),
			.NE(gen[2372]),

			.O(gen[2430]),
			.E(gen[2432]),

			.SO(gen[2490]),
			.S(gen[2491]),
			.SE(gen[2492]),

			.SELF(gen[2431]),
			.cell_state(gen[2431])
		); 

/******************* CELL 2432 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2432 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2371]),
			.N(gen[2372]),
			.NE(gen[2373]),

			.O(gen[2431]),
			.E(gen[2433]),

			.SO(gen[2491]),
			.S(gen[2492]),
			.SE(gen[2493]),

			.SELF(gen[2432]),
			.cell_state(gen[2432])
		); 

/******************* CELL 2433 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2433 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2372]),
			.N(gen[2373]),
			.NE(gen[2374]),

			.O(gen[2432]),
			.E(gen[2434]),

			.SO(gen[2492]),
			.S(gen[2493]),
			.SE(gen[2494]),

			.SELF(gen[2433]),
			.cell_state(gen[2433])
		); 

/******************* CELL 2434 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2434 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2373]),
			.N(gen[2374]),
			.NE(gen[2375]),

			.O(gen[2433]),
			.E(gen[2435]),

			.SO(gen[2493]),
			.S(gen[2494]),
			.SE(gen[2495]),

			.SELF(gen[2434]),
			.cell_state(gen[2434])
		); 

/******************* CELL 2435 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2435 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2374]),
			.N(gen[2375]),
			.NE(gen[2376]),

			.O(gen[2434]),
			.E(gen[2436]),

			.SO(gen[2494]),
			.S(gen[2495]),
			.SE(gen[2496]),

			.SELF(gen[2435]),
			.cell_state(gen[2435])
		); 

/******************* CELL 2436 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2436 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2375]),
			.N(gen[2376]),
			.NE(gen[2377]),

			.O(gen[2435]),
			.E(gen[2437]),

			.SO(gen[2495]),
			.S(gen[2496]),
			.SE(gen[2497]),

			.SELF(gen[2436]),
			.cell_state(gen[2436])
		); 

/******************* CELL 2437 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2437 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2376]),
			.N(gen[2377]),
			.NE(gen[2378]),

			.O(gen[2436]),
			.E(gen[2438]),

			.SO(gen[2496]),
			.S(gen[2497]),
			.SE(gen[2498]),

			.SELF(gen[2437]),
			.cell_state(gen[2437])
		); 

/******************* CELL 2438 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2438 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2377]),
			.N(gen[2378]),
			.NE(gen[2379]),

			.O(gen[2437]),
			.E(gen[2439]),

			.SO(gen[2497]),
			.S(gen[2498]),
			.SE(gen[2499]),

			.SELF(gen[2438]),
			.cell_state(gen[2438])
		); 

/******************* CELL 2439 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2439 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2378]),
			.N(gen[2379]),
			.NE(gen[2380]),

			.O(gen[2438]),
			.E(gen[2440]),

			.SO(gen[2498]),
			.S(gen[2499]),
			.SE(gen[2500]),

			.SELF(gen[2439]),
			.cell_state(gen[2439])
		); 

/******************* CELL 2440 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2440 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2379]),
			.N(gen[2380]),
			.NE(gen[2381]),

			.O(gen[2439]),
			.E(gen[2441]),

			.SO(gen[2499]),
			.S(gen[2500]),
			.SE(gen[2501]),

			.SELF(gen[2440]),
			.cell_state(gen[2440])
		); 

/******************* CELL 2441 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2441 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2380]),
			.N(gen[2381]),
			.NE(gen[2382]),

			.O(gen[2440]),
			.E(gen[2442]),

			.SO(gen[2500]),
			.S(gen[2501]),
			.SE(gen[2502]),

			.SELF(gen[2441]),
			.cell_state(gen[2441])
		); 

/******************* CELL 2442 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2442 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2381]),
			.N(gen[2382]),
			.NE(gen[2383]),

			.O(gen[2441]),
			.E(gen[2443]),

			.SO(gen[2501]),
			.S(gen[2502]),
			.SE(gen[2503]),

			.SELF(gen[2442]),
			.cell_state(gen[2442])
		); 

/******************* CELL 2443 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2443 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2382]),
			.N(gen[2383]),
			.NE(gen[2384]),

			.O(gen[2442]),
			.E(gen[2444]),

			.SO(gen[2502]),
			.S(gen[2503]),
			.SE(gen[2504]),

			.SELF(gen[2443]),
			.cell_state(gen[2443])
		); 

/******************* CELL 2444 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2444 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2383]),
			.N(gen[2384]),
			.NE(gen[2385]),

			.O(gen[2443]),
			.E(gen[2445]),

			.SO(gen[2503]),
			.S(gen[2504]),
			.SE(gen[2505]),

			.SELF(gen[2444]),
			.cell_state(gen[2444])
		); 

/******************* CELL 2445 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2445 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2384]),
			.N(gen[2385]),
			.NE(gen[2386]),

			.O(gen[2444]),
			.E(gen[2446]),

			.SO(gen[2504]),
			.S(gen[2505]),
			.SE(gen[2506]),

			.SELF(gen[2445]),
			.cell_state(gen[2445])
		); 

/******************* CELL 2446 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2446 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2385]),
			.N(gen[2386]),
			.NE(gen[2387]),

			.O(gen[2445]),
			.E(gen[2447]),

			.SO(gen[2505]),
			.S(gen[2506]),
			.SE(gen[2507]),

			.SELF(gen[2446]),
			.cell_state(gen[2446])
		); 

/******************* CELL 2447 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2447 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2386]),
			.N(gen[2387]),
			.NE(gen[2388]),

			.O(gen[2446]),
			.E(gen[2448]),

			.SO(gen[2506]),
			.S(gen[2507]),
			.SE(gen[2508]),

			.SELF(gen[2447]),
			.cell_state(gen[2447])
		); 

/******************* CELL 2448 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2448 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2387]),
			.N(gen[2388]),
			.NE(gen[2389]),

			.O(gen[2447]),
			.E(gen[2449]),

			.SO(gen[2507]),
			.S(gen[2508]),
			.SE(gen[2509]),

			.SELF(gen[2448]),
			.cell_state(gen[2448])
		); 

/******************* CELL 2449 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2449 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2388]),
			.N(gen[2389]),
			.NE(gen[2390]),

			.O(gen[2448]),
			.E(gen[2450]),

			.SO(gen[2508]),
			.S(gen[2509]),
			.SE(gen[2510]),

			.SELF(gen[2449]),
			.cell_state(gen[2449])
		); 

/******************* CELL 2450 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2450 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2389]),
			.N(gen[2390]),
			.NE(gen[2391]),

			.O(gen[2449]),
			.E(gen[2451]),

			.SO(gen[2509]),
			.S(gen[2510]),
			.SE(gen[2511]),

			.SELF(gen[2450]),
			.cell_state(gen[2450])
		); 

/******************* CELL 2451 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2451 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2390]),
			.N(gen[2391]),
			.NE(gen[2392]),

			.O(gen[2450]),
			.E(gen[2452]),

			.SO(gen[2510]),
			.S(gen[2511]),
			.SE(gen[2512]),

			.SELF(gen[2451]),
			.cell_state(gen[2451])
		); 

/******************* CELL 2452 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2452 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2391]),
			.N(gen[2392]),
			.NE(gen[2393]),

			.O(gen[2451]),
			.E(gen[2453]),

			.SO(gen[2511]),
			.S(gen[2512]),
			.SE(gen[2513]),

			.SELF(gen[2452]),
			.cell_state(gen[2452])
		); 

/******************* CELL 2453 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2453 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2392]),
			.N(gen[2393]),
			.NE(gen[2394]),

			.O(gen[2452]),
			.E(gen[2454]),

			.SO(gen[2512]),
			.S(gen[2513]),
			.SE(gen[2514]),

			.SELF(gen[2453]),
			.cell_state(gen[2453])
		); 

/******************* CELL 2454 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2454 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2393]),
			.N(gen[2394]),
			.NE(gen[2395]),

			.O(gen[2453]),
			.E(gen[2455]),

			.SO(gen[2513]),
			.S(gen[2514]),
			.SE(gen[2515]),

			.SELF(gen[2454]),
			.cell_state(gen[2454])
		); 

/******************* CELL 2455 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2455 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2394]),
			.N(gen[2395]),
			.NE(gen[2396]),

			.O(gen[2454]),
			.E(gen[2456]),

			.SO(gen[2514]),
			.S(gen[2515]),
			.SE(gen[2516]),

			.SELF(gen[2455]),
			.cell_state(gen[2455])
		); 

/******************* CELL 2456 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2456 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2395]),
			.N(gen[2396]),
			.NE(gen[2397]),

			.O(gen[2455]),
			.E(gen[2457]),

			.SO(gen[2515]),
			.S(gen[2516]),
			.SE(gen[2517]),

			.SELF(gen[2456]),
			.cell_state(gen[2456])
		); 

/******************* CELL 2457 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2457 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2396]),
			.N(gen[2397]),
			.NE(gen[2398]),

			.O(gen[2456]),
			.E(gen[2458]),

			.SO(gen[2516]),
			.S(gen[2517]),
			.SE(gen[2518]),

			.SELF(gen[2457]),
			.cell_state(gen[2457])
		); 

/******************* CELL 2458 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2458 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2397]),
			.N(gen[2398]),
			.NE(gen[2399]),

			.O(gen[2457]),
			.E(gen[2459]),

			.SO(gen[2517]),
			.S(gen[2518]),
			.SE(gen[2519]),

			.SELF(gen[2458]),
			.cell_state(gen[2458])
		); 

/******************* CELL 2459 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2459 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2398]),
			.N(gen[2399]),
			.NE(gen[2398]),

			.O(gen[2458]),
			.E(gen[2458]),

			.SO(gen[2518]),
			.S(gen[2519]),
			.SE(gen[2518]),

			.SELF(gen[2459]),
			.cell_state(gen[2459])
		); 

/******************* CELL 2460 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2460 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2401]),
			.N(gen[2400]),
			.NE(gen[2401]),

			.O(gen[2461]),
			.E(gen[2461]),

			.SO(gen[2521]),
			.S(gen[2520]),
			.SE(gen[2521]),

			.SELF(gen[2460]),
			.cell_state(gen[2460])
		); 

/******************* CELL 2461 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2461 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2400]),
			.N(gen[2401]),
			.NE(gen[2402]),

			.O(gen[2460]),
			.E(gen[2462]),

			.SO(gen[2520]),
			.S(gen[2521]),
			.SE(gen[2522]),

			.SELF(gen[2461]),
			.cell_state(gen[2461])
		); 

/******************* CELL 2462 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2462 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2401]),
			.N(gen[2402]),
			.NE(gen[2403]),

			.O(gen[2461]),
			.E(gen[2463]),

			.SO(gen[2521]),
			.S(gen[2522]),
			.SE(gen[2523]),

			.SELF(gen[2462]),
			.cell_state(gen[2462])
		); 

/******************* CELL 2463 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2463 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2402]),
			.N(gen[2403]),
			.NE(gen[2404]),

			.O(gen[2462]),
			.E(gen[2464]),

			.SO(gen[2522]),
			.S(gen[2523]),
			.SE(gen[2524]),

			.SELF(gen[2463]),
			.cell_state(gen[2463])
		); 

/******************* CELL 2464 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2464 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2403]),
			.N(gen[2404]),
			.NE(gen[2405]),

			.O(gen[2463]),
			.E(gen[2465]),

			.SO(gen[2523]),
			.S(gen[2524]),
			.SE(gen[2525]),

			.SELF(gen[2464]),
			.cell_state(gen[2464])
		); 

/******************* CELL 2465 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2465 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2404]),
			.N(gen[2405]),
			.NE(gen[2406]),

			.O(gen[2464]),
			.E(gen[2466]),

			.SO(gen[2524]),
			.S(gen[2525]),
			.SE(gen[2526]),

			.SELF(gen[2465]),
			.cell_state(gen[2465])
		); 

/******************* CELL 2466 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2466 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2405]),
			.N(gen[2406]),
			.NE(gen[2407]),

			.O(gen[2465]),
			.E(gen[2467]),

			.SO(gen[2525]),
			.S(gen[2526]),
			.SE(gen[2527]),

			.SELF(gen[2466]),
			.cell_state(gen[2466])
		); 

/******************* CELL 2467 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2467 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2406]),
			.N(gen[2407]),
			.NE(gen[2408]),

			.O(gen[2466]),
			.E(gen[2468]),

			.SO(gen[2526]),
			.S(gen[2527]),
			.SE(gen[2528]),

			.SELF(gen[2467]),
			.cell_state(gen[2467])
		); 

/******************* CELL 2468 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2468 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2407]),
			.N(gen[2408]),
			.NE(gen[2409]),

			.O(gen[2467]),
			.E(gen[2469]),

			.SO(gen[2527]),
			.S(gen[2528]),
			.SE(gen[2529]),

			.SELF(gen[2468]),
			.cell_state(gen[2468])
		); 

/******************* CELL 2469 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2469 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2408]),
			.N(gen[2409]),
			.NE(gen[2410]),

			.O(gen[2468]),
			.E(gen[2470]),

			.SO(gen[2528]),
			.S(gen[2529]),
			.SE(gen[2530]),

			.SELF(gen[2469]),
			.cell_state(gen[2469])
		); 

/******************* CELL 2470 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2470 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2409]),
			.N(gen[2410]),
			.NE(gen[2411]),

			.O(gen[2469]),
			.E(gen[2471]),

			.SO(gen[2529]),
			.S(gen[2530]),
			.SE(gen[2531]),

			.SELF(gen[2470]),
			.cell_state(gen[2470])
		); 

/******************* CELL 2471 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2471 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2410]),
			.N(gen[2411]),
			.NE(gen[2412]),

			.O(gen[2470]),
			.E(gen[2472]),

			.SO(gen[2530]),
			.S(gen[2531]),
			.SE(gen[2532]),

			.SELF(gen[2471]),
			.cell_state(gen[2471])
		); 

/******************* CELL 2472 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2472 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2411]),
			.N(gen[2412]),
			.NE(gen[2413]),

			.O(gen[2471]),
			.E(gen[2473]),

			.SO(gen[2531]),
			.S(gen[2532]),
			.SE(gen[2533]),

			.SELF(gen[2472]),
			.cell_state(gen[2472])
		); 

/******************* CELL 2473 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2473 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2412]),
			.N(gen[2413]),
			.NE(gen[2414]),

			.O(gen[2472]),
			.E(gen[2474]),

			.SO(gen[2532]),
			.S(gen[2533]),
			.SE(gen[2534]),

			.SELF(gen[2473]),
			.cell_state(gen[2473])
		); 

/******************* CELL 2474 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2474 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2413]),
			.N(gen[2414]),
			.NE(gen[2415]),

			.O(gen[2473]),
			.E(gen[2475]),

			.SO(gen[2533]),
			.S(gen[2534]),
			.SE(gen[2535]),

			.SELF(gen[2474]),
			.cell_state(gen[2474])
		); 

/******************* CELL 2475 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2475 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2414]),
			.N(gen[2415]),
			.NE(gen[2416]),

			.O(gen[2474]),
			.E(gen[2476]),

			.SO(gen[2534]),
			.S(gen[2535]),
			.SE(gen[2536]),

			.SELF(gen[2475]),
			.cell_state(gen[2475])
		); 

/******************* CELL 2476 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2476 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2415]),
			.N(gen[2416]),
			.NE(gen[2417]),

			.O(gen[2475]),
			.E(gen[2477]),

			.SO(gen[2535]),
			.S(gen[2536]),
			.SE(gen[2537]),

			.SELF(gen[2476]),
			.cell_state(gen[2476])
		); 

/******************* CELL 2477 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2477 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2416]),
			.N(gen[2417]),
			.NE(gen[2418]),

			.O(gen[2476]),
			.E(gen[2478]),

			.SO(gen[2536]),
			.S(gen[2537]),
			.SE(gen[2538]),

			.SELF(gen[2477]),
			.cell_state(gen[2477])
		); 

/******************* CELL 2478 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2478 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2417]),
			.N(gen[2418]),
			.NE(gen[2419]),

			.O(gen[2477]),
			.E(gen[2479]),

			.SO(gen[2537]),
			.S(gen[2538]),
			.SE(gen[2539]),

			.SELF(gen[2478]),
			.cell_state(gen[2478])
		); 

/******************* CELL 2479 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2479 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2418]),
			.N(gen[2419]),
			.NE(gen[2420]),

			.O(gen[2478]),
			.E(gen[2480]),

			.SO(gen[2538]),
			.S(gen[2539]),
			.SE(gen[2540]),

			.SELF(gen[2479]),
			.cell_state(gen[2479])
		); 

/******************* CELL 2480 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2480 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2419]),
			.N(gen[2420]),
			.NE(gen[2421]),

			.O(gen[2479]),
			.E(gen[2481]),

			.SO(gen[2539]),
			.S(gen[2540]),
			.SE(gen[2541]),

			.SELF(gen[2480]),
			.cell_state(gen[2480])
		); 

/******************* CELL 2481 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2481 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2420]),
			.N(gen[2421]),
			.NE(gen[2422]),

			.O(gen[2480]),
			.E(gen[2482]),

			.SO(gen[2540]),
			.S(gen[2541]),
			.SE(gen[2542]),

			.SELF(gen[2481]),
			.cell_state(gen[2481])
		); 

/******************* CELL 2482 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2482 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2421]),
			.N(gen[2422]),
			.NE(gen[2423]),

			.O(gen[2481]),
			.E(gen[2483]),

			.SO(gen[2541]),
			.S(gen[2542]),
			.SE(gen[2543]),

			.SELF(gen[2482]),
			.cell_state(gen[2482])
		); 

/******************* CELL 2483 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2483 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2422]),
			.N(gen[2423]),
			.NE(gen[2424]),

			.O(gen[2482]),
			.E(gen[2484]),

			.SO(gen[2542]),
			.S(gen[2543]),
			.SE(gen[2544]),

			.SELF(gen[2483]),
			.cell_state(gen[2483])
		); 

/******************* CELL 2484 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2484 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2423]),
			.N(gen[2424]),
			.NE(gen[2425]),

			.O(gen[2483]),
			.E(gen[2485]),

			.SO(gen[2543]),
			.S(gen[2544]),
			.SE(gen[2545]),

			.SELF(gen[2484]),
			.cell_state(gen[2484])
		); 

/******************* CELL 2485 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2485 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2424]),
			.N(gen[2425]),
			.NE(gen[2426]),

			.O(gen[2484]),
			.E(gen[2486]),

			.SO(gen[2544]),
			.S(gen[2545]),
			.SE(gen[2546]),

			.SELF(gen[2485]),
			.cell_state(gen[2485])
		); 

/******************* CELL 2486 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2486 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2425]),
			.N(gen[2426]),
			.NE(gen[2427]),

			.O(gen[2485]),
			.E(gen[2487]),

			.SO(gen[2545]),
			.S(gen[2546]),
			.SE(gen[2547]),

			.SELF(gen[2486]),
			.cell_state(gen[2486])
		); 

/******************* CELL 2487 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2487 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2426]),
			.N(gen[2427]),
			.NE(gen[2428]),

			.O(gen[2486]),
			.E(gen[2488]),

			.SO(gen[2546]),
			.S(gen[2547]),
			.SE(gen[2548]),

			.SELF(gen[2487]),
			.cell_state(gen[2487])
		); 

/******************* CELL 2488 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2488 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2427]),
			.N(gen[2428]),
			.NE(gen[2429]),

			.O(gen[2487]),
			.E(gen[2489]),

			.SO(gen[2547]),
			.S(gen[2548]),
			.SE(gen[2549]),

			.SELF(gen[2488]),
			.cell_state(gen[2488])
		); 

/******************* CELL 2489 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2489 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2428]),
			.N(gen[2429]),
			.NE(gen[2430]),

			.O(gen[2488]),
			.E(gen[2490]),

			.SO(gen[2548]),
			.S(gen[2549]),
			.SE(gen[2550]),

			.SELF(gen[2489]),
			.cell_state(gen[2489])
		); 

/******************* CELL 2490 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2490 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2429]),
			.N(gen[2430]),
			.NE(gen[2431]),

			.O(gen[2489]),
			.E(gen[2491]),

			.SO(gen[2549]),
			.S(gen[2550]),
			.SE(gen[2551]),

			.SELF(gen[2490]),
			.cell_state(gen[2490])
		); 

/******************* CELL 2491 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2491 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2430]),
			.N(gen[2431]),
			.NE(gen[2432]),

			.O(gen[2490]),
			.E(gen[2492]),

			.SO(gen[2550]),
			.S(gen[2551]),
			.SE(gen[2552]),

			.SELF(gen[2491]),
			.cell_state(gen[2491])
		); 

/******************* CELL 2492 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2492 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2431]),
			.N(gen[2432]),
			.NE(gen[2433]),

			.O(gen[2491]),
			.E(gen[2493]),

			.SO(gen[2551]),
			.S(gen[2552]),
			.SE(gen[2553]),

			.SELF(gen[2492]),
			.cell_state(gen[2492])
		); 

/******************* CELL 2493 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2493 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2432]),
			.N(gen[2433]),
			.NE(gen[2434]),

			.O(gen[2492]),
			.E(gen[2494]),

			.SO(gen[2552]),
			.S(gen[2553]),
			.SE(gen[2554]),

			.SELF(gen[2493]),
			.cell_state(gen[2493])
		); 

/******************* CELL 2494 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2494 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2433]),
			.N(gen[2434]),
			.NE(gen[2435]),

			.O(gen[2493]),
			.E(gen[2495]),

			.SO(gen[2553]),
			.S(gen[2554]),
			.SE(gen[2555]),

			.SELF(gen[2494]),
			.cell_state(gen[2494])
		); 

/******************* CELL 2495 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2495 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2434]),
			.N(gen[2435]),
			.NE(gen[2436]),

			.O(gen[2494]),
			.E(gen[2496]),

			.SO(gen[2554]),
			.S(gen[2555]),
			.SE(gen[2556]),

			.SELF(gen[2495]),
			.cell_state(gen[2495])
		); 

/******************* CELL 2496 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2496 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2435]),
			.N(gen[2436]),
			.NE(gen[2437]),

			.O(gen[2495]),
			.E(gen[2497]),

			.SO(gen[2555]),
			.S(gen[2556]),
			.SE(gen[2557]),

			.SELF(gen[2496]),
			.cell_state(gen[2496])
		); 

/******************* CELL 2497 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2497 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2436]),
			.N(gen[2437]),
			.NE(gen[2438]),

			.O(gen[2496]),
			.E(gen[2498]),

			.SO(gen[2556]),
			.S(gen[2557]),
			.SE(gen[2558]),

			.SELF(gen[2497]),
			.cell_state(gen[2497])
		); 

/******************* CELL 2498 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2498 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2437]),
			.N(gen[2438]),
			.NE(gen[2439]),

			.O(gen[2497]),
			.E(gen[2499]),

			.SO(gen[2557]),
			.S(gen[2558]),
			.SE(gen[2559]),

			.SELF(gen[2498]),
			.cell_state(gen[2498])
		); 

/******************* CELL 2499 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2499 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2438]),
			.N(gen[2439]),
			.NE(gen[2440]),

			.O(gen[2498]),
			.E(gen[2500]),

			.SO(gen[2558]),
			.S(gen[2559]),
			.SE(gen[2560]),

			.SELF(gen[2499]),
			.cell_state(gen[2499])
		); 

/******************* CELL 2500 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2500 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2439]),
			.N(gen[2440]),
			.NE(gen[2441]),

			.O(gen[2499]),
			.E(gen[2501]),

			.SO(gen[2559]),
			.S(gen[2560]),
			.SE(gen[2561]),

			.SELF(gen[2500]),
			.cell_state(gen[2500])
		); 

/******************* CELL 2501 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2501 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2440]),
			.N(gen[2441]),
			.NE(gen[2442]),

			.O(gen[2500]),
			.E(gen[2502]),

			.SO(gen[2560]),
			.S(gen[2561]),
			.SE(gen[2562]),

			.SELF(gen[2501]),
			.cell_state(gen[2501])
		); 

/******************* CELL 2502 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2502 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2441]),
			.N(gen[2442]),
			.NE(gen[2443]),

			.O(gen[2501]),
			.E(gen[2503]),

			.SO(gen[2561]),
			.S(gen[2562]),
			.SE(gen[2563]),

			.SELF(gen[2502]),
			.cell_state(gen[2502])
		); 

/******************* CELL 2503 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2503 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2442]),
			.N(gen[2443]),
			.NE(gen[2444]),

			.O(gen[2502]),
			.E(gen[2504]),

			.SO(gen[2562]),
			.S(gen[2563]),
			.SE(gen[2564]),

			.SELF(gen[2503]),
			.cell_state(gen[2503])
		); 

/******************* CELL 2504 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2504 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2443]),
			.N(gen[2444]),
			.NE(gen[2445]),

			.O(gen[2503]),
			.E(gen[2505]),

			.SO(gen[2563]),
			.S(gen[2564]),
			.SE(gen[2565]),

			.SELF(gen[2504]),
			.cell_state(gen[2504])
		); 

/******************* CELL 2505 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2505 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2444]),
			.N(gen[2445]),
			.NE(gen[2446]),

			.O(gen[2504]),
			.E(gen[2506]),

			.SO(gen[2564]),
			.S(gen[2565]),
			.SE(gen[2566]),

			.SELF(gen[2505]),
			.cell_state(gen[2505])
		); 

/******************* CELL 2506 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2506 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2445]),
			.N(gen[2446]),
			.NE(gen[2447]),

			.O(gen[2505]),
			.E(gen[2507]),

			.SO(gen[2565]),
			.S(gen[2566]),
			.SE(gen[2567]),

			.SELF(gen[2506]),
			.cell_state(gen[2506])
		); 

/******************* CELL 2507 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2507 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2446]),
			.N(gen[2447]),
			.NE(gen[2448]),

			.O(gen[2506]),
			.E(gen[2508]),

			.SO(gen[2566]),
			.S(gen[2567]),
			.SE(gen[2568]),

			.SELF(gen[2507]),
			.cell_state(gen[2507])
		); 

/******************* CELL 2508 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2508 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2447]),
			.N(gen[2448]),
			.NE(gen[2449]),

			.O(gen[2507]),
			.E(gen[2509]),

			.SO(gen[2567]),
			.S(gen[2568]),
			.SE(gen[2569]),

			.SELF(gen[2508]),
			.cell_state(gen[2508])
		); 

/******************* CELL 2509 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2509 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2448]),
			.N(gen[2449]),
			.NE(gen[2450]),

			.O(gen[2508]),
			.E(gen[2510]),

			.SO(gen[2568]),
			.S(gen[2569]),
			.SE(gen[2570]),

			.SELF(gen[2509]),
			.cell_state(gen[2509])
		); 

/******************* CELL 2510 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2510 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2449]),
			.N(gen[2450]),
			.NE(gen[2451]),

			.O(gen[2509]),
			.E(gen[2511]),

			.SO(gen[2569]),
			.S(gen[2570]),
			.SE(gen[2571]),

			.SELF(gen[2510]),
			.cell_state(gen[2510])
		); 

/******************* CELL 2511 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2511 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2450]),
			.N(gen[2451]),
			.NE(gen[2452]),

			.O(gen[2510]),
			.E(gen[2512]),

			.SO(gen[2570]),
			.S(gen[2571]),
			.SE(gen[2572]),

			.SELF(gen[2511]),
			.cell_state(gen[2511])
		); 

/******************* CELL 2512 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2512 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2451]),
			.N(gen[2452]),
			.NE(gen[2453]),

			.O(gen[2511]),
			.E(gen[2513]),

			.SO(gen[2571]),
			.S(gen[2572]),
			.SE(gen[2573]),

			.SELF(gen[2512]),
			.cell_state(gen[2512])
		); 

/******************* CELL 2513 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2513 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2452]),
			.N(gen[2453]),
			.NE(gen[2454]),

			.O(gen[2512]),
			.E(gen[2514]),

			.SO(gen[2572]),
			.S(gen[2573]),
			.SE(gen[2574]),

			.SELF(gen[2513]),
			.cell_state(gen[2513])
		); 

/******************* CELL 2514 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2514 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2453]),
			.N(gen[2454]),
			.NE(gen[2455]),

			.O(gen[2513]),
			.E(gen[2515]),

			.SO(gen[2573]),
			.S(gen[2574]),
			.SE(gen[2575]),

			.SELF(gen[2514]),
			.cell_state(gen[2514])
		); 

/******************* CELL 2515 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2515 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2454]),
			.N(gen[2455]),
			.NE(gen[2456]),

			.O(gen[2514]),
			.E(gen[2516]),

			.SO(gen[2574]),
			.S(gen[2575]),
			.SE(gen[2576]),

			.SELF(gen[2515]),
			.cell_state(gen[2515])
		); 

/******************* CELL 2516 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2516 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2455]),
			.N(gen[2456]),
			.NE(gen[2457]),

			.O(gen[2515]),
			.E(gen[2517]),

			.SO(gen[2575]),
			.S(gen[2576]),
			.SE(gen[2577]),

			.SELF(gen[2516]),
			.cell_state(gen[2516])
		); 

/******************* CELL 2517 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2517 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2456]),
			.N(gen[2457]),
			.NE(gen[2458]),

			.O(gen[2516]),
			.E(gen[2518]),

			.SO(gen[2576]),
			.S(gen[2577]),
			.SE(gen[2578]),

			.SELF(gen[2517]),
			.cell_state(gen[2517])
		); 

/******************* CELL 2518 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2518 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2457]),
			.N(gen[2458]),
			.NE(gen[2459]),

			.O(gen[2517]),
			.E(gen[2519]),

			.SO(gen[2577]),
			.S(gen[2578]),
			.SE(gen[2579]),

			.SELF(gen[2518]),
			.cell_state(gen[2518])
		); 

/******************* CELL 2519 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2519 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2458]),
			.N(gen[2459]),
			.NE(gen[2458]),

			.O(gen[2518]),
			.E(gen[2518]),

			.SO(gen[2578]),
			.S(gen[2579]),
			.SE(gen[2578]),

			.SELF(gen[2519]),
			.cell_state(gen[2519])
		); 

/******************* CELL 2520 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2520 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2461]),
			.N(gen[2460]),
			.NE(gen[2461]),

			.O(gen[2521]),
			.E(gen[2521]),

			.SO(gen[2581]),
			.S(gen[2580]),
			.SE(gen[2581]),

			.SELF(gen[2520]),
			.cell_state(gen[2520])
		); 

/******************* CELL 2521 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2521 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2460]),
			.N(gen[2461]),
			.NE(gen[2462]),

			.O(gen[2520]),
			.E(gen[2522]),

			.SO(gen[2580]),
			.S(gen[2581]),
			.SE(gen[2582]),

			.SELF(gen[2521]),
			.cell_state(gen[2521])
		); 

/******************* CELL 2522 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2522 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2461]),
			.N(gen[2462]),
			.NE(gen[2463]),

			.O(gen[2521]),
			.E(gen[2523]),

			.SO(gen[2581]),
			.S(gen[2582]),
			.SE(gen[2583]),

			.SELF(gen[2522]),
			.cell_state(gen[2522])
		); 

/******************* CELL 2523 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2523 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2462]),
			.N(gen[2463]),
			.NE(gen[2464]),

			.O(gen[2522]),
			.E(gen[2524]),

			.SO(gen[2582]),
			.S(gen[2583]),
			.SE(gen[2584]),

			.SELF(gen[2523]),
			.cell_state(gen[2523])
		); 

/******************* CELL 2524 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2524 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2463]),
			.N(gen[2464]),
			.NE(gen[2465]),

			.O(gen[2523]),
			.E(gen[2525]),

			.SO(gen[2583]),
			.S(gen[2584]),
			.SE(gen[2585]),

			.SELF(gen[2524]),
			.cell_state(gen[2524])
		); 

/******************* CELL 2525 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2525 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2464]),
			.N(gen[2465]),
			.NE(gen[2466]),

			.O(gen[2524]),
			.E(gen[2526]),

			.SO(gen[2584]),
			.S(gen[2585]),
			.SE(gen[2586]),

			.SELF(gen[2525]),
			.cell_state(gen[2525])
		); 

/******************* CELL 2526 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2526 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2465]),
			.N(gen[2466]),
			.NE(gen[2467]),

			.O(gen[2525]),
			.E(gen[2527]),

			.SO(gen[2585]),
			.S(gen[2586]),
			.SE(gen[2587]),

			.SELF(gen[2526]),
			.cell_state(gen[2526])
		); 

/******************* CELL 2527 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2527 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2466]),
			.N(gen[2467]),
			.NE(gen[2468]),

			.O(gen[2526]),
			.E(gen[2528]),

			.SO(gen[2586]),
			.S(gen[2587]),
			.SE(gen[2588]),

			.SELF(gen[2527]),
			.cell_state(gen[2527])
		); 

/******************* CELL 2528 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2528 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2467]),
			.N(gen[2468]),
			.NE(gen[2469]),

			.O(gen[2527]),
			.E(gen[2529]),

			.SO(gen[2587]),
			.S(gen[2588]),
			.SE(gen[2589]),

			.SELF(gen[2528]),
			.cell_state(gen[2528])
		); 

/******************* CELL 2529 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2529 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2468]),
			.N(gen[2469]),
			.NE(gen[2470]),

			.O(gen[2528]),
			.E(gen[2530]),

			.SO(gen[2588]),
			.S(gen[2589]),
			.SE(gen[2590]),

			.SELF(gen[2529]),
			.cell_state(gen[2529])
		); 

/******************* CELL 2530 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2530 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2469]),
			.N(gen[2470]),
			.NE(gen[2471]),

			.O(gen[2529]),
			.E(gen[2531]),

			.SO(gen[2589]),
			.S(gen[2590]),
			.SE(gen[2591]),

			.SELF(gen[2530]),
			.cell_state(gen[2530])
		); 

/******************* CELL 2531 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2531 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2470]),
			.N(gen[2471]),
			.NE(gen[2472]),

			.O(gen[2530]),
			.E(gen[2532]),

			.SO(gen[2590]),
			.S(gen[2591]),
			.SE(gen[2592]),

			.SELF(gen[2531]),
			.cell_state(gen[2531])
		); 

/******************* CELL 2532 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2532 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2471]),
			.N(gen[2472]),
			.NE(gen[2473]),

			.O(gen[2531]),
			.E(gen[2533]),

			.SO(gen[2591]),
			.S(gen[2592]),
			.SE(gen[2593]),

			.SELF(gen[2532]),
			.cell_state(gen[2532])
		); 

/******************* CELL 2533 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2533 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2472]),
			.N(gen[2473]),
			.NE(gen[2474]),

			.O(gen[2532]),
			.E(gen[2534]),

			.SO(gen[2592]),
			.S(gen[2593]),
			.SE(gen[2594]),

			.SELF(gen[2533]),
			.cell_state(gen[2533])
		); 

/******************* CELL 2534 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2534 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2473]),
			.N(gen[2474]),
			.NE(gen[2475]),

			.O(gen[2533]),
			.E(gen[2535]),

			.SO(gen[2593]),
			.S(gen[2594]),
			.SE(gen[2595]),

			.SELF(gen[2534]),
			.cell_state(gen[2534])
		); 

/******************* CELL 2535 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2535 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2474]),
			.N(gen[2475]),
			.NE(gen[2476]),

			.O(gen[2534]),
			.E(gen[2536]),

			.SO(gen[2594]),
			.S(gen[2595]),
			.SE(gen[2596]),

			.SELF(gen[2535]),
			.cell_state(gen[2535])
		); 

/******************* CELL 2536 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2536 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2475]),
			.N(gen[2476]),
			.NE(gen[2477]),

			.O(gen[2535]),
			.E(gen[2537]),

			.SO(gen[2595]),
			.S(gen[2596]),
			.SE(gen[2597]),

			.SELF(gen[2536]),
			.cell_state(gen[2536])
		); 

/******************* CELL 2537 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2537 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2476]),
			.N(gen[2477]),
			.NE(gen[2478]),

			.O(gen[2536]),
			.E(gen[2538]),

			.SO(gen[2596]),
			.S(gen[2597]),
			.SE(gen[2598]),

			.SELF(gen[2537]),
			.cell_state(gen[2537])
		); 

/******************* CELL 2538 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2538 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2477]),
			.N(gen[2478]),
			.NE(gen[2479]),

			.O(gen[2537]),
			.E(gen[2539]),

			.SO(gen[2597]),
			.S(gen[2598]),
			.SE(gen[2599]),

			.SELF(gen[2538]),
			.cell_state(gen[2538])
		); 

/******************* CELL 2539 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2539 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2478]),
			.N(gen[2479]),
			.NE(gen[2480]),

			.O(gen[2538]),
			.E(gen[2540]),

			.SO(gen[2598]),
			.S(gen[2599]),
			.SE(gen[2600]),

			.SELF(gen[2539]),
			.cell_state(gen[2539])
		); 

/******************* CELL 2540 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2540 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2479]),
			.N(gen[2480]),
			.NE(gen[2481]),

			.O(gen[2539]),
			.E(gen[2541]),

			.SO(gen[2599]),
			.S(gen[2600]),
			.SE(gen[2601]),

			.SELF(gen[2540]),
			.cell_state(gen[2540])
		); 

/******************* CELL 2541 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2541 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2480]),
			.N(gen[2481]),
			.NE(gen[2482]),

			.O(gen[2540]),
			.E(gen[2542]),

			.SO(gen[2600]),
			.S(gen[2601]),
			.SE(gen[2602]),

			.SELF(gen[2541]),
			.cell_state(gen[2541])
		); 

/******************* CELL 2542 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2542 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2481]),
			.N(gen[2482]),
			.NE(gen[2483]),

			.O(gen[2541]),
			.E(gen[2543]),

			.SO(gen[2601]),
			.S(gen[2602]),
			.SE(gen[2603]),

			.SELF(gen[2542]),
			.cell_state(gen[2542])
		); 

/******************* CELL 2543 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2543 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2482]),
			.N(gen[2483]),
			.NE(gen[2484]),

			.O(gen[2542]),
			.E(gen[2544]),

			.SO(gen[2602]),
			.S(gen[2603]),
			.SE(gen[2604]),

			.SELF(gen[2543]),
			.cell_state(gen[2543])
		); 

/******************* CELL 2544 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2544 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2483]),
			.N(gen[2484]),
			.NE(gen[2485]),

			.O(gen[2543]),
			.E(gen[2545]),

			.SO(gen[2603]),
			.S(gen[2604]),
			.SE(gen[2605]),

			.SELF(gen[2544]),
			.cell_state(gen[2544])
		); 

/******************* CELL 2545 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2545 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2484]),
			.N(gen[2485]),
			.NE(gen[2486]),

			.O(gen[2544]),
			.E(gen[2546]),

			.SO(gen[2604]),
			.S(gen[2605]),
			.SE(gen[2606]),

			.SELF(gen[2545]),
			.cell_state(gen[2545])
		); 

/******************* CELL 2546 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2546 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2485]),
			.N(gen[2486]),
			.NE(gen[2487]),

			.O(gen[2545]),
			.E(gen[2547]),

			.SO(gen[2605]),
			.S(gen[2606]),
			.SE(gen[2607]),

			.SELF(gen[2546]),
			.cell_state(gen[2546])
		); 

/******************* CELL 2547 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2547 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2486]),
			.N(gen[2487]),
			.NE(gen[2488]),

			.O(gen[2546]),
			.E(gen[2548]),

			.SO(gen[2606]),
			.S(gen[2607]),
			.SE(gen[2608]),

			.SELF(gen[2547]),
			.cell_state(gen[2547])
		); 

/******************* CELL 2548 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2548 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2487]),
			.N(gen[2488]),
			.NE(gen[2489]),

			.O(gen[2547]),
			.E(gen[2549]),

			.SO(gen[2607]),
			.S(gen[2608]),
			.SE(gen[2609]),

			.SELF(gen[2548]),
			.cell_state(gen[2548])
		); 

/******************* CELL 2549 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2549 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2488]),
			.N(gen[2489]),
			.NE(gen[2490]),

			.O(gen[2548]),
			.E(gen[2550]),

			.SO(gen[2608]),
			.S(gen[2609]),
			.SE(gen[2610]),

			.SELF(gen[2549]),
			.cell_state(gen[2549])
		); 

/******************* CELL 2550 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2550 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2489]),
			.N(gen[2490]),
			.NE(gen[2491]),

			.O(gen[2549]),
			.E(gen[2551]),

			.SO(gen[2609]),
			.S(gen[2610]),
			.SE(gen[2611]),

			.SELF(gen[2550]),
			.cell_state(gen[2550])
		); 

/******************* CELL 2551 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2551 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2490]),
			.N(gen[2491]),
			.NE(gen[2492]),

			.O(gen[2550]),
			.E(gen[2552]),

			.SO(gen[2610]),
			.S(gen[2611]),
			.SE(gen[2612]),

			.SELF(gen[2551]),
			.cell_state(gen[2551])
		); 

/******************* CELL 2552 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2552 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2491]),
			.N(gen[2492]),
			.NE(gen[2493]),

			.O(gen[2551]),
			.E(gen[2553]),

			.SO(gen[2611]),
			.S(gen[2612]),
			.SE(gen[2613]),

			.SELF(gen[2552]),
			.cell_state(gen[2552])
		); 

/******************* CELL 2553 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2553 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2492]),
			.N(gen[2493]),
			.NE(gen[2494]),

			.O(gen[2552]),
			.E(gen[2554]),

			.SO(gen[2612]),
			.S(gen[2613]),
			.SE(gen[2614]),

			.SELF(gen[2553]),
			.cell_state(gen[2553])
		); 

/******************* CELL 2554 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2554 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2493]),
			.N(gen[2494]),
			.NE(gen[2495]),

			.O(gen[2553]),
			.E(gen[2555]),

			.SO(gen[2613]),
			.S(gen[2614]),
			.SE(gen[2615]),

			.SELF(gen[2554]),
			.cell_state(gen[2554])
		); 

/******************* CELL 2555 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2555 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2494]),
			.N(gen[2495]),
			.NE(gen[2496]),

			.O(gen[2554]),
			.E(gen[2556]),

			.SO(gen[2614]),
			.S(gen[2615]),
			.SE(gen[2616]),

			.SELF(gen[2555]),
			.cell_state(gen[2555])
		); 

/******************* CELL 2556 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2556 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2495]),
			.N(gen[2496]),
			.NE(gen[2497]),

			.O(gen[2555]),
			.E(gen[2557]),

			.SO(gen[2615]),
			.S(gen[2616]),
			.SE(gen[2617]),

			.SELF(gen[2556]),
			.cell_state(gen[2556])
		); 

/******************* CELL 2557 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2557 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2496]),
			.N(gen[2497]),
			.NE(gen[2498]),

			.O(gen[2556]),
			.E(gen[2558]),

			.SO(gen[2616]),
			.S(gen[2617]),
			.SE(gen[2618]),

			.SELF(gen[2557]),
			.cell_state(gen[2557])
		); 

/******************* CELL 2558 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2558 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2497]),
			.N(gen[2498]),
			.NE(gen[2499]),

			.O(gen[2557]),
			.E(gen[2559]),

			.SO(gen[2617]),
			.S(gen[2618]),
			.SE(gen[2619]),

			.SELF(gen[2558]),
			.cell_state(gen[2558])
		); 

/******************* CELL 2559 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2559 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2498]),
			.N(gen[2499]),
			.NE(gen[2500]),

			.O(gen[2558]),
			.E(gen[2560]),

			.SO(gen[2618]),
			.S(gen[2619]),
			.SE(gen[2620]),

			.SELF(gen[2559]),
			.cell_state(gen[2559])
		); 

/******************* CELL 2560 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2560 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2499]),
			.N(gen[2500]),
			.NE(gen[2501]),

			.O(gen[2559]),
			.E(gen[2561]),

			.SO(gen[2619]),
			.S(gen[2620]),
			.SE(gen[2621]),

			.SELF(gen[2560]),
			.cell_state(gen[2560])
		); 

/******************* CELL 2561 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2561 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2500]),
			.N(gen[2501]),
			.NE(gen[2502]),

			.O(gen[2560]),
			.E(gen[2562]),

			.SO(gen[2620]),
			.S(gen[2621]),
			.SE(gen[2622]),

			.SELF(gen[2561]),
			.cell_state(gen[2561])
		); 

/******************* CELL 2562 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2562 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2501]),
			.N(gen[2502]),
			.NE(gen[2503]),

			.O(gen[2561]),
			.E(gen[2563]),

			.SO(gen[2621]),
			.S(gen[2622]),
			.SE(gen[2623]),

			.SELF(gen[2562]),
			.cell_state(gen[2562])
		); 

/******************* CELL 2563 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2563 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2502]),
			.N(gen[2503]),
			.NE(gen[2504]),

			.O(gen[2562]),
			.E(gen[2564]),

			.SO(gen[2622]),
			.S(gen[2623]),
			.SE(gen[2624]),

			.SELF(gen[2563]),
			.cell_state(gen[2563])
		); 

/******************* CELL 2564 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2564 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2503]),
			.N(gen[2504]),
			.NE(gen[2505]),

			.O(gen[2563]),
			.E(gen[2565]),

			.SO(gen[2623]),
			.S(gen[2624]),
			.SE(gen[2625]),

			.SELF(gen[2564]),
			.cell_state(gen[2564])
		); 

/******************* CELL 2565 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2565 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2504]),
			.N(gen[2505]),
			.NE(gen[2506]),

			.O(gen[2564]),
			.E(gen[2566]),

			.SO(gen[2624]),
			.S(gen[2625]),
			.SE(gen[2626]),

			.SELF(gen[2565]),
			.cell_state(gen[2565])
		); 

/******************* CELL 2566 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2566 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2505]),
			.N(gen[2506]),
			.NE(gen[2507]),

			.O(gen[2565]),
			.E(gen[2567]),

			.SO(gen[2625]),
			.S(gen[2626]),
			.SE(gen[2627]),

			.SELF(gen[2566]),
			.cell_state(gen[2566])
		); 

/******************* CELL 2567 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2567 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2506]),
			.N(gen[2507]),
			.NE(gen[2508]),

			.O(gen[2566]),
			.E(gen[2568]),

			.SO(gen[2626]),
			.S(gen[2627]),
			.SE(gen[2628]),

			.SELF(gen[2567]),
			.cell_state(gen[2567])
		); 

/******************* CELL 2568 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2568 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2507]),
			.N(gen[2508]),
			.NE(gen[2509]),

			.O(gen[2567]),
			.E(gen[2569]),

			.SO(gen[2627]),
			.S(gen[2628]),
			.SE(gen[2629]),

			.SELF(gen[2568]),
			.cell_state(gen[2568])
		); 

/******************* CELL 2569 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2569 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2508]),
			.N(gen[2509]),
			.NE(gen[2510]),

			.O(gen[2568]),
			.E(gen[2570]),

			.SO(gen[2628]),
			.S(gen[2629]),
			.SE(gen[2630]),

			.SELF(gen[2569]),
			.cell_state(gen[2569])
		); 

/******************* CELL 2570 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2570 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2509]),
			.N(gen[2510]),
			.NE(gen[2511]),

			.O(gen[2569]),
			.E(gen[2571]),

			.SO(gen[2629]),
			.S(gen[2630]),
			.SE(gen[2631]),

			.SELF(gen[2570]),
			.cell_state(gen[2570])
		); 

/******************* CELL 2571 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2571 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2510]),
			.N(gen[2511]),
			.NE(gen[2512]),

			.O(gen[2570]),
			.E(gen[2572]),

			.SO(gen[2630]),
			.S(gen[2631]),
			.SE(gen[2632]),

			.SELF(gen[2571]),
			.cell_state(gen[2571])
		); 

/******************* CELL 2572 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2572 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2511]),
			.N(gen[2512]),
			.NE(gen[2513]),

			.O(gen[2571]),
			.E(gen[2573]),

			.SO(gen[2631]),
			.S(gen[2632]),
			.SE(gen[2633]),

			.SELF(gen[2572]),
			.cell_state(gen[2572])
		); 

/******************* CELL 2573 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2573 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2512]),
			.N(gen[2513]),
			.NE(gen[2514]),

			.O(gen[2572]),
			.E(gen[2574]),

			.SO(gen[2632]),
			.S(gen[2633]),
			.SE(gen[2634]),

			.SELF(gen[2573]),
			.cell_state(gen[2573])
		); 

/******************* CELL 2574 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2574 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2513]),
			.N(gen[2514]),
			.NE(gen[2515]),

			.O(gen[2573]),
			.E(gen[2575]),

			.SO(gen[2633]),
			.S(gen[2634]),
			.SE(gen[2635]),

			.SELF(gen[2574]),
			.cell_state(gen[2574])
		); 

/******************* CELL 2575 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2575 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2514]),
			.N(gen[2515]),
			.NE(gen[2516]),

			.O(gen[2574]),
			.E(gen[2576]),

			.SO(gen[2634]),
			.S(gen[2635]),
			.SE(gen[2636]),

			.SELF(gen[2575]),
			.cell_state(gen[2575])
		); 

/******************* CELL 2576 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2576 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2515]),
			.N(gen[2516]),
			.NE(gen[2517]),

			.O(gen[2575]),
			.E(gen[2577]),

			.SO(gen[2635]),
			.S(gen[2636]),
			.SE(gen[2637]),

			.SELF(gen[2576]),
			.cell_state(gen[2576])
		); 

/******************* CELL 2577 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2577 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2516]),
			.N(gen[2517]),
			.NE(gen[2518]),

			.O(gen[2576]),
			.E(gen[2578]),

			.SO(gen[2636]),
			.S(gen[2637]),
			.SE(gen[2638]),

			.SELF(gen[2577]),
			.cell_state(gen[2577])
		); 

/******************* CELL 2578 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2578 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2517]),
			.N(gen[2518]),
			.NE(gen[2519]),

			.O(gen[2577]),
			.E(gen[2579]),

			.SO(gen[2637]),
			.S(gen[2638]),
			.SE(gen[2639]),

			.SELF(gen[2578]),
			.cell_state(gen[2578])
		); 

/******************* CELL 2579 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2579 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2518]),
			.N(gen[2519]),
			.NE(gen[2518]),

			.O(gen[2578]),
			.E(gen[2578]),

			.SO(gen[2638]),
			.S(gen[2639]),
			.SE(gen[2638]),

			.SELF(gen[2579]),
			.cell_state(gen[2579])
		); 

/******************* CELL 2580 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2580 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2521]),
			.N(gen[2520]),
			.NE(gen[2521]),

			.O(gen[2581]),
			.E(gen[2581]),

			.SO(gen[2641]),
			.S(gen[2640]),
			.SE(gen[2641]),

			.SELF(gen[2580]),
			.cell_state(gen[2580])
		); 

/******************* CELL 2581 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2581 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2520]),
			.N(gen[2521]),
			.NE(gen[2522]),

			.O(gen[2580]),
			.E(gen[2582]),

			.SO(gen[2640]),
			.S(gen[2641]),
			.SE(gen[2642]),

			.SELF(gen[2581]),
			.cell_state(gen[2581])
		); 

/******************* CELL 2582 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2582 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2521]),
			.N(gen[2522]),
			.NE(gen[2523]),

			.O(gen[2581]),
			.E(gen[2583]),

			.SO(gen[2641]),
			.S(gen[2642]),
			.SE(gen[2643]),

			.SELF(gen[2582]),
			.cell_state(gen[2582])
		); 

/******************* CELL 2583 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2583 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2522]),
			.N(gen[2523]),
			.NE(gen[2524]),

			.O(gen[2582]),
			.E(gen[2584]),

			.SO(gen[2642]),
			.S(gen[2643]),
			.SE(gen[2644]),

			.SELF(gen[2583]),
			.cell_state(gen[2583])
		); 

/******************* CELL 2584 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2584 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2523]),
			.N(gen[2524]),
			.NE(gen[2525]),

			.O(gen[2583]),
			.E(gen[2585]),

			.SO(gen[2643]),
			.S(gen[2644]),
			.SE(gen[2645]),

			.SELF(gen[2584]),
			.cell_state(gen[2584])
		); 

/******************* CELL 2585 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2585 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2524]),
			.N(gen[2525]),
			.NE(gen[2526]),

			.O(gen[2584]),
			.E(gen[2586]),

			.SO(gen[2644]),
			.S(gen[2645]),
			.SE(gen[2646]),

			.SELF(gen[2585]),
			.cell_state(gen[2585])
		); 

/******************* CELL 2586 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2586 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2525]),
			.N(gen[2526]),
			.NE(gen[2527]),

			.O(gen[2585]),
			.E(gen[2587]),

			.SO(gen[2645]),
			.S(gen[2646]),
			.SE(gen[2647]),

			.SELF(gen[2586]),
			.cell_state(gen[2586])
		); 

/******************* CELL 2587 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2587 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2526]),
			.N(gen[2527]),
			.NE(gen[2528]),

			.O(gen[2586]),
			.E(gen[2588]),

			.SO(gen[2646]),
			.S(gen[2647]),
			.SE(gen[2648]),

			.SELF(gen[2587]),
			.cell_state(gen[2587])
		); 

/******************* CELL 2588 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2588 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2527]),
			.N(gen[2528]),
			.NE(gen[2529]),

			.O(gen[2587]),
			.E(gen[2589]),

			.SO(gen[2647]),
			.S(gen[2648]),
			.SE(gen[2649]),

			.SELF(gen[2588]),
			.cell_state(gen[2588])
		); 

/******************* CELL 2589 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2589 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2528]),
			.N(gen[2529]),
			.NE(gen[2530]),

			.O(gen[2588]),
			.E(gen[2590]),

			.SO(gen[2648]),
			.S(gen[2649]),
			.SE(gen[2650]),

			.SELF(gen[2589]),
			.cell_state(gen[2589])
		); 

/******************* CELL 2590 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2590 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2529]),
			.N(gen[2530]),
			.NE(gen[2531]),

			.O(gen[2589]),
			.E(gen[2591]),

			.SO(gen[2649]),
			.S(gen[2650]),
			.SE(gen[2651]),

			.SELF(gen[2590]),
			.cell_state(gen[2590])
		); 

/******************* CELL 2591 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2591 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2530]),
			.N(gen[2531]),
			.NE(gen[2532]),

			.O(gen[2590]),
			.E(gen[2592]),

			.SO(gen[2650]),
			.S(gen[2651]),
			.SE(gen[2652]),

			.SELF(gen[2591]),
			.cell_state(gen[2591])
		); 

/******************* CELL 2592 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2592 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2531]),
			.N(gen[2532]),
			.NE(gen[2533]),

			.O(gen[2591]),
			.E(gen[2593]),

			.SO(gen[2651]),
			.S(gen[2652]),
			.SE(gen[2653]),

			.SELF(gen[2592]),
			.cell_state(gen[2592])
		); 

/******************* CELL 2593 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2593 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2532]),
			.N(gen[2533]),
			.NE(gen[2534]),

			.O(gen[2592]),
			.E(gen[2594]),

			.SO(gen[2652]),
			.S(gen[2653]),
			.SE(gen[2654]),

			.SELF(gen[2593]),
			.cell_state(gen[2593])
		); 

/******************* CELL 2594 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2594 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2533]),
			.N(gen[2534]),
			.NE(gen[2535]),

			.O(gen[2593]),
			.E(gen[2595]),

			.SO(gen[2653]),
			.S(gen[2654]),
			.SE(gen[2655]),

			.SELF(gen[2594]),
			.cell_state(gen[2594])
		); 

/******************* CELL 2595 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2595 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2534]),
			.N(gen[2535]),
			.NE(gen[2536]),

			.O(gen[2594]),
			.E(gen[2596]),

			.SO(gen[2654]),
			.S(gen[2655]),
			.SE(gen[2656]),

			.SELF(gen[2595]),
			.cell_state(gen[2595])
		); 

/******************* CELL 2596 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2596 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2535]),
			.N(gen[2536]),
			.NE(gen[2537]),

			.O(gen[2595]),
			.E(gen[2597]),

			.SO(gen[2655]),
			.S(gen[2656]),
			.SE(gen[2657]),

			.SELF(gen[2596]),
			.cell_state(gen[2596])
		); 

/******************* CELL 2597 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2597 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2536]),
			.N(gen[2537]),
			.NE(gen[2538]),

			.O(gen[2596]),
			.E(gen[2598]),

			.SO(gen[2656]),
			.S(gen[2657]),
			.SE(gen[2658]),

			.SELF(gen[2597]),
			.cell_state(gen[2597])
		); 

/******************* CELL 2598 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2598 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2537]),
			.N(gen[2538]),
			.NE(gen[2539]),

			.O(gen[2597]),
			.E(gen[2599]),

			.SO(gen[2657]),
			.S(gen[2658]),
			.SE(gen[2659]),

			.SELF(gen[2598]),
			.cell_state(gen[2598])
		); 

/******************* CELL 2599 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2599 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2538]),
			.N(gen[2539]),
			.NE(gen[2540]),

			.O(gen[2598]),
			.E(gen[2600]),

			.SO(gen[2658]),
			.S(gen[2659]),
			.SE(gen[2660]),

			.SELF(gen[2599]),
			.cell_state(gen[2599])
		); 

/******************* CELL 2600 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2600 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2539]),
			.N(gen[2540]),
			.NE(gen[2541]),

			.O(gen[2599]),
			.E(gen[2601]),

			.SO(gen[2659]),
			.S(gen[2660]),
			.SE(gen[2661]),

			.SELF(gen[2600]),
			.cell_state(gen[2600])
		); 

/******************* CELL 2601 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2601 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2540]),
			.N(gen[2541]),
			.NE(gen[2542]),

			.O(gen[2600]),
			.E(gen[2602]),

			.SO(gen[2660]),
			.S(gen[2661]),
			.SE(gen[2662]),

			.SELF(gen[2601]),
			.cell_state(gen[2601])
		); 

/******************* CELL 2602 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2602 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2541]),
			.N(gen[2542]),
			.NE(gen[2543]),

			.O(gen[2601]),
			.E(gen[2603]),

			.SO(gen[2661]),
			.S(gen[2662]),
			.SE(gen[2663]),

			.SELF(gen[2602]),
			.cell_state(gen[2602])
		); 

/******************* CELL 2603 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2603 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2542]),
			.N(gen[2543]),
			.NE(gen[2544]),

			.O(gen[2602]),
			.E(gen[2604]),

			.SO(gen[2662]),
			.S(gen[2663]),
			.SE(gen[2664]),

			.SELF(gen[2603]),
			.cell_state(gen[2603])
		); 

/******************* CELL 2604 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2604 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2543]),
			.N(gen[2544]),
			.NE(gen[2545]),

			.O(gen[2603]),
			.E(gen[2605]),

			.SO(gen[2663]),
			.S(gen[2664]),
			.SE(gen[2665]),

			.SELF(gen[2604]),
			.cell_state(gen[2604])
		); 

/******************* CELL 2605 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2605 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2544]),
			.N(gen[2545]),
			.NE(gen[2546]),

			.O(gen[2604]),
			.E(gen[2606]),

			.SO(gen[2664]),
			.S(gen[2665]),
			.SE(gen[2666]),

			.SELF(gen[2605]),
			.cell_state(gen[2605])
		); 

/******************* CELL 2606 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2606 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2545]),
			.N(gen[2546]),
			.NE(gen[2547]),

			.O(gen[2605]),
			.E(gen[2607]),

			.SO(gen[2665]),
			.S(gen[2666]),
			.SE(gen[2667]),

			.SELF(gen[2606]),
			.cell_state(gen[2606])
		); 

/******************* CELL 2607 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2607 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2546]),
			.N(gen[2547]),
			.NE(gen[2548]),

			.O(gen[2606]),
			.E(gen[2608]),

			.SO(gen[2666]),
			.S(gen[2667]),
			.SE(gen[2668]),

			.SELF(gen[2607]),
			.cell_state(gen[2607])
		); 

/******************* CELL 2608 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2608 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2547]),
			.N(gen[2548]),
			.NE(gen[2549]),

			.O(gen[2607]),
			.E(gen[2609]),

			.SO(gen[2667]),
			.S(gen[2668]),
			.SE(gen[2669]),

			.SELF(gen[2608]),
			.cell_state(gen[2608])
		); 

/******************* CELL 2609 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2609 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2548]),
			.N(gen[2549]),
			.NE(gen[2550]),

			.O(gen[2608]),
			.E(gen[2610]),

			.SO(gen[2668]),
			.S(gen[2669]),
			.SE(gen[2670]),

			.SELF(gen[2609]),
			.cell_state(gen[2609])
		); 

/******************* CELL 2610 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2610 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2549]),
			.N(gen[2550]),
			.NE(gen[2551]),

			.O(gen[2609]),
			.E(gen[2611]),

			.SO(gen[2669]),
			.S(gen[2670]),
			.SE(gen[2671]),

			.SELF(gen[2610]),
			.cell_state(gen[2610])
		); 

/******************* CELL 2611 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2611 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2550]),
			.N(gen[2551]),
			.NE(gen[2552]),

			.O(gen[2610]),
			.E(gen[2612]),

			.SO(gen[2670]),
			.S(gen[2671]),
			.SE(gen[2672]),

			.SELF(gen[2611]),
			.cell_state(gen[2611])
		); 

/******************* CELL 2612 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2612 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2551]),
			.N(gen[2552]),
			.NE(gen[2553]),

			.O(gen[2611]),
			.E(gen[2613]),

			.SO(gen[2671]),
			.S(gen[2672]),
			.SE(gen[2673]),

			.SELF(gen[2612]),
			.cell_state(gen[2612])
		); 

/******************* CELL 2613 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2613 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2552]),
			.N(gen[2553]),
			.NE(gen[2554]),

			.O(gen[2612]),
			.E(gen[2614]),

			.SO(gen[2672]),
			.S(gen[2673]),
			.SE(gen[2674]),

			.SELF(gen[2613]),
			.cell_state(gen[2613])
		); 

/******************* CELL 2614 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2614 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2553]),
			.N(gen[2554]),
			.NE(gen[2555]),

			.O(gen[2613]),
			.E(gen[2615]),

			.SO(gen[2673]),
			.S(gen[2674]),
			.SE(gen[2675]),

			.SELF(gen[2614]),
			.cell_state(gen[2614])
		); 

/******************* CELL 2615 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2615 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2554]),
			.N(gen[2555]),
			.NE(gen[2556]),

			.O(gen[2614]),
			.E(gen[2616]),

			.SO(gen[2674]),
			.S(gen[2675]),
			.SE(gen[2676]),

			.SELF(gen[2615]),
			.cell_state(gen[2615])
		); 

/******************* CELL 2616 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2616 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2555]),
			.N(gen[2556]),
			.NE(gen[2557]),

			.O(gen[2615]),
			.E(gen[2617]),

			.SO(gen[2675]),
			.S(gen[2676]),
			.SE(gen[2677]),

			.SELF(gen[2616]),
			.cell_state(gen[2616])
		); 

/******************* CELL 2617 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2617 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2556]),
			.N(gen[2557]),
			.NE(gen[2558]),

			.O(gen[2616]),
			.E(gen[2618]),

			.SO(gen[2676]),
			.S(gen[2677]),
			.SE(gen[2678]),

			.SELF(gen[2617]),
			.cell_state(gen[2617])
		); 

/******************* CELL 2618 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2618 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2557]),
			.N(gen[2558]),
			.NE(gen[2559]),

			.O(gen[2617]),
			.E(gen[2619]),

			.SO(gen[2677]),
			.S(gen[2678]),
			.SE(gen[2679]),

			.SELF(gen[2618]),
			.cell_state(gen[2618])
		); 

/******************* CELL 2619 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2619 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2558]),
			.N(gen[2559]),
			.NE(gen[2560]),

			.O(gen[2618]),
			.E(gen[2620]),

			.SO(gen[2678]),
			.S(gen[2679]),
			.SE(gen[2680]),

			.SELF(gen[2619]),
			.cell_state(gen[2619])
		); 

/******************* CELL 2620 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2620 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2559]),
			.N(gen[2560]),
			.NE(gen[2561]),

			.O(gen[2619]),
			.E(gen[2621]),

			.SO(gen[2679]),
			.S(gen[2680]),
			.SE(gen[2681]),

			.SELF(gen[2620]),
			.cell_state(gen[2620])
		); 

/******************* CELL 2621 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2621 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2560]),
			.N(gen[2561]),
			.NE(gen[2562]),

			.O(gen[2620]),
			.E(gen[2622]),

			.SO(gen[2680]),
			.S(gen[2681]),
			.SE(gen[2682]),

			.SELF(gen[2621]),
			.cell_state(gen[2621])
		); 

/******************* CELL 2622 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2622 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2561]),
			.N(gen[2562]),
			.NE(gen[2563]),

			.O(gen[2621]),
			.E(gen[2623]),

			.SO(gen[2681]),
			.S(gen[2682]),
			.SE(gen[2683]),

			.SELF(gen[2622]),
			.cell_state(gen[2622])
		); 

/******************* CELL 2623 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2623 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2562]),
			.N(gen[2563]),
			.NE(gen[2564]),

			.O(gen[2622]),
			.E(gen[2624]),

			.SO(gen[2682]),
			.S(gen[2683]),
			.SE(gen[2684]),

			.SELF(gen[2623]),
			.cell_state(gen[2623])
		); 

/******************* CELL 2624 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2624 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2563]),
			.N(gen[2564]),
			.NE(gen[2565]),

			.O(gen[2623]),
			.E(gen[2625]),

			.SO(gen[2683]),
			.S(gen[2684]),
			.SE(gen[2685]),

			.SELF(gen[2624]),
			.cell_state(gen[2624])
		); 

/******************* CELL 2625 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2625 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2564]),
			.N(gen[2565]),
			.NE(gen[2566]),

			.O(gen[2624]),
			.E(gen[2626]),

			.SO(gen[2684]),
			.S(gen[2685]),
			.SE(gen[2686]),

			.SELF(gen[2625]),
			.cell_state(gen[2625])
		); 

/******************* CELL 2626 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2626 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2565]),
			.N(gen[2566]),
			.NE(gen[2567]),

			.O(gen[2625]),
			.E(gen[2627]),

			.SO(gen[2685]),
			.S(gen[2686]),
			.SE(gen[2687]),

			.SELF(gen[2626]),
			.cell_state(gen[2626])
		); 

/******************* CELL 2627 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2627 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2566]),
			.N(gen[2567]),
			.NE(gen[2568]),

			.O(gen[2626]),
			.E(gen[2628]),

			.SO(gen[2686]),
			.S(gen[2687]),
			.SE(gen[2688]),

			.SELF(gen[2627]),
			.cell_state(gen[2627])
		); 

/******************* CELL 2628 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2628 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2567]),
			.N(gen[2568]),
			.NE(gen[2569]),

			.O(gen[2627]),
			.E(gen[2629]),

			.SO(gen[2687]),
			.S(gen[2688]),
			.SE(gen[2689]),

			.SELF(gen[2628]),
			.cell_state(gen[2628])
		); 

/******************* CELL 2629 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2629 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2568]),
			.N(gen[2569]),
			.NE(gen[2570]),

			.O(gen[2628]),
			.E(gen[2630]),

			.SO(gen[2688]),
			.S(gen[2689]),
			.SE(gen[2690]),

			.SELF(gen[2629]),
			.cell_state(gen[2629])
		); 

/******************* CELL 2630 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2630 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2569]),
			.N(gen[2570]),
			.NE(gen[2571]),

			.O(gen[2629]),
			.E(gen[2631]),

			.SO(gen[2689]),
			.S(gen[2690]),
			.SE(gen[2691]),

			.SELF(gen[2630]),
			.cell_state(gen[2630])
		); 

/******************* CELL 2631 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2631 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2570]),
			.N(gen[2571]),
			.NE(gen[2572]),

			.O(gen[2630]),
			.E(gen[2632]),

			.SO(gen[2690]),
			.S(gen[2691]),
			.SE(gen[2692]),

			.SELF(gen[2631]),
			.cell_state(gen[2631])
		); 

/******************* CELL 2632 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2632 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2571]),
			.N(gen[2572]),
			.NE(gen[2573]),

			.O(gen[2631]),
			.E(gen[2633]),

			.SO(gen[2691]),
			.S(gen[2692]),
			.SE(gen[2693]),

			.SELF(gen[2632]),
			.cell_state(gen[2632])
		); 

/******************* CELL 2633 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2633 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2572]),
			.N(gen[2573]),
			.NE(gen[2574]),

			.O(gen[2632]),
			.E(gen[2634]),

			.SO(gen[2692]),
			.S(gen[2693]),
			.SE(gen[2694]),

			.SELF(gen[2633]),
			.cell_state(gen[2633])
		); 

/******************* CELL 2634 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2634 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2573]),
			.N(gen[2574]),
			.NE(gen[2575]),

			.O(gen[2633]),
			.E(gen[2635]),

			.SO(gen[2693]),
			.S(gen[2694]),
			.SE(gen[2695]),

			.SELF(gen[2634]),
			.cell_state(gen[2634])
		); 

/******************* CELL 2635 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2635 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2574]),
			.N(gen[2575]),
			.NE(gen[2576]),

			.O(gen[2634]),
			.E(gen[2636]),

			.SO(gen[2694]),
			.S(gen[2695]),
			.SE(gen[2696]),

			.SELF(gen[2635]),
			.cell_state(gen[2635])
		); 

/******************* CELL 2636 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2636 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2575]),
			.N(gen[2576]),
			.NE(gen[2577]),

			.O(gen[2635]),
			.E(gen[2637]),

			.SO(gen[2695]),
			.S(gen[2696]),
			.SE(gen[2697]),

			.SELF(gen[2636]),
			.cell_state(gen[2636])
		); 

/******************* CELL 2637 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2637 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2576]),
			.N(gen[2577]),
			.NE(gen[2578]),

			.O(gen[2636]),
			.E(gen[2638]),

			.SO(gen[2696]),
			.S(gen[2697]),
			.SE(gen[2698]),

			.SELF(gen[2637]),
			.cell_state(gen[2637])
		); 

/******************* CELL 2638 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2638 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2577]),
			.N(gen[2578]),
			.NE(gen[2579]),

			.O(gen[2637]),
			.E(gen[2639]),

			.SO(gen[2697]),
			.S(gen[2698]),
			.SE(gen[2699]),

			.SELF(gen[2638]),
			.cell_state(gen[2638])
		); 

/******************* CELL 2639 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2639 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2578]),
			.N(gen[2579]),
			.NE(gen[2578]),

			.O(gen[2638]),
			.E(gen[2638]),

			.SO(gen[2698]),
			.S(gen[2699]),
			.SE(gen[2698]),

			.SELF(gen[2639]),
			.cell_state(gen[2639])
		); 

/******************* CELL 2640 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2640 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2581]),
			.N(gen[2580]),
			.NE(gen[2581]),

			.O(gen[2641]),
			.E(gen[2641]),

			.SO(gen[2701]),
			.S(gen[2700]),
			.SE(gen[2701]),

			.SELF(gen[2640]),
			.cell_state(gen[2640])
		); 

/******************* CELL 2641 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2641 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2580]),
			.N(gen[2581]),
			.NE(gen[2582]),

			.O(gen[2640]),
			.E(gen[2642]),

			.SO(gen[2700]),
			.S(gen[2701]),
			.SE(gen[2702]),

			.SELF(gen[2641]),
			.cell_state(gen[2641])
		); 

/******************* CELL 2642 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2642 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2581]),
			.N(gen[2582]),
			.NE(gen[2583]),

			.O(gen[2641]),
			.E(gen[2643]),

			.SO(gen[2701]),
			.S(gen[2702]),
			.SE(gen[2703]),

			.SELF(gen[2642]),
			.cell_state(gen[2642])
		); 

/******************* CELL 2643 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2643 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2582]),
			.N(gen[2583]),
			.NE(gen[2584]),

			.O(gen[2642]),
			.E(gen[2644]),

			.SO(gen[2702]),
			.S(gen[2703]),
			.SE(gen[2704]),

			.SELF(gen[2643]),
			.cell_state(gen[2643])
		); 

/******************* CELL 2644 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2644 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2583]),
			.N(gen[2584]),
			.NE(gen[2585]),

			.O(gen[2643]),
			.E(gen[2645]),

			.SO(gen[2703]),
			.S(gen[2704]),
			.SE(gen[2705]),

			.SELF(gen[2644]),
			.cell_state(gen[2644])
		); 

/******************* CELL 2645 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2645 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2584]),
			.N(gen[2585]),
			.NE(gen[2586]),

			.O(gen[2644]),
			.E(gen[2646]),

			.SO(gen[2704]),
			.S(gen[2705]),
			.SE(gen[2706]),

			.SELF(gen[2645]),
			.cell_state(gen[2645])
		); 

/******************* CELL 2646 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2646 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2585]),
			.N(gen[2586]),
			.NE(gen[2587]),

			.O(gen[2645]),
			.E(gen[2647]),

			.SO(gen[2705]),
			.S(gen[2706]),
			.SE(gen[2707]),

			.SELF(gen[2646]),
			.cell_state(gen[2646])
		); 

/******************* CELL 2647 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2647 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2586]),
			.N(gen[2587]),
			.NE(gen[2588]),

			.O(gen[2646]),
			.E(gen[2648]),

			.SO(gen[2706]),
			.S(gen[2707]),
			.SE(gen[2708]),

			.SELF(gen[2647]),
			.cell_state(gen[2647])
		); 

/******************* CELL 2648 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2648 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2587]),
			.N(gen[2588]),
			.NE(gen[2589]),

			.O(gen[2647]),
			.E(gen[2649]),

			.SO(gen[2707]),
			.S(gen[2708]),
			.SE(gen[2709]),

			.SELF(gen[2648]),
			.cell_state(gen[2648])
		); 

/******************* CELL 2649 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2649 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2588]),
			.N(gen[2589]),
			.NE(gen[2590]),

			.O(gen[2648]),
			.E(gen[2650]),

			.SO(gen[2708]),
			.S(gen[2709]),
			.SE(gen[2710]),

			.SELF(gen[2649]),
			.cell_state(gen[2649])
		); 

/******************* CELL 2650 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2650 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2589]),
			.N(gen[2590]),
			.NE(gen[2591]),

			.O(gen[2649]),
			.E(gen[2651]),

			.SO(gen[2709]),
			.S(gen[2710]),
			.SE(gen[2711]),

			.SELF(gen[2650]),
			.cell_state(gen[2650])
		); 

/******************* CELL 2651 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2651 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2590]),
			.N(gen[2591]),
			.NE(gen[2592]),

			.O(gen[2650]),
			.E(gen[2652]),

			.SO(gen[2710]),
			.S(gen[2711]),
			.SE(gen[2712]),

			.SELF(gen[2651]),
			.cell_state(gen[2651])
		); 

/******************* CELL 2652 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2652 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2591]),
			.N(gen[2592]),
			.NE(gen[2593]),

			.O(gen[2651]),
			.E(gen[2653]),

			.SO(gen[2711]),
			.S(gen[2712]),
			.SE(gen[2713]),

			.SELF(gen[2652]),
			.cell_state(gen[2652])
		); 

/******************* CELL 2653 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2653 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2592]),
			.N(gen[2593]),
			.NE(gen[2594]),

			.O(gen[2652]),
			.E(gen[2654]),

			.SO(gen[2712]),
			.S(gen[2713]),
			.SE(gen[2714]),

			.SELF(gen[2653]),
			.cell_state(gen[2653])
		); 

/******************* CELL 2654 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2654 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2593]),
			.N(gen[2594]),
			.NE(gen[2595]),

			.O(gen[2653]),
			.E(gen[2655]),

			.SO(gen[2713]),
			.S(gen[2714]),
			.SE(gen[2715]),

			.SELF(gen[2654]),
			.cell_state(gen[2654])
		); 

/******************* CELL 2655 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2655 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2594]),
			.N(gen[2595]),
			.NE(gen[2596]),

			.O(gen[2654]),
			.E(gen[2656]),

			.SO(gen[2714]),
			.S(gen[2715]),
			.SE(gen[2716]),

			.SELF(gen[2655]),
			.cell_state(gen[2655])
		); 

/******************* CELL 2656 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2656 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2595]),
			.N(gen[2596]),
			.NE(gen[2597]),

			.O(gen[2655]),
			.E(gen[2657]),

			.SO(gen[2715]),
			.S(gen[2716]),
			.SE(gen[2717]),

			.SELF(gen[2656]),
			.cell_state(gen[2656])
		); 

/******************* CELL 2657 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2657 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2596]),
			.N(gen[2597]),
			.NE(gen[2598]),

			.O(gen[2656]),
			.E(gen[2658]),

			.SO(gen[2716]),
			.S(gen[2717]),
			.SE(gen[2718]),

			.SELF(gen[2657]),
			.cell_state(gen[2657])
		); 

/******************* CELL 2658 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2658 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2597]),
			.N(gen[2598]),
			.NE(gen[2599]),

			.O(gen[2657]),
			.E(gen[2659]),

			.SO(gen[2717]),
			.S(gen[2718]),
			.SE(gen[2719]),

			.SELF(gen[2658]),
			.cell_state(gen[2658])
		); 

/******************* CELL 2659 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2659 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2598]),
			.N(gen[2599]),
			.NE(gen[2600]),

			.O(gen[2658]),
			.E(gen[2660]),

			.SO(gen[2718]),
			.S(gen[2719]),
			.SE(gen[2720]),

			.SELF(gen[2659]),
			.cell_state(gen[2659])
		); 

/******************* CELL 2660 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2660 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2599]),
			.N(gen[2600]),
			.NE(gen[2601]),

			.O(gen[2659]),
			.E(gen[2661]),

			.SO(gen[2719]),
			.S(gen[2720]),
			.SE(gen[2721]),

			.SELF(gen[2660]),
			.cell_state(gen[2660])
		); 

/******************* CELL 2661 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2661 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2600]),
			.N(gen[2601]),
			.NE(gen[2602]),

			.O(gen[2660]),
			.E(gen[2662]),

			.SO(gen[2720]),
			.S(gen[2721]),
			.SE(gen[2722]),

			.SELF(gen[2661]),
			.cell_state(gen[2661])
		); 

/******************* CELL 2662 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2662 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2601]),
			.N(gen[2602]),
			.NE(gen[2603]),

			.O(gen[2661]),
			.E(gen[2663]),

			.SO(gen[2721]),
			.S(gen[2722]),
			.SE(gen[2723]),

			.SELF(gen[2662]),
			.cell_state(gen[2662])
		); 

/******************* CELL 2663 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2663 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2602]),
			.N(gen[2603]),
			.NE(gen[2604]),

			.O(gen[2662]),
			.E(gen[2664]),

			.SO(gen[2722]),
			.S(gen[2723]),
			.SE(gen[2724]),

			.SELF(gen[2663]),
			.cell_state(gen[2663])
		); 

/******************* CELL 2664 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2664 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2603]),
			.N(gen[2604]),
			.NE(gen[2605]),

			.O(gen[2663]),
			.E(gen[2665]),

			.SO(gen[2723]),
			.S(gen[2724]),
			.SE(gen[2725]),

			.SELF(gen[2664]),
			.cell_state(gen[2664])
		); 

/******************* CELL 2665 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2665 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2604]),
			.N(gen[2605]),
			.NE(gen[2606]),

			.O(gen[2664]),
			.E(gen[2666]),

			.SO(gen[2724]),
			.S(gen[2725]),
			.SE(gen[2726]),

			.SELF(gen[2665]),
			.cell_state(gen[2665])
		); 

/******************* CELL 2666 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2666 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2605]),
			.N(gen[2606]),
			.NE(gen[2607]),

			.O(gen[2665]),
			.E(gen[2667]),

			.SO(gen[2725]),
			.S(gen[2726]),
			.SE(gen[2727]),

			.SELF(gen[2666]),
			.cell_state(gen[2666])
		); 

/******************* CELL 2667 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2667 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2606]),
			.N(gen[2607]),
			.NE(gen[2608]),

			.O(gen[2666]),
			.E(gen[2668]),

			.SO(gen[2726]),
			.S(gen[2727]),
			.SE(gen[2728]),

			.SELF(gen[2667]),
			.cell_state(gen[2667])
		); 

/******************* CELL 2668 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2668 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2607]),
			.N(gen[2608]),
			.NE(gen[2609]),

			.O(gen[2667]),
			.E(gen[2669]),

			.SO(gen[2727]),
			.S(gen[2728]),
			.SE(gen[2729]),

			.SELF(gen[2668]),
			.cell_state(gen[2668])
		); 

/******************* CELL 2669 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2669 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2608]),
			.N(gen[2609]),
			.NE(gen[2610]),

			.O(gen[2668]),
			.E(gen[2670]),

			.SO(gen[2728]),
			.S(gen[2729]),
			.SE(gen[2730]),

			.SELF(gen[2669]),
			.cell_state(gen[2669])
		); 

/******************* CELL 2670 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2670 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2609]),
			.N(gen[2610]),
			.NE(gen[2611]),

			.O(gen[2669]),
			.E(gen[2671]),

			.SO(gen[2729]),
			.S(gen[2730]),
			.SE(gen[2731]),

			.SELF(gen[2670]),
			.cell_state(gen[2670])
		); 

/******************* CELL 2671 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2671 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2610]),
			.N(gen[2611]),
			.NE(gen[2612]),

			.O(gen[2670]),
			.E(gen[2672]),

			.SO(gen[2730]),
			.S(gen[2731]),
			.SE(gen[2732]),

			.SELF(gen[2671]),
			.cell_state(gen[2671])
		); 

/******************* CELL 2672 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2672 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2611]),
			.N(gen[2612]),
			.NE(gen[2613]),

			.O(gen[2671]),
			.E(gen[2673]),

			.SO(gen[2731]),
			.S(gen[2732]),
			.SE(gen[2733]),

			.SELF(gen[2672]),
			.cell_state(gen[2672])
		); 

/******************* CELL 2673 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2673 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2612]),
			.N(gen[2613]),
			.NE(gen[2614]),

			.O(gen[2672]),
			.E(gen[2674]),

			.SO(gen[2732]),
			.S(gen[2733]),
			.SE(gen[2734]),

			.SELF(gen[2673]),
			.cell_state(gen[2673])
		); 

/******************* CELL 2674 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2674 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2613]),
			.N(gen[2614]),
			.NE(gen[2615]),

			.O(gen[2673]),
			.E(gen[2675]),

			.SO(gen[2733]),
			.S(gen[2734]),
			.SE(gen[2735]),

			.SELF(gen[2674]),
			.cell_state(gen[2674])
		); 

/******************* CELL 2675 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2675 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2614]),
			.N(gen[2615]),
			.NE(gen[2616]),

			.O(gen[2674]),
			.E(gen[2676]),

			.SO(gen[2734]),
			.S(gen[2735]),
			.SE(gen[2736]),

			.SELF(gen[2675]),
			.cell_state(gen[2675])
		); 

/******************* CELL 2676 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2676 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2615]),
			.N(gen[2616]),
			.NE(gen[2617]),

			.O(gen[2675]),
			.E(gen[2677]),

			.SO(gen[2735]),
			.S(gen[2736]),
			.SE(gen[2737]),

			.SELF(gen[2676]),
			.cell_state(gen[2676])
		); 

/******************* CELL 2677 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2677 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2616]),
			.N(gen[2617]),
			.NE(gen[2618]),

			.O(gen[2676]),
			.E(gen[2678]),

			.SO(gen[2736]),
			.S(gen[2737]),
			.SE(gen[2738]),

			.SELF(gen[2677]),
			.cell_state(gen[2677])
		); 

/******************* CELL 2678 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2678 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2617]),
			.N(gen[2618]),
			.NE(gen[2619]),

			.O(gen[2677]),
			.E(gen[2679]),

			.SO(gen[2737]),
			.S(gen[2738]),
			.SE(gen[2739]),

			.SELF(gen[2678]),
			.cell_state(gen[2678])
		); 

/******************* CELL 2679 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2679 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2618]),
			.N(gen[2619]),
			.NE(gen[2620]),

			.O(gen[2678]),
			.E(gen[2680]),

			.SO(gen[2738]),
			.S(gen[2739]),
			.SE(gen[2740]),

			.SELF(gen[2679]),
			.cell_state(gen[2679])
		); 

/******************* CELL 2680 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2680 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2619]),
			.N(gen[2620]),
			.NE(gen[2621]),

			.O(gen[2679]),
			.E(gen[2681]),

			.SO(gen[2739]),
			.S(gen[2740]),
			.SE(gen[2741]),

			.SELF(gen[2680]),
			.cell_state(gen[2680])
		); 

/******************* CELL 2681 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2681 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2620]),
			.N(gen[2621]),
			.NE(gen[2622]),

			.O(gen[2680]),
			.E(gen[2682]),

			.SO(gen[2740]),
			.S(gen[2741]),
			.SE(gen[2742]),

			.SELF(gen[2681]),
			.cell_state(gen[2681])
		); 

/******************* CELL 2682 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2682 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2621]),
			.N(gen[2622]),
			.NE(gen[2623]),

			.O(gen[2681]),
			.E(gen[2683]),

			.SO(gen[2741]),
			.S(gen[2742]),
			.SE(gen[2743]),

			.SELF(gen[2682]),
			.cell_state(gen[2682])
		); 

/******************* CELL 2683 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2683 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2622]),
			.N(gen[2623]),
			.NE(gen[2624]),

			.O(gen[2682]),
			.E(gen[2684]),

			.SO(gen[2742]),
			.S(gen[2743]),
			.SE(gen[2744]),

			.SELF(gen[2683]),
			.cell_state(gen[2683])
		); 

/******************* CELL 2684 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2684 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2623]),
			.N(gen[2624]),
			.NE(gen[2625]),

			.O(gen[2683]),
			.E(gen[2685]),

			.SO(gen[2743]),
			.S(gen[2744]),
			.SE(gen[2745]),

			.SELF(gen[2684]),
			.cell_state(gen[2684])
		); 

/******************* CELL 2685 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2685 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2624]),
			.N(gen[2625]),
			.NE(gen[2626]),

			.O(gen[2684]),
			.E(gen[2686]),

			.SO(gen[2744]),
			.S(gen[2745]),
			.SE(gen[2746]),

			.SELF(gen[2685]),
			.cell_state(gen[2685])
		); 

/******************* CELL 2686 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2686 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2625]),
			.N(gen[2626]),
			.NE(gen[2627]),

			.O(gen[2685]),
			.E(gen[2687]),

			.SO(gen[2745]),
			.S(gen[2746]),
			.SE(gen[2747]),

			.SELF(gen[2686]),
			.cell_state(gen[2686])
		); 

/******************* CELL 2687 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2687 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2626]),
			.N(gen[2627]),
			.NE(gen[2628]),

			.O(gen[2686]),
			.E(gen[2688]),

			.SO(gen[2746]),
			.S(gen[2747]),
			.SE(gen[2748]),

			.SELF(gen[2687]),
			.cell_state(gen[2687])
		); 

/******************* CELL 2688 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2688 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2627]),
			.N(gen[2628]),
			.NE(gen[2629]),

			.O(gen[2687]),
			.E(gen[2689]),

			.SO(gen[2747]),
			.S(gen[2748]),
			.SE(gen[2749]),

			.SELF(gen[2688]),
			.cell_state(gen[2688])
		); 

/******************* CELL 2689 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2689 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2628]),
			.N(gen[2629]),
			.NE(gen[2630]),

			.O(gen[2688]),
			.E(gen[2690]),

			.SO(gen[2748]),
			.S(gen[2749]),
			.SE(gen[2750]),

			.SELF(gen[2689]),
			.cell_state(gen[2689])
		); 

/******************* CELL 2690 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2690 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2629]),
			.N(gen[2630]),
			.NE(gen[2631]),

			.O(gen[2689]),
			.E(gen[2691]),

			.SO(gen[2749]),
			.S(gen[2750]),
			.SE(gen[2751]),

			.SELF(gen[2690]),
			.cell_state(gen[2690])
		); 

/******************* CELL 2691 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2691 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2630]),
			.N(gen[2631]),
			.NE(gen[2632]),

			.O(gen[2690]),
			.E(gen[2692]),

			.SO(gen[2750]),
			.S(gen[2751]),
			.SE(gen[2752]),

			.SELF(gen[2691]),
			.cell_state(gen[2691])
		); 

/******************* CELL 2692 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2692 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2631]),
			.N(gen[2632]),
			.NE(gen[2633]),

			.O(gen[2691]),
			.E(gen[2693]),

			.SO(gen[2751]),
			.S(gen[2752]),
			.SE(gen[2753]),

			.SELF(gen[2692]),
			.cell_state(gen[2692])
		); 

/******************* CELL 2693 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2693 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2632]),
			.N(gen[2633]),
			.NE(gen[2634]),

			.O(gen[2692]),
			.E(gen[2694]),

			.SO(gen[2752]),
			.S(gen[2753]),
			.SE(gen[2754]),

			.SELF(gen[2693]),
			.cell_state(gen[2693])
		); 

/******************* CELL 2694 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2694 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2633]),
			.N(gen[2634]),
			.NE(gen[2635]),

			.O(gen[2693]),
			.E(gen[2695]),

			.SO(gen[2753]),
			.S(gen[2754]),
			.SE(gen[2755]),

			.SELF(gen[2694]),
			.cell_state(gen[2694])
		); 

/******************* CELL 2695 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2695 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2634]),
			.N(gen[2635]),
			.NE(gen[2636]),

			.O(gen[2694]),
			.E(gen[2696]),

			.SO(gen[2754]),
			.S(gen[2755]),
			.SE(gen[2756]),

			.SELF(gen[2695]),
			.cell_state(gen[2695])
		); 

/******************* CELL 2696 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2696 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2635]),
			.N(gen[2636]),
			.NE(gen[2637]),

			.O(gen[2695]),
			.E(gen[2697]),

			.SO(gen[2755]),
			.S(gen[2756]),
			.SE(gen[2757]),

			.SELF(gen[2696]),
			.cell_state(gen[2696])
		); 

/******************* CELL 2697 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2697 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2636]),
			.N(gen[2637]),
			.NE(gen[2638]),

			.O(gen[2696]),
			.E(gen[2698]),

			.SO(gen[2756]),
			.S(gen[2757]),
			.SE(gen[2758]),

			.SELF(gen[2697]),
			.cell_state(gen[2697])
		); 

/******************* CELL 2698 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2698 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2637]),
			.N(gen[2638]),
			.NE(gen[2639]),

			.O(gen[2697]),
			.E(gen[2699]),

			.SO(gen[2757]),
			.S(gen[2758]),
			.SE(gen[2759]),

			.SELF(gen[2698]),
			.cell_state(gen[2698])
		); 

/******************* CELL 2699 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2699 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2638]),
			.N(gen[2639]),
			.NE(gen[2638]),

			.O(gen[2698]),
			.E(gen[2698]),

			.SO(gen[2758]),
			.S(gen[2759]),
			.SE(gen[2758]),

			.SELF(gen[2699]),
			.cell_state(gen[2699])
		); 

/******************* CELL 2700 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2700 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2641]),
			.N(gen[2640]),
			.NE(gen[2641]),

			.O(gen[2701]),
			.E(gen[2701]),

			.SO(gen[2761]),
			.S(gen[2760]),
			.SE(gen[2761]),

			.SELF(gen[2700]),
			.cell_state(gen[2700])
		); 

/******************* CELL 2701 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2701 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2640]),
			.N(gen[2641]),
			.NE(gen[2642]),

			.O(gen[2700]),
			.E(gen[2702]),

			.SO(gen[2760]),
			.S(gen[2761]),
			.SE(gen[2762]),

			.SELF(gen[2701]),
			.cell_state(gen[2701])
		); 

/******************* CELL 2702 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2702 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2641]),
			.N(gen[2642]),
			.NE(gen[2643]),

			.O(gen[2701]),
			.E(gen[2703]),

			.SO(gen[2761]),
			.S(gen[2762]),
			.SE(gen[2763]),

			.SELF(gen[2702]),
			.cell_state(gen[2702])
		); 

/******************* CELL 2703 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2703 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2642]),
			.N(gen[2643]),
			.NE(gen[2644]),

			.O(gen[2702]),
			.E(gen[2704]),

			.SO(gen[2762]),
			.S(gen[2763]),
			.SE(gen[2764]),

			.SELF(gen[2703]),
			.cell_state(gen[2703])
		); 

/******************* CELL 2704 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2704 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2643]),
			.N(gen[2644]),
			.NE(gen[2645]),

			.O(gen[2703]),
			.E(gen[2705]),

			.SO(gen[2763]),
			.S(gen[2764]),
			.SE(gen[2765]),

			.SELF(gen[2704]),
			.cell_state(gen[2704])
		); 

/******************* CELL 2705 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2705 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2644]),
			.N(gen[2645]),
			.NE(gen[2646]),

			.O(gen[2704]),
			.E(gen[2706]),

			.SO(gen[2764]),
			.S(gen[2765]),
			.SE(gen[2766]),

			.SELF(gen[2705]),
			.cell_state(gen[2705])
		); 

/******************* CELL 2706 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2706 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2645]),
			.N(gen[2646]),
			.NE(gen[2647]),

			.O(gen[2705]),
			.E(gen[2707]),

			.SO(gen[2765]),
			.S(gen[2766]),
			.SE(gen[2767]),

			.SELF(gen[2706]),
			.cell_state(gen[2706])
		); 

/******************* CELL 2707 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2707 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2646]),
			.N(gen[2647]),
			.NE(gen[2648]),

			.O(gen[2706]),
			.E(gen[2708]),

			.SO(gen[2766]),
			.S(gen[2767]),
			.SE(gen[2768]),

			.SELF(gen[2707]),
			.cell_state(gen[2707])
		); 

/******************* CELL 2708 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2708 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2647]),
			.N(gen[2648]),
			.NE(gen[2649]),

			.O(gen[2707]),
			.E(gen[2709]),

			.SO(gen[2767]),
			.S(gen[2768]),
			.SE(gen[2769]),

			.SELF(gen[2708]),
			.cell_state(gen[2708])
		); 

/******************* CELL 2709 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2709 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2648]),
			.N(gen[2649]),
			.NE(gen[2650]),

			.O(gen[2708]),
			.E(gen[2710]),

			.SO(gen[2768]),
			.S(gen[2769]),
			.SE(gen[2770]),

			.SELF(gen[2709]),
			.cell_state(gen[2709])
		); 

/******************* CELL 2710 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2710 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2649]),
			.N(gen[2650]),
			.NE(gen[2651]),

			.O(gen[2709]),
			.E(gen[2711]),

			.SO(gen[2769]),
			.S(gen[2770]),
			.SE(gen[2771]),

			.SELF(gen[2710]),
			.cell_state(gen[2710])
		); 

/******************* CELL 2711 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2711 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2650]),
			.N(gen[2651]),
			.NE(gen[2652]),

			.O(gen[2710]),
			.E(gen[2712]),

			.SO(gen[2770]),
			.S(gen[2771]),
			.SE(gen[2772]),

			.SELF(gen[2711]),
			.cell_state(gen[2711])
		); 

/******************* CELL 2712 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2712 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2651]),
			.N(gen[2652]),
			.NE(gen[2653]),

			.O(gen[2711]),
			.E(gen[2713]),

			.SO(gen[2771]),
			.S(gen[2772]),
			.SE(gen[2773]),

			.SELF(gen[2712]),
			.cell_state(gen[2712])
		); 

/******************* CELL 2713 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2713 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2652]),
			.N(gen[2653]),
			.NE(gen[2654]),

			.O(gen[2712]),
			.E(gen[2714]),

			.SO(gen[2772]),
			.S(gen[2773]),
			.SE(gen[2774]),

			.SELF(gen[2713]),
			.cell_state(gen[2713])
		); 

/******************* CELL 2714 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2714 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2653]),
			.N(gen[2654]),
			.NE(gen[2655]),

			.O(gen[2713]),
			.E(gen[2715]),

			.SO(gen[2773]),
			.S(gen[2774]),
			.SE(gen[2775]),

			.SELF(gen[2714]),
			.cell_state(gen[2714])
		); 

/******************* CELL 2715 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2715 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2654]),
			.N(gen[2655]),
			.NE(gen[2656]),

			.O(gen[2714]),
			.E(gen[2716]),

			.SO(gen[2774]),
			.S(gen[2775]),
			.SE(gen[2776]),

			.SELF(gen[2715]),
			.cell_state(gen[2715])
		); 

/******************* CELL 2716 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2716 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2655]),
			.N(gen[2656]),
			.NE(gen[2657]),

			.O(gen[2715]),
			.E(gen[2717]),

			.SO(gen[2775]),
			.S(gen[2776]),
			.SE(gen[2777]),

			.SELF(gen[2716]),
			.cell_state(gen[2716])
		); 

/******************* CELL 2717 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2717 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2656]),
			.N(gen[2657]),
			.NE(gen[2658]),

			.O(gen[2716]),
			.E(gen[2718]),

			.SO(gen[2776]),
			.S(gen[2777]),
			.SE(gen[2778]),

			.SELF(gen[2717]),
			.cell_state(gen[2717])
		); 

/******************* CELL 2718 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2718 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2657]),
			.N(gen[2658]),
			.NE(gen[2659]),

			.O(gen[2717]),
			.E(gen[2719]),

			.SO(gen[2777]),
			.S(gen[2778]),
			.SE(gen[2779]),

			.SELF(gen[2718]),
			.cell_state(gen[2718])
		); 

/******************* CELL 2719 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2719 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2658]),
			.N(gen[2659]),
			.NE(gen[2660]),

			.O(gen[2718]),
			.E(gen[2720]),

			.SO(gen[2778]),
			.S(gen[2779]),
			.SE(gen[2780]),

			.SELF(gen[2719]),
			.cell_state(gen[2719])
		); 

/******************* CELL 2720 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2720 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2659]),
			.N(gen[2660]),
			.NE(gen[2661]),

			.O(gen[2719]),
			.E(gen[2721]),

			.SO(gen[2779]),
			.S(gen[2780]),
			.SE(gen[2781]),

			.SELF(gen[2720]),
			.cell_state(gen[2720])
		); 

/******************* CELL 2721 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2721 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2660]),
			.N(gen[2661]),
			.NE(gen[2662]),

			.O(gen[2720]),
			.E(gen[2722]),

			.SO(gen[2780]),
			.S(gen[2781]),
			.SE(gen[2782]),

			.SELF(gen[2721]),
			.cell_state(gen[2721])
		); 

/******************* CELL 2722 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2722 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2661]),
			.N(gen[2662]),
			.NE(gen[2663]),

			.O(gen[2721]),
			.E(gen[2723]),

			.SO(gen[2781]),
			.S(gen[2782]),
			.SE(gen[2783]),

			.SELF(gen[2722]),
			.cell_state(gen[2722])
		); 

/******************* CELL 2723 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2723 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2662]),
			.N(gen[2663]),
			.NE(gen[2664]),

			.O(gen[2722]),
			.E(gen[2724]),

			.SO(gen[2782]),
			.S(gen[2783]),
			.SE(gen[2784]),

			.SELF(gen[2723]),
			.cell_state(gen[2723])
		); 

/******************* CELL 2724 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2724 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2663]),
			.N(gen[2664]),
			.NE(gen[2665]),

			.O(gen[2723]),
			.E(gen[2725]),

			.SO(gen[2783]),
			.S(gen[2784]),
			.SE(gen[2785]),

			.SELF(gen[2724]),
			.cell_state(gen[2724])
		); 

/******************* CELL 2725 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2725 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2664]),
			.N(gen[2665]),
			.NE(gen[2666]),

			.O(gen[2724]),
			.E(gen[2726]),

			.SO(gen[2784]),
			.S(gen[2785]),
			.SE(gen[2786]),

			.SELF(gen[2725]),
			.cell_state(gen[2725])
		); 

/******************* CELL 2726 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2726 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2665]),
			.N(gen[2666]),
			.NE(gen[2667]),

			.O(gen[2725]),
			.E(gen[2727]),

			.SO(gen[2785]),
			.S(gen[2786]),
			.SE(gen[2787]),

			.SELF(gen[2726]),
			.cell_state(gen[2726])
		); 

/******************* CELL 2727 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2727 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2666]),
			.N(gen[2667]),
			.NE(gen[2668]),

			.O(gen[2726]),
			.E(gen[2728]),

			.SO(gen[2786]),
			.S(gen[2787]),
			.SE(gen[2788]),

			.SELF(gen[2727]),
			.cell_state(gen[2727])
		); 

/******************* CELL 2728 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2728 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2667]),
			.N(gen[2668]),
			.NE(gen[2669]),

			.O(gen[2727]),
			.E(gen[2729]),

			.SO(gen[2787]),
			.S(gen[2788]),
			.SE(gen[2789]),

			.SELF(gen[2728]),
			.cell_state(gen[2728])
		); 

/******************* CELL 2729 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2729 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2668]),
			.N(gen[2669]),
			.NE(gen[2670]),

			.O(gen[2728]),
			.E(gen[2730]),

			.SO(gen[2788]),
			.S(gen[2789]),
			.SE(gen[2790]),

			.SELF(gen[2729]),
			.cell_state(gen[2729])
		); 

/******************* CELL 2730 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2730 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2669]),
			.N(gen[2670]),
			.NE(gen[2671]),

			.O(gen[2729]),
			.E(gen[2731]),

			.SO(gen[2789]),
			.S(gen[2790]),
			.SE(gen[2791]),

			.SELF(gen[2730]),
			.cell_state(gen[2730])
		); 

/******************* CELL 2731 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2731 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2670]),
			.N(gen[2671]),
			.NE(gen[2672]),

			.O(gen[2730]),
			.E(gen[2732]),

			.SO(gen[2790]),
			.S(gen[2791]),
			.SE(gen[2792]),

			.SELF(gen[2731]),
			.cell_state(gen[2731])
		); 

/******************* CELL 2732 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2732 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2671]),
			.N(gen[2672]),
			.NE(gen[2673]),

			.O(gen[2731]),
			.E(gen[2733]),

			.SO(gen[2791]),
			.S(gen[2792]),
			.SE(gen[2793]),

			.SELF(gen[2732]),
			.cell_state(gen[2732])
		); 

/******************* CELL 2733 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2733 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2672]),
			.N(gen[2673]),
			.NE(gen[2674]),

			.O(gen[2732]),
			.E(gen[2734]),

			.SO(gen[2792]),
			.S(gen[2793]),
			.SE(gen[2794]),

			.SELF(gen[2733]),
			.cell_state(gen[2733])
		); 

/******************* CELL 2734 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2734 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2673]),
			.N(gen[2674]),
			.NE(gen[2675]),

			.O(gen[2733]),
			.E(gen[2735]),

			.SO(gen[2793]),
			.S(gen[2794]),
			.SE(gen[2795]),

			.SELF(gen[2734]),
			.cell_state(gen[2734])
		); 

/******************* CELL 2735 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2735 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2674]),
			.N(gen[2675]),
			.NE(gen[2676]),

			.O(gen[2734]),
			.E(gen[2736]),

			.SO(gen[2794]),
			.S(gen[2795]),
			.SE(gen[2796]),

			.SELF(gen[2735]),
			.cell_state(gen[2735])
		); 

/******************* CELL 2736 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2736 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2675]),
			.N(gen[2676]),
			.NE(gen[2677]),

			.O(gen[2735]),
			.E(gen[2737]),

			.SO(gen[2795]),
			.S(gen[2796]),
			.SE(gen[2797]),

			.SELF(gen[2736]),
			.cell_state(gen[2736])
		); 

/******************* CELL 2737 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2737 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2676]),
			.N(gen[2677]),
			.NE(gen[2678]),

			.O(gen[2736]),
			.E(gen[2738]),

			.SO(gen[2796]),
			.S(gen[2797]),
			.SE(gen[2798]),

			.SELF(gen[2737]),
			.cell_state(gen[2737])
		); 

/******************* CELL 2738 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2738 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2677]),
			.N(gen[2678]),
			.NE(gen[2679]),

			.O(gen[2737]),
			.E(gen[2739]),

			.SO(gen[2797]),
			.S(gen[2798]),
			.SE(gen[2799]),

			.SELF(gen[2738]),
			.cell_state(gen[2738])
		); 

/******************* CELL 2739 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2739 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2678]),
			.N(gen[2679]),
			.NE(gen[2680]),

			.O(gen[2738]),
			.E(gen[2740]),

			.SO(gen[2798]),
			.S(gen[2799]),
			.SE(gen[2800]),

			.SELF(gen[2739]),
			.cell_state(gen[2739])
		); 

/******************* CELL 2740 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2740 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2679]),
			.N(gen[2680]),
			.NE(gen[2681]),

			.O(gen[2739]),
			.E(gen[2741]),

			.SO(gen[2799]),
			.S(gen[2800]),
			.SE(gen[2801]),

			.SELF(gen[2740]),
			.cell_state(gen[2740])
		); 

/******************* CELL 2741 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2741 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2680]),
			.N(gen[2681]),
			.NE(gen[2682]),

			.O(gen[2740]),
			.E(gen[2742]),

			.SO(gen[2800]),
			.S(gen[2801]),
			.SE(gen[2802]),

			.SELF(gen[2741]),
			.cell_state(gen[2741])
		); 

/******************* CELL 2742 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2742 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2681]),
			.N(gen[2682]),
			.NE(gen[2683]),

			.O(gen[2741]),
			.E(gen[2743]),

			.SO(gen[2801]),
			.S(gen[2802]),
			.SE(gen[2803]),

			.SELF(gen[2742]),
			.cell_state(gen[2742])
		); 

/******************* CELL 2743 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2743 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2682]),
			.N(gen[2683]),
			.NE(gen[2684]),

			.O(gen[2742]),
			.E(gen[2744]),

			.SO(gen[2802]),
			.S(gen[2803]),
			.SE(gen[2804]),

			.SELF(gen[2743]),
			.cell_state(gen[2743])
		); 

/******************* CELL 2744 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2744 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2683]),
			.N(gen[2684]),
			.NE(gen[2685]),

			.O(gen[2743]),
			.E(gen[2745]),

			.SO(gen[2803]),
			.S(gen[2804]),
			.SE(gen[2805]),

			.SELF(gen[2744]),
			.cell_state(gen[2744])
		); 

/******************* CELL 2745 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2745 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2684]),
			.N(gen[2685]),
			.NE(gen[2686]),

			.O(gen[2744]),
			.E(gen[2746]),

			.SO(gen[2804]),
			.S(gen[2805]),
			.SE(gen[2806]),

			.SELF(gen[2745]),
			.cell_state(gen[2745])
		); 

/******************* CELL 2746 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2746 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2685]),
			.N(gen[2686]),
			.NE(gen[2687]),

			.O(gen[2745]),
			.E(gen[2747]),

			.SO(gen[2805]),
			.S(gen[2806]),
			.SE(gen[2807]),

			.SELF(gen[2746]),
			.cell_state(gen[2746])
		); 

/******************* CELL 2747 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2747 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2686]),
			.N(gen[2687]),
			.NE(gen[2688]),

			.O(gen[2746]),
			.E(gen[2748]),

			.SO(gen[2806]),
			.S(gen[2807]),
			.SE(gen[2808]),

			.SELF(gen[2747]),
			.cell_state(gen[2747])
		); 

/******************* CELL 2748 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2748 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2687]),
			.N(gen[2688]),
			.NE(gen[2689]),

			.O(gen[2747]),
			.E(gen[2749]),

			.SO(gen[2807]),
			.S(gen[2808]),
			.SE(gen[2809]),

			.SELF(gen[2748]),
			.cell_state(gen[2748])
		); 

/******************* CELL 2749 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2749 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2688]),
			.N(gen[2689]),
			.NE(gen[2690]),

			.O(gen[2748]),
			.E(gen[2750]),

			.SO(gen[2808]),
			.S(gen[2809]),
			.SE(gen[2810]),

			.SELF(gen[2749]),
			.cell_state(gen[2749])
		); 

/******************* CELL 2750 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2750 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2689]),
			.N(gen[2690]),
			.NE(gen[2691]),

			.O(gen[2749]),
			.E(gen[2751]),

			.SO(gen[2809]),
			.S(gen[2810]),
			.SE(gen[2811]),

			.SELF(gen[2750]),
			.cell_state(gen[2750])
		); 

/******************* CELL 2751 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2751 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2690]),
			.N(gen[2691]),
			.NE(gen[2692]),

			.O(gen[2750]),
			.E(gen[2752]),

			.SO(gen[2810]),
			.S(gen[2811]),
			.SE(gen[2812]),

			.SELF(gen[2751]),
			.cell_state(gen[2751])
		); 

/******************* CELL 2752 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2752 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2691]),
			.N(gen[2692]),
			.NE(gen[2693]),

			.O(gen[2751]),
			.E(gen[2753]),

			.SO(gen[2811]),
			.S(gen[2812]),
			.SE(gen[2813]),

			.SELF(gen[2752]),
			.cell_state(gen[2752])
		); 

/******************* CELL 2753 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2753 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2692]),
			.N(gen[2693]),
			.NE(gen[2694]),

			.O(gen[2752]),
			.E(gen[2754]),

			.SO(gen[2812]),
			.S(gen[2813]),
			.SE(gen[2814]),

			.SELF(gen[2753]),
			.cell_state(gen[2753])
		); 

/******************* CELL 2754 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2754 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2693]),
			.N(gen[2694]),
			.NE(gen[2695]),

			.O(gen[2753]),
			.E(gen[2755]),

			.SO(gen[2813]),
			.S(gen[2814]),
			.SE(gen[2815]),

			.SELF(gen[2754]),
			.cell_state(gen[2754])
		); 

/******************* CELL 2755 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2755 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2694]),
			.N(gen[2695]),
			.NE(gen[2696]),

			.O(gen[2754]),
			.E(gen[2756]),

			.SO(gen[2814]),
			.S(gen[2815]),
			.SE(gen[2816]),

			.SELF(gen[2755]),
			.cell_state(gen[2755])
		); 

/******************* CELL 2756 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2756 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2695]),
			.N(gen[2696]),
			.NE(gen[2697]),

			.O(gen[2755]),
			.E(gen[2757]),

			.SO(gen[2815]),
			.S(gen[2816]),
			.SE(gen[2817]),

			.SELF(gen[2756]),
			.cell_state(gen[2756])
		); 

/******************* CELL 2757 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2757 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2696]),
			.N(gen[2697]),
			.NE(gen[2698]),

			.O(gen[2756]),
			.E(gen[2758]),

			.SO(gen[2816]),
			.S(gen[2817]),
			.SE(gen[2818]),

			.SELF(gen[2757]),
			.cell_state(gen[2757])
		); 

/******************* CELL 2758 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2758 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2697]),
			.N(gen[2698]),
			.NE(gen[2699]),

			.O(gen[2757]),
			.E(gen[2759]),

			.SO(gen[2817]),
			.S(gen[2818]),
			.SE(gen[2819]),

			.SELF(gen[2758]),
			.cell_state(gen[2758])
		); 

/******************* CELL 2759 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2759 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2698]),
			.N(gen[2699]),
			.NE(gen[2698]),

			.O(gen[2758]),
			.E(gen[2758]),

			.SO(gen[2818]),
			.S(gen[2819]),
			.SE(gen[2818]),

			.SELF(gen[2759]),
			.cell_state(gen[2759])
		); 

/******************* CELL 2760 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2760 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2701]),
			.N(gen[2700]),
			.NE(gen[2701]),

			.O(gen[2761]),
			.E(gen[2761]),

			.SO(gen[2821]),
			.S(gen[2820]),
			.SE(gen[2821]),

			.SELF(gen[2760]),
			.cell_state(gen[2760])
		); 

/******************* CELL 2761 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2761 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2700]),
			.N(gen[2701]),
			.NE(gen[2702]),

			.O(gen[2760]),
			.E(gen[2762]),

			.SO(gen[2820]),
			.S(gen[2821]),
			.SE(gen[2822]),

			.SELF(gen[2761]),
			.cell_state(gen[2761])
		); 

/******************* CELL 2762 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2762 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2701]),
			.N(gen[2702]),
			.NE(gen[2703]),

			.O(gen[2761]),
			.E(gen[2763]),

			.SO(gen[2821]),
			.S(gen[2822]),
			.SE(gen[2823]),

			.SELF(gen[2762]),
			.cell_state(gen[2762])
		); 

/******************* CELL 2763 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2763 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2702]),
			.N(gen[2703]),
			.NE(gen[2704]),

			.O(gen[2762]),
			.E(gen[2764]),

			.SO(gen[2822]),
			.S(gen[2823]),
			.SE(gen[2824]),

			.SELF(gen[2763]),
			.cell_state(gen[2763])
		); 

/******************* CELL 2764 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2764 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2703]),
			.N(gen[2704]),
			.NE(gen[2705]),

			.O(gen[2763]),
			.E(gen[2765]),

			.SO(gen[2823]),
			.S(gen[2824]),
			.SE(gen[2825]),

			.SELF(gen[2764]),
			.cell_state(gen[2764])
		); 

/******************* CELL 2765 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2765 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2704]),
			.N(gen[2705]),
			.NE(gen[2706]),

			.O(gen[2764]),
			.E(gen[2766]),

			.SO(gen[2824]),
			.S(gen[2825]),
			.SE(gen[2826]),

			.SELF(gen[2765]),
			.cell_state(gen[2765])
		); 

/******************* CELL 2766 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2766 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2705]),
			.N(gen[2706]),
			.NE(gen[2707]),

			.O(gen[2765]),
			.E(gen[2767]),

			.SO(gen[2825]),
			.S(gen[2826]),
			.SE(gen[2827]),

			.SELF(gen[2766]),
			.cell_state(gen[2766])
		); 

/******************* CELL 2767 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2767 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2706]),
			.N(gen[2707]),
			.NE(gen[2708]),

			.O(gen[2766]),
			.E(gen[2768]),

			.SO(gen[2826]),
			.S(gen[2827]),
			.SE(gen[2828]),

			.SELF(gen[2767]),
			.cell_state(gen[2767])
		); 

/******************* CELL 2768 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2768 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2707]),
			.N(gen[2708]),
			.NE(gen[2709]),

			.O(gen[2767]),
			.E(gen[2769]),

			.SO(gen[2827]),
			.S(gen[2828]),
			.SE(gen[2829]),

			.SELF(gen[2768]),
			.cell_state(gen[2768])
		); 

/******************* CELL 2769 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2769 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2708]),
			.N(gen[2709]),
			.NE(gen[2710]),

			.O(gen[2768]),
			.E(gen[2770]),

			.SO(gen[2828]),
			.S(gen[2829]),
			.SE(gen[2830]),

			.SELF(gen[2769]),
			.cell_state(gen[2769])
		); 

/******************* CELL 2770 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2770 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2709]),
			.N(gen[2710]),
			.NE(gen[2711]),

			.O(gen[2769]),
			.E(gen[2771]),

			.SO(gen[2829]),
			.S(gen[2830]),
			.SE(gen[2831]),

			.SELF(gen[2770]),
			.cell_state(gen[2770])
		); 

/******************* CELL 2771 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2771 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2710]),
			.N(gen[2711]),
			.NE(gen[2712]),

			.O(gen[2770]),
			.E(gen[2772]),

			.SO(gen[2830]),
			.S(gen[2831]),
			.SE(gen[2832]),

			.SELF(gen[2771]),
			.cell_state(gen[2771])
		); 

/******************* CELL 2772 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2772 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2711]),
			.N(gen[2712]),
			.NE(gen[2713]),

			.O(gen[2771]),
			.E(gen[2773]),

			.SO(gen[2831]),
			.S(gen[2832]),
			.SE(gen[2833]),

			.SELF(gen[2772]),
			.cell_state(gen[2772])
		); 

/******************* CELL 2773 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2773 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2712]),
			.N(gen[2713]),
			.NE(gen[2714]),

			.O(gen[2772]),
			.E(gen[2774]),

			.SO(gen[2832]),
			.S(gen[2833]),
			.SE(gen[2834]),

			.SELF(gen[2773]),
			.cell_state(gen[2773])
		); 

/******************* CELL 2774 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2774 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2713]),
			.N(gen[2714]),
			.NE(gen[2715]),

			.O(gen[2773]),
			.E(gen[2775]),

			.SO(gen[2833]),
			.S(gen[2834]),
			.SE(gen[2835]),

			.SELF(gen[2774]),
			.cell_state(gen[2774])
		); 

/******************* CELL 2775 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2775 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2714]),
			.N(gen[2715]),
			.NE(gen[2716]),

			.O(gen[2774]),
			.E(gen[2776]),

			.SO(gen[2834]),
			.S(gen[2835]),
			.SE(gen[2836]),

			.SELF(gen[2775]),
			.cell_state(gen[2775])
		); 

/******************* CELL 2776 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2776 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2715]),
			.N(gen[2716]),
			.NE(gen[2717]),

			.O(gen[2775]),
			.E(gen[2777]),

			.SO(gen[2835]),
			.S(gen[2836]),
			.SE(gen[2837]),

			.SELF(gen[2776]),
			.cell_state(gen[2776])
		); 

/******************* CELL 2777 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2777 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2716]),
			.N(gen[2717]),
			.NE(gen[2718]),

			.O(gen[2776]),
			.E(gen[2778]),

			.SO(gen[2836]),
			.S(gen[2837]),
			.SE(gen[2838]),

			.SELF(gen[2777]),
			.cell_state(gen[2777])
		); 

/******************* CELL 2778 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2778 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2717]),
			.N(gen[2718]),
			.NE(gen[2719]),

			.O(gen[2777]),
			.E(gen[2779]),

			.SO(gen[2837]),
			.S(gen[2838]),
			.SE(gen[2839]),

			.SELF(gen[2778]),
			.cell_state(gen[2778])
		); 

/******************* CELL 2779 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2779 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2718]),
			.N(gen[2719]),
			.NE(gen[2720]),

			.O(gen[2778]),
			.E(gen[2780]),

			.SO(gen[2838]),
			.S(gen[2839]),
			.SE(gen[2840]),

			.SELF(gen[2779]),
			.cell_state(gen[2779])
		); 

/******************* CELL 2780 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2780 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2719]),
			.N(gen[2720]),
			.NE(gen[2721]),

			.O(gen[2779]),
			.E(gen[2781]),

			.SO(gen[2839]),
			.S(gen[2840]),
			.SE(gen[2841]),

			.SELF(gen[2780]),
			.cell_state(gen[2780])
		); 

/******************* CELL 2781 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2781 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2720]),
			.N(gen[2721]),
			.NE(gen[2722]),

			.O(gen[2780]),
			.E(gen[2782]),

			.SO(gen[2840]),
			.S(gen[2841]),
			.SE(gen[2842]),

			.SELF(gen[2781]),
			.cell_state(gen[2781])
		); 

/******************* CELL 2782 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2782 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2721]),
			.N(gen[2722]),
			.NE(gen[2723]),

			.O(gen[2781]),
			.E(gen[2783]),

			.SO(gen[2841]),
			.S(gen[2842]),
			.SE(gen[2843]),

			.SELF(gen[2782]),
			.cell_state(gen[2782])
		); 

/******************* CELL 2783 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2783 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2722]),
			.N(gen[2723]),
			.NE(gen[2724]),

			.O(gen[2782]),
			.E(gen[2784]),

			.SO(gen[2842]),
			.S(gen[2843]),
			.SE(gen[2844]),

			.SELF(gen[2783]),
			.cell_state(gen[2783])
		); 

/******************* CELL 2784 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2784 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2723]),
			.N(gen[2724]),
			.NE(gen[2725]),

			.O(gen[2783]),
			.E(gen[2785]),

			.SO(gen[2843]),
			.S(gen[2844]),
			.SE(gen[2845]),

			.SELF(gen[2784]),
			.cell_state(gen[2784])
		); 

/******************* CELL 2785 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2785 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2724]),
			.N(gen[2725]),
			.NE(gen[2726]),

			.O(gen[2784]),
			.E(gen[2786]),

			.SO(gen[2844]),
			.S(gen[2845]),
			.SE(gen[2846]),

			.SELF(gen[2785]),
			.cell_state(gen[2785])
		); 

/******************* CELL 2786 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2786 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2725]),
			.N(gen[2726]),
			.NE(gen[2727]),

			.O(gen[2785]),
			.E(gen[2787]),

			.SO(gen[2845]),
			.S(gen[2846]),
			.SE(gen[2847]),

			.SELF(gen[2786]),
			.cell_state(gen[2786])
		); 

/******************* CELL 2787 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2787 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2726]),
			.N(gen[2727]),
			.NE(gen[2728]),

			.O(gen[2786]),
			.E(gen[2788]),

			.SO(gen[2846]),
			.S(gen[2847]),
			.SE(gen[2848]),

			.SELF(gen[2787]),
			.cell_state(gen[2787])
		); 

/******************* CELL 2788 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2788 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2727]),
			.N(gen[2728]),
			.NE(gen[2729]),

			.O(gen[2787]),
			.E(gen[2789]),

			.SO(gen[2847]),
			.S(gen[2848]),
			.SE(gen[2849]),

			.SELF(gen[2788]),
			.cell_state(gen[2788])
		); 

/******************* CELL 2789 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2789 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2728]),
			.N(gen[2729]),
			.NE(gen[2730]),

			.O(gen[2788]),
			.E(gen[2790]),

			.SO(gen[2848]),
			.S(gen[2849]),
			.SE(gen[2850]),

			.SELF(gen[2789]),
			.cell_state(gen[2789])
		); 

/******************* CELL 2790 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2790 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2729]),
			.N(gen[2730]),
			.NE(gen[2731]),

			.O(gen[2789]),
			.E(gen[2791]),

			.SO(gen[2849]),
			.S(gen[2850]),
			.SE(gen[2851]),

			.SELF(gen[2790]),
			.cell_state(gen[2790])
		); 

/******************* CELL 2791 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2791 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2730]),
			.N(gen[2731]),
			.NE(gen[2732]),

			.O(gen[2790]),
			.E(gen[2792]),

			.SO(gen[2850]),
			.S(gen[2851]),
			.SE(gen[2852]),

			.SELF(gen[2791]),
			.cell_state(gen[2791])
		); 

/******************* CELL 2792 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2792 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2731]),
			.N(gen[2732]),
			.NE(gen[2733]),

			.O(gen[2791]),
			.E(gen[2793]),

			.SO(gen[2851]),
			.S(gen[2852]),
			.SE(gen[2853]),

			.SELF(gen[2792]),
			.cell_state(gen[2792])
		); 

/******************* CELL 2793 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2793 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2732]),
			.N(gen[2733]),
			.NE(gen[2734]),

			.O(gen[2792]),
			.E(gen[2794]),

			.SO(gen[2852]),
			.S(gen[2853]),
			.SE(gen[2854]),

			.SELF(gen[2793]),
			.cell_state(gen[2793])
		); 

/******************* CELL 2794 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2794 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2733]),
			.N(gen[2734]),
			.NE(gen[2735]),

			.O(gen[2793]),
			.E(gen[2795]),

			.SO(gen[2853]),
			.S(gen[2854]),
			.SE(gen[2855]),

			.SELF(gen[2794]),
			.cell_state(gen[2794])
		); 

/******************* CELL 2795 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2795 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2734]),
			.N(gen[2735]),
			.NE(gen[2736]),

			.O(gen[2794]),
			.E(gen[2796]),

			.SO(gen[2854]),
			.S(gen[2855]),
			.SE(gen[2856]),

			.SELF(gen[2795]),
			.cell_state(gen[2795])
		); 

/******************* CELL 2796 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2796 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2735]),
			.N(gen[2736]),
			.NE(gen[2737]),

			.O(gen[2795]),
			.E(gen[2797]),

			.SO(gen[2855]),
			.S(gen[2856]),
			.SE(gen[2857]),

			.SELF(gen[2796]),
			.cell_state(gen[2796])
		); 

/******************* CELL 2797 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2797 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2736]),
			.N(gen[2737]),
			.NE(gen[2738]),

			.O(gen[2796]),
			.E(gen[2798]),

			.SO(gen[2856]),
			.S(gen[2857]),
			.SE(gen[2858]),

			.SELF(gen[2797]),
			.cell_state(gen[2797])
		); 

/******************* CELL 2798 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2798 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2737]),
			.N(gen[2738]),
			.NE(gen[2739]),

			.O(gen[2797]),
			.E(gen[2799]),

			.SO(gen[2857]),
			.S(gen[2858]),
			.SE(gen[2859]),

			.SELF(gen[2798]),
			.cell_state(gen[2798])
		); 

/******************* CELL 2799 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2799 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2738]),
			.N(gen[2739]),
			.NE(gen[2740]),

			.O(gen[2798]),
			.E(gen[2800]),

			.SO(gen[2858]),
			.S(gen[2859]),
			.SE(gen[2860]),

			.SELF(gen[2799]),
			.cell_state(gen[2799])
		); 

/******************* CELL 2800 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2800 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2739]),
			.N(gen[2740]),
			.NE(gen[2741]),

			.O(gen[2799]),
			.E(gen[2801]),

			.SO(gen[2859]),
			.S(gen[2860]),
			.SE(gen[2861]),

			.SELF(gen[2800]),
			.cell_state(gen[2800])
		); 

/******************* CELL 2801 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2801 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2740]),
			.N(gen[2741]),
			.NE(gen[2742]),

			.O(gen[2800]),
			.E(gen[2802]),

			.SO(gen[2860]),
			.S(gen[2861]),
			.SE(gen[2862]),

			.SELF(gen[2801]),
			.cell_state(gen[2801])
		); 

/******************* CELL 2802 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2802 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2741]),
			.N(gen[2742]),
			.NE(gen[2743]),

			.O(gen[2801]),
			.E(gen[2803]),

			.SO(gen[2861]),
			.S(gen[2862]),
			.SE(gen[2863]),

			.SELF(gen[2802]),
			.cell_state(gen[2802])
		); 

/******************* CELL 2803 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2803 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2742]),
			.N(gen[2743]),
			.NE(gen[2744]),

			.O(gen[2802]),
			.E(gen[2804]),

			.SO(gen[2862]),
			.S(gen[2863]),
			.SE(gen[2864]),

			.SELF(gen[2803]),
			.cell_state(gen[2803])
		); 

/******************* CELL 2804 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2804 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2743]),
			.N(gen[2744]),
			.NE(gen[2745]),

			.O(gen[2803]),
			.E(gen[2805]),

			.SO(gen[2863]),
			.S(gen[2864]),
			.SE(gen[2865]),

			.SELF(gen[2804]),
			.cell_state(gen[2804])
		); 

/******************* CELL 2805 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2805 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2744]),
			.N(gen[2745]),
			.NE(gen[2746]),

			.O(gen[2804]),
			.E(gen[2806]),

			.SO(gen[2864]),
			.S(gen[2865]),
			.SE(gen[2866]),

			.SELF(gen[2805]),
			.cell_state(gen[2805])
		); 

/******************* CELL 2806 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2806 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2745]),
			.N(gen[2746]),
			.NE(gen[2747]),

			.O(gen[2805]),
			.E(gen[2807]),

			.SO(gen[2865]),
			.S(gen[2866]),
			.SE(gen[2867]),

			.SELF(gen[2806]),
			.cell_state(gen[2806])
		); 

/******************* CELL 2807 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2807 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2746]),
			.N(gen[2747]),
			.NE(gen[2748]),

			.O(gen[2806]),
			.E(gen[2808]),

			.SO(gen[2866]),
			.S(gen[2867]),
			.SE(gen[2868]),

			.SELF(gen[2807]),
			.cell_state(gen[2807])
		); 

/******************* CELL 2808 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2808 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2747]),
			.N(gen[2748]),
			.NE(gen[2749]),

			.O(gen[2807]),
			.E(gen[2809]),

			.SO(gen[2867]),
			.S(gen[2868]),
			.SE(gen[2869]),

			.SELF(gen[2808]),
			.cell_state(gen[2808])
		); 

/******************* CELL 2809 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2809 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2748]),
			.N(gen[2749]),
			.NE(gen[2750]),

			.O(gen[2808]),
			.E(gen[2810]),

			.SO(gen[2868]),
			.S(gen[2869]),
			.SE(gen[2870]),

			.SELF(gen[2809]),
			.cell_state(gen[2809])
		); 

/******************* CELL 2810 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2810 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2749]),
			.N(gen[2750]),
			.NE(gen[2751]),

			.O(gen[2809]),
			.E(gen[2811]),

			.SO(gen[2869]),
			.S(gen[2870]),
			.SE(gen[2871]),

			.SELF(gen[2810]),
			.cell_state(gen[2810])
		); 

/******************* CELL 2811 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2811 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2750]),
			.N(gen[2751]),
			.NE(gen[2752]),

			.O(gen[2810]),
			.E(gen[2812]),

			.SO(gen[2870]),
			.S(gen[2871]),
			.SE(gen[2872]),

			.SELF(gen[2811]),
			.cell_state(gen[2811])
		); 

/******************* CELL 2812 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2812 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2751]),
			.N(gen[2752]),
			.NE(gen[2753]),

			.O(gen[2811]),
			.E(gen[2813]),

			.SO(gen[2871]),
			.S(gen[2872]),
			.SE(gen[2873]),

			.SELF(gen[2812]),
			.cell_state(gen[2812])
		); 

/******************* CELL 2813 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2813 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2752]),
			.N(gen[2753]),
			.NE(gen[2754]),

			.O(gen[2812]),
			.E(gen[2814]),

			.SO(gen[2872]),
			.S(gen[2873]),
			.SE(gen[2874]),

			.SELF(gen[2813]),
			.cell_state(gen[2813])
		); 

/******************* CELL 2814 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2814 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2753]),
			.N(gen[2754]),
			.NE(gen[2755]),

			.O(gen[2813]),
			.E(gen[2815]),

			.SO(gen[2873]),
			.S(gen[2874]),
			.SE(gen[2875]),

			.SELF(gen[2814]),
			.cell_state(gen[2814])
		); 

/******************* CELL 2815 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2815 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2754]),
			.N(gen[2755]),
			.NE(gen[2756]),

			.O(gen[2814]),
			.E(gen[2816]),

			.SO(gen[2874]),
			.S(gen[2875]),
			.SE(gen[2876]),

			.SELF(gen[2815]),
			.cell_state(gen[2815])
		); 

/******************* CELL 2816 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2816 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2755]),
			.N(gen[2756]),
			.NE(gen[2757]),

			.O(gen[2815]),
			.E(gen[2817]),

			.SO(gen[2875]),
			.S(gen[2876]),
			.SE(gen[2877]),

			.SELF(gen[2816]),
			.cell_state(gen[2816])
		); 

/******************* CELL 2817 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2817 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2756]),
			.N(gen[2757]),
			.NE(gen[2758]),

			.O(gen[2816]),
			.E(gen[2818]),

			.SO(gen[2876]),
			.S(gen[2877]),
			.SE(gen[2878]),

			.SELF(gen[2817]),
			.cell_state(gen[2817])
		); 

/******************* CELL 2818 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2818 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2757]),
			.N(gen[2758]),
			.NE(gen[2759]),

			.O(gen[2817]),
			.E(gen[2819]),

			.SO(gen[2877]),
			.S(gen[2878]),
			.SE(gen[2879]),

			.SELF(gen[2818]),
			.cell_state(gen[2818])
		); 

/******************* CELL 2819 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2819 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2758]),
			.N(gen[2759]),
			.NE(gen[2758]),

			.O(gen[2818]),
			.E(gen[2818]),

			.SO(gen[2878]),
			.S(gen[2879]),
			.SE(gen[2878]),

			.SELF(gen[2819]),
			.cell_state(gen[2819])
		); 

/******************* CELL 2820 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2820 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2761]),
			.N(gen[2760]),
			.NE(gen[2761]),

			.O(gen[2821]),
			.E(gen[2821]),

			.SO(gen[2881]),
			.S(gen[2880]),
			.SE(gen[2881]),

			.SELF(gen[2820]),
			.cell_state(gen[2820])
		); 

/******************* CELL 2821 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2821 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2760]),
			.N(gen[2761]),
			.NE(gen[2762]),

			.O(gen[2820]),
			.E(gen[2822]),

			.SO(gen[2880]),
			.S(gen[2881]),
			.SE(gen[2882]),

			.SELF(gen[2821]),
			.cell_state(gen[2821])
		); 

/******************* CELL 2822 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2822 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2761]),
			.N(gen[2762]),
			.NE(gen[2763]),

			.O(gen[2821]),
			.E(gen[2823]),

			.SO(gen[2881]),
			.S(gen[2882]),
			.SE(gen[2883]),

			.SELF(gen[2822]),
			.cell_state(gen[2822])
		); 

/******************* CELL 2823 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2823 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2762]),
			.N(gen[2763]),
			.NE(gen[2764]),

			.O(gen[2822]),
			.E(gen[2824]),

			.SO(gen[2882]),
			.S(gen[2883]),
			.SE(gen[2884]),

			.SELF(gen[2823]),
			.cell_state(gen[2823])
		); 

/******************* CELL 2824 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2824 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2763]),
			.N(gen[2764]),
			.NE(gen[2765]),

			.O(gen[2823]),
			.E(gen[2825]),

			.SO(gen[2883]),
			.S(gen[2884]),
			.SE(gen[2885]),

			.SELF(gen[2824]),
			.cell_state(gen[2824])
		); 

/******************* CELL 2825 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2825 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2764]),
			.N(gen[2765]),
			.NE(gen[2766]),

			.O(gen[2824]),
			.E(gen[2826]),

			.SO(gen[2884]),
			.S(gen[2885]),
			.SE(gen[2886]),

			.SELF(gen[2825]),
			.cell_state(gen[2825])
		); 

/******************* CELL 2826 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2826 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2765]),
			.N(gen[2766]),
			.NE(gen[2767]),

			.O(gen[2825]),
			.E(gen[2827]),

			.SO(gen[2885]),
			.S(gen[2886]),
			.SE(gen[2887]),

			.SELF(gen[2826]),
			.cell_state(gen[2826])
		); 

/******************* CELL 2827 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2827 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2766]),
			.N(gen[2767]),
			.NE(gen[2768]),

			.O(gen[2826]),
			.E(gen[2828]),

			.SO(gen[2886]),
			.S(gen[2887]),
			.SE(gen[2888]),

			.SELF(gen[2827]),
			.cell_state(gen[2827])
		); 

/******************* CELL 2828 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2828 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2767]),
			.N(gen[2768]),
			.NE(gen[2769]),

			.O(gen[2827]),
			.E(gen[2829]),

			.SO(gen[2887]),
			.S(gen[2888]),
			.SE(gen[2889]),

			.SELF(gen[2828]),
			.cell_state(gen[2828])
		); 

/******************* CELL 2829 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2829 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2768]),
			.N(gen[2769]),
			.NE(gen[2770]),

			.O(gen[2828]),
			.E(gen[2830]),

			.SO(gen[2888]),
			.S(gen[2889]),
			.SE(gen[2890]),

			.SELF(gen[2829]),
			.cell_state(gen[2829])
		); 

/******************* CELL 2830 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2830 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2769]),
			.N(gen[2770]),
			.NE(gen[2771]),

			.O(gen[2829]),
			.E(gen[2831]),

			.SO(gen[2889]),
			.S(gen[2890]),
			.SE(gen[2891]),

			.SELF(gen[2830]),
			.cell_state(gen[2830])
		); 

/******************* CELL 2831 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2831 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2770]),
			.N(gen[2771]),
			.NE(gen[2772]),

			.O(gen[2830]),
			.E(gen[2832]),

			.SO(gen[2890]),
			.S(gen[2891]),
			.SE(gen[2892]),

			.SELF(gen[2831]),
			.cell_state(gen[2831])
		); 

/******************* CELL 2832 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2832 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2771]),
			.N(gen[2772]),
			.NE(gen[2773]),

			.O(gen[2831]),
			.E(gen[2833]),

			.SO(gen[2891]),
			.S(gen[2892]),
			.SE(gen[2893]),

			.SELF(gen[2832]),
			.cell_state(gen[2832])
		); 

/******************* CELL 2833 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2833 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2772]),
			.N(gen[2773]),
			.NE(gen[2774]),

			.O(gen[2832]),
			.E(gen[2834]),

			.SO(gen[2892]),
			.S(gen[2893]),
			.SE(gen[2894]),

			.SELF(gen[2833]),
			.cell_state(gen[2833])
		); 

/******************* CELL 2834 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2834 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2773]),
			.N(gen[2774]),
			.NE(gen[2775]),

			.O(gen[2833]),
			.E(gen[2835]),

			.SO(gen[2893]),
			.S(gen[2894]),
			.SE(gen[2895]),

			.SELF(gen[2834]),
			.cell_state(gen[2834])
		); 

/******************* CELL 2835 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2835 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2774]),
			.N(gen[2775]),
			.NE(gen[2776]),

			.O(gen[2834]),
			.E(gen[2836]),

			.SO(gen[2894]),
			.S(gen[2895]),
			.SE(gen[2896]),

			.SELF(gen[2835]),
			.cell_state(gen[2835])
		); 

/******************* CELL 2836 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2836 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2775]),
			.N(gen[2776]),
			.NE(gen[2777]),

			.O(gen[2835]),
			.E(gen[2837]),

			.SO(gen[2895]),
			.S(gen[2896]),
			.SE(gen[2897]),

			.SELF(gen[2836]),
			.cell_state(gen[2836])
		); 

/******************* CELL 2837 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2837 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2776]),
			.N(gen[2777]),
			.NE(gen[2778]),

			.O(gen[2836]),
			.E(gen[2838]),

			.SO(gen[2896]),
			.S(gen[2897]),
			.SE(gen[2898]),

			.SELF(gen[2837]),
			.cell_state(gen[2837])
		); 

/******************* CELL 2838 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2838 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2777]),
			.N(gen[2778]),
			.NE(gen[2779]),

			.O(gen[2837]),
			.E(gen[2839]),

			.SO(gen[2897]),
			.S(gen[2898]),
			.SE(gen[2899]),

			.SELF(gen[2838]),
			.cell_state(gen[2838])
		); 

/******************* CELL 2839 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2839 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2778]),
			.N(gen[2779]),
			.NE(gen[2780]),

			.O(gen[2838]),
			.E(gen[2840]),

			.SO(gen[2898]),
			.S(gen[2899]),
			.SE(gen[2900]),

			.SELF(gen[2839]),
			.cell_state(gen[2839])
		); 

/******************* CELL 2840 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2840 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2779]),
			.N(gen[2780]),
			.NE(gen[2781]),

			.O(gen[2839]),
			.E(gen[2841]),

			.SO(gen[2899]),
			.S(gen[2900]),
			.SE(gen[2901]),

			.SELF(gen[2840]),
			.cell_state(gen[2840])
		); 

/******************* CELL 2841 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2841 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2780]),
			.N(gen[2781]),
			.NE(gen[2782]),

			.O(gen[2840]),
			.E(gen[2842]),

			.SO(gen[2900]),
			.S(gen[2901]),
			.SE(gen[2902]),

			.SELF(gen[2841]),
			.cell_state(gen[2841])
		); 

/******************* CELL 2842 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2842 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2781]),
			.N(gen[2782]),
			.NE(gen[2783]),

			.O(gen[2841]),
			.E(gen[2843]),

			.SO(gen[2901]),
			.S(gen[2902]),
			.SE(gen[2903]),

			.SELF(gen[2842]),
			.cell_state(gen[2842])
		); 

/******************* CELL 2843 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2843 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2782]),
			.N(gen[2783]),
			.NE(gen[2784]),

			.O(gen[2842]),
			.E(gen[2844]),

			.SO(gen[2902]),
			.S(gen[2903]),
			.SE(gen[2904]),

			.SELF(gen[2843]),
			.cell_state(gen[2843])
		); 

/******************* CELL 2844 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2844 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2783]),
			.N(gen[2784]),
			.NE(gen[2785]),

			.O(gen[2843]),
			.E(gen[2845]),

			.SO(gen[2903]),
			.S(gen[2904]),
			.SE(gen[2905]),

			.SELF(gen[2844]),
			.cell_state(gen[2844])
		); 

/******************* CELL 2845 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2845 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2784]),
			.N(gen[2785]),
			.NE(gen[2786]),

			.O(gen[2844]),
			.E(gen[2846]),

			.SO(gen[2904]),
			.S(gen[2905]),
			.SE(gen[2906]),

			.SELF(gen[2845]),
			.cell_state(gen[2845])
		); 

/******************* CELL 2846 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2846 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2785]),
			.N(gen[2786]),
			.NE(gen[2787]),

			.O(gen[2845]),
			.E(gen[2847]),

			.SO(gen[2905]),
			.S(gen[2906]),
			.SE(gen[2907]),

			.SELF(gen[2846]),
			.cell_state(gen[2846])
		); 

/******************* CELL 2847 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2847 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2786]),
			.N(gen[2787]),
			.NE(gen[2788]),

			.O(gen[2846]),
			.E(gen[2848]),

			.SO(gen[2906]),
			.S(gen[2907]),
			.SE(gen[2908]),

			.SELF(gen[2847]),
			.cell_state(gen[2847])
		); 

/******************* CELL 2848 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2848 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2787]),
			.N(gen[2788]),
			.NE(gen[2789]),

			.O(gen[2847]),
			.E(gen[2849]),

			.SO(gen[2907]),
			.S(gen[2908]),
			.SE(gen[2909]),

			.SELF(gen[2848]),
			.cell_state(gen[2848])
		); 

/******************* CELL 2849 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2849 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2788]),
			.N(gen[2789]),
			.NE(gen[2790]),

			.O(gen[2848]),
			.E(gen[2850]),

			.SO(gen[2908]),
			.S(gen[2909]),
			.SE(gen[2910]),

			.SELF(gen[2849]),
			.cell_state(gen[2849])
		); 

/******************* CELL 2850 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2850 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2789]),
			.N(gen[2790]),
			.NE(gen[2791]),

			.O(gen[2849]),
			.E(gen[2851]),

			.SO(gen[2909]),
			.S(gen[2910]),
			.SE(gen[2911]),

			.SELF(gen[2850]),
			.cell_state(gen[2850])
		); 

/******************* CELL 2851 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2851 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2790]),
			.N(gen[2791]),
			.NE(gen[2792]),

			.O(gen[2850]),
			.E(gen[2852]),

			.SO(gen[2910]),
			.S(gen[2911]),
			.SE(gen[2912]),

			.SELF(gen[2851]),
			.cell_state(gen[2851])
		); 

/******************* CELL 2852 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2852 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2791]),
			.N(gen[2792]),
			.NE(gen[2793]),

			.O(gen[2851]),
			.E(gen[2853]),

			.SO(gen[2911]),
			.S(gen[2912]),
			.SE(gen[2913]),

			.SELF(gen[2852]),
			.cell_state(gen[2852])
		); 

/******************* CELL 2853 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2853 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2792]),
			.N(gen[2793]),
			.NE(gen[2794]),

			.O(gen[2852]),
			.E(gen[2854]),

			.SO(gen[2912]),
			.S(gen[2913]),
			.SE(gen[2914]),

			.SELF(gen[2853]),
			.cell_state(gen[2853])
		); 

/******************* CELL 2854 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2854 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2793]),
			.N(gen[2794]),
			.NE(gen[2795]),

			.O(gen[2853]),
			.E(gen[2855]),

			.SO(gen[2913]),
			.S(gen[2914]),
			.SE(gen[2915]),

			.SELF(gen[2854]),
			.cell_state(gen[2854])
		); 

/******************* CELL 2855 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2855 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2794]),
			.N(gen[2795]),
			.NE(gen[2796]),

			.O(gen[2854]),
			.E(gen[2856]),

			.SO(gen[2914]),
			.S(gen[2915]),
			.SE(gen[2916]),

			.SELF(gen[2855]),
			.cell_state(gen[2855])
		); 

/******************* CELL 2856 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2856 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2795]),
			.N(gen[2796]),
			.NE(gen[2797]),

			.O(gen[2855]),
			.E(gen[2857]),

			.SO(gen[2915]),
			.S(gen[2916]),
			.SE(gen[2917]),

			.SELF(gen[2856]),
			.cell_state(gen[2856])
		); 

/******************* CELL 2857 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2857 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2796]),
			.N(gen[2797]),
			.NE(gen[2798]),

			.O(gen[2856]),
			.E(gen[2858]),

			.SO(gen[2916]),
			.S(gen[2917]),
			.SE(gen[2918]),

			.SELF(gen[2857]),
			.cell_state(gen[2857])
		); 

/******************* CELL 2858 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2858 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2797]),
			.N(gen[2798]),
			.NE(gen[2799]),

			.O(gen[2857]),
			.E(gen[2859]),

			.SO(gen[2917]),
			.S(gen[2918]),
			.SE(gen[2919]),

			.SELF(gen[2858]),
			.cell_state(gen[2858])
		); 

/******************* CELL 2859 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2859 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2798]),
			.N(gen[2799]),
			.NE(gen[2800]),

			.O(gen[2858]),
			.E(gen[2860]),

			.SO(gen[2918]),
			.S(gen[2919]),
			.SE(gen[2920]),

			.SELF(gen[2859]),
			.cell_state(gen[2859])
		); 

/******************* CELL 2860 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2860 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2799]),
			.N(gen[2800]),
			.NE(gen[2801]),

			.O(gen[2859]),
			.E(gen[2861]),

			.SO(gen[2919]),
			.S(gen[2920]),
			.SE(gen[2921]),

			.SELF(gen[2860]),
			.cell_state(gen[2860])
		); 

/******************* CELL 2861 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2861 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2800]),
			.N(gen[2801]),
			.NE(gen[2802]),

			.O(gen[2860]),
			.E(gen[2862]),

			.SO(gen[2920]),
			.S(gen[2921]),
			.SE(gen[2922]),

			.SELF(gen[2861]),
			.cell_state(gen[2861])
		); 

/******************* CELL 2862 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2862 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2801]),
			.N(gen[2802]),
			.NE(gen[2803]),

			.O(gen[2861]),
			.E(gen[2863]),

			.SO(gen[2921]),
			.S(gen[2922]),
			.SE(gen[2923]),

			.SELF(gen[2862]),
			.cell_state(gen[2862])
		); 

/******************* CELL 2863 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2863 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2802]),
			.N(gen[2803]),
			.NE(gen[2804]),

			.O(gen[2862]),
			.E(gen[2864]),

			.SO(gen[2922]),
			.S(gen[2923]),
			.SE(gen[2924]),

			.SELF(gen[2863]),
			.cell_state(gen[2863])
		); 

/******************* CELL 2864 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2864 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2803]),
			.N(gen[2804]),
			.NE(gen[2805]),

			.O(gen[2863]),
			.E(gen[2865]),

			.SO(gen[2923]),
			.S(gen[2924]),
			.SE(gen[2925]),

			.SELF(gen[2864]),
			.cell_state(gen[2864])
		); 

/******************* CELL 2865 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2865 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2804]),
			.N(gen[2805]),
			.NE(gen[2806]),

			.O(gen[2864]),
			.E(gen[2866]),

			.SO(gen[2924]),
			.S(gen[2925]),
			.SE(gen[2926]),

			.SELF(gen[2865]),
			.cell_state(gen[2865])
		); 

/******************* CELL 2866 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2866 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2805]),
			.N(gen[2806]),
			.NE(gen[2807]),

			.O(gen[2865]),
			.E(gen[2867]),

			.SO(gen[2925]),
			.S(gen[2926]),
			.SE(gen[2927]),

			.SELF(gen[2866]),
			.cell_state(gen[2866])
		); 

/******************* CELL 2867 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2867 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2806]),
			.N(gen[2807]),
			.NE(gen[2808]),

			.O(gen[2866]),
			.E(gen[2868]),

			.SO(gen[2926]),
			.S(gen[2927]),
			.SE(gen[2928]),

			.SELF(gen[2867]),
			.cell_state(gen[2867])
		); 

/******************* CELL 2868 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2868 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2807]),
			.N(gen[2808]),
			.NE(gen[2809]),

			.O(gen[2867]),
			.E(gen[2869]),

			.SO(gen[2927]),
			.S(gen[2928]),
			.SE(gen[2929]),

			.SELF(gen[2868]),
			.cell_state(gen[2868])
		); 

/******************* CELL 2869 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2869 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2808]),
			.N(gen[2809]),
			.NE(gen[2810]),

			.O(gen[2868]),
			.E(gen[2870]),

			.SO(gen[2928]),
			.S(gen[2929]),
			.SE(gen[2930]),

			.SELF(gen[2869]),
			.cell_state(gen[2869])
		); 

/******************* CELL 2870 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2870 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2809]),
			.N(gen[2810]),
			.NE(gen[2811]),

			.O(gen[2869]),
			.E(gen[2871]),

			.SO(gen[2929]),
			.S(gen[2930]),
			.SE(gen[2931]),

			.SELF(gen[2870]),
			.cell_state(gen[2870])
		); 

/******************* CELL 2871 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2871 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2810]),
			.N(gen[2811]),
			.NE(gen[2812]),

			.O(gen[2870]),
			.E(gen[2872]),

			.SO(gen[2930]),
			.S(gen[2931]),
			.SE(gen[2932]),

			.SELF(gen[2871]),
			.cell_state(gen[2871])
		); 

/******************* CELL 2872 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2872 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2811]),
			.N(gen[2812]),
			.NE(gen[2813]),

			.O(gen[2871]),
			.E(gen[2873]),

			.SO(gen[2931]),
			.S(gen[2932]),
			.SE(gen[2933]),

			.SELF(gen[2872]),
			.cell_state(gen[2872])
		); 

/******************* CELL 2873 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2873 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2812]),
			.N(gen[2813]),
			.NE(gen[2814]),

			.O(gen[2872]),
			.E(gen[2874]),

			.SO(gen[2932]),
			.S(gen[2933]),
			.SE(gen[2934]),

			.SELF(gen[2873]),
			.cell_state(gen[2873])
		); 

/******************* CELL 2874 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2874 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2813]),
			.N(gen[2814]),
			.NE(gen[2815]),

			.O(gen[2873]),
			.E(gen[2875]),

			.SO(gen[2933]),
			.S(gen[2934]),
			.SE(gen[2935]),

			.SELF(gen[2874]),
			.cell_state(gen[2874])
		); 

/******************* CELL 2875 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2875 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2814]),
			.N(gen[2815]),
			.NE(gen[2816]),

			.O(gen[2874]),
			.E(gen[2876]),

			.SO(gen[2934]),
			.S(gen[2935]),
			.SE(gen[2936]),

			.SELF(gen[2875]),
			.cell_state(gen[2875])
		); 

/******************* CELL 2876 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2876 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2815]),
			.N(gen[2816]),
			.NE(gen[2817]),

			.O(gen[2875]),
			.E(gen[2877]),

			.SO(gen[2935]),
			.S(gen[2936]),
			.SE(gen[2937]),

			.SELF(gen[2876]),
			.cell_state(gen[2876])
		); 

/******************* CELL 2877 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2877 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2816]),
			.N(gen[2817]),
			.NE(gen[2818]),

			.O(gen[2876]),
			.E(gen[2878]),

			.SO(gen[2936]),
			.S(gen[2937]),
			.SE(gen[2938]),

			.SELF(gen[2877]),
			.cell_state(gen[2877])
		); 

/******************* CELL 2878 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2878 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2817]),
			.N(gen[2818]),
			.NE(gen[2819]),

			.O(gen[2877]),
			.E(gen[2879]),

			.SO(gen[2937]),
			.S(gen[2938]),
			.SE(gen[2939]),

			.SELF(gen[2878]),
			.cell_state(gen[2878])
		); 

/******************* CELL 2879 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2879 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2818]),
			.N(gen[2819]),
			.NE(gen[2818]),

			.O(gen[2878]),
			.E(gen[2878]),

			.SO(gen[2938]),
			.S(gen[2939]),
			.SE(gen[2938]),

			.SELF(gen[2879]),
			.cell_state(gen[2879])
		); 

/******************* CELL 2880 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2880 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2821]),
			.N(gen[2820]),
			.NE(gen[2821]),

			.O(gen[2881]),
			.E(gen[2881]),

			.SO(gen[2941]),
			.S(gen[2940]),
			.SE(gen[2941]),

			.SELF(gen[2880]),
			.cell_state(gen[2880])
		); 

/******************* CELL 2881 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2881 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2820]),
			.N(gen[2821]),
			.NE(gen[2822]),

			.O(gen[2880]),
			.E(gen[2882]),

			.SO(gen[2940]),
			.S(gen[2941]),
			.SE(gen[2942]),

			.SELF(gen[2881]),
			.cell_state(gen[2881])
		); 

/******************* CELL 2882 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2882 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2821]),
			.N(gen[2822]),
			.NE(gen[2823]),

			.O(gen[2881]),
			.E(gen[2883]),

			.SO(gen[2941]),
			.S(gen[2942]),
			.SE(gen[2943]),

			.SELF(gen[2882]),
			.cell_state(gen[2882])
		); 

/******************* CELL 2883 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2883 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2822]),
			.N(gen[2823]),
			.NE(gen[2824]),

			.O(gen[2882]),
			.E(gen[2884]),

			.SO(gen[2942]),
			.S(gen[2943]),
			.SE(gen[2944]),

			.SELF(gen[2883]),
			.cell_state(gen[2883])
		); 

/******************* CELL 2884 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2884 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2823]),
			.N(gen[2824]),
			.NE(gen[2825]),

			.O(gen[2883]),
			.E(gen[2885]),

			.SO(gen[2943]),
			.S(gen[2944]),
			.SE(gen[2945]),

			.SELF(gen[2884]),
			.cell_state(gen[2884])
		); 

/******************* CELL 2885 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2885 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2824]),
			.N(gen[2825]),
			.NE(gen[2826]),

			.O(gen[2884]),
			.E(gen[2886]),

			.SO(gen[2944]),
			.S(gen[2945]),
			.SE(gen[2946]),

			.SELF(gen[2885]),
			.cell_state(gen[2885])
		); 

/******************* CELL 2886 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2886 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2825]),
			.N(gen[2826]),
			.NE(gen[2827]),

			.O(gen[2885]),
			.E(gen[2887]),

			.SO(gen[2945]),
			.S(gen[2946]),
			.SE(gen[2947]),

			.SELF(gen[2886]),
			.cell_state(gen[2886])
		); 

/******************* CELL 2887 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2887 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2826]),
			.N(gen[2827]),
			.NE(gen[2828]),

			.O(gen[2886]),
			.E(gen[2888]),

			.SO(gen[2946]),
			.S(gen[2947]),
			.SE(gen[2948]),

			.SELF(gen[2887]),
			.cell_state(gen[2887])
		); 

/******************* CELL 2888 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2888 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2827]),
			.N(gen[2828]),
			.NE(gen[2829]),

			.O(gen[2887]),
			.E(gen[2889]),

			.SO(gen[2947]),
			.S(gen[2948]),
			.SE(gen[2949]),

			.SELF(gen[2888]),
			.cell_state(gen[2888])
		); 

/******************* CELL 2889 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2889 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2828]),
			.N(gen[2829]),
			.NE(gen[2830]),

			.O(gen[2888]),
			.E(gen[2890]),

			.SO(gen[2948]),
			.S(gen[2949]),
			.SE(gen[2950]),

			.SELF(gen[2889]),
			.cell_state(gen[2889])
		); 

/******************* CELL 2890 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2890 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2829]),
			.N(gen[2830]),
			.NE(gen[2831]),

			.O(gen[2889]),
			.E(gen[2891]),

			.SO(gen[2949]),
			.S(gen[2950]),
			.SE(gen[2951]),

			.SELF(gen[2890]),
			.cell_state(gen[2890])
		); 

/******************* CELL 2891 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2891 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2830]),
			.N(gen[2831]),
			.NE(gen[2832]),

			.O(gen[2890]),
			.E(gen[2892]),

			.SO(gen[2950]),
			.S(gen[2951]),
			.SE(gen[2952]),

			.SELF(gen[2891]),
			.cell_state(gen[2891])
		); 

/******************* CELL 2892 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2892 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2831]),
			.N(gen[2832]),
			.NE(gen[2833]),

			.O(gen[2891]),
			.E(gen[2893]),

			.SO(gen[2951]),
			.S(gen[2952]),
			.SE(gen[2953]),

			.SELF(gen[2892]),
			.cell_state(gen[2892])
		); 

/******************* CELL 2893 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2893 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2832]),
			.N(gen[2833]),
			.NE(gen[2834]),

			.O(gen[2892]),
			.E(gen[2894]),

			.SO(gen[2952]),
			.S(gen[2953]),
			.SE(gen[2954]),

			.SELF(gen[2893]),
			.cell_state(gen[2893])
		); 

/******************* CELL 2894 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2894 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2833]),
			.N(gen[2834]),
			.NE(gen[2835]),

			.O(gen[2893]),
			.E(gen[2895]),

			.SO(gen[2953]),
			.S(gen[2954]),
			.SE(gen[2955]),

			.SELF(gen[2894]),
			.cell_state(gen[2894])
		); 

/******************* CELL 2895 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2895 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2834]),
			.N(gen[2835]),
			.NE(gen[2836]),

			.O(gen[2894]),
			.E(gen[2896]),

			.SO(gen[2954]),
			.S(gen[2955]),
			.SE(gen[2956]),

			.SELF(gen[2895]),
			.cell_state(gen[2895])
		); 

/******************* CELL 2896 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2896 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2835]),
			.N(gen[2836]),
			.NE(gen[2837]),

			.O(gen[2895]),
			.E(gen[2897]),

			.SO(gen[2955]),
			.S(gen[2956]),
			.SE(gen[2957]),

			.SELF(gen[2896]),
			.cell_state(gen[2896])
		); 

/******************* CELL 2897 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2897 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2836]),
			.N(gen[2837]),
			.NE(gen[2838]),

			.O(gen[2896]),
			.E(gen[2898]),

			.SO(gen[2956]),
			.S(gen[2957]),
			.SE(gen[2958]),

			.SELF(gen[2897]),
			.cell_state(gen[2897])
		); 

/******************* CELL 2898 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2898 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2837]),
			.N(gen[2838]),
			.NE(gen[2839]),

			.O(gen[2897]),
			.E(gen[2899]),

			.SO(gen[2957]),
			.S(gen[2958]),
			.SE(gen[2959]),

			.SELF(gen[2898]),
			.cell_state(gen[2898])
		); 

/******************* CELL 2899 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2899 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2838]),
			.N(gen[2839]),
			.NE(gen[2840]),

			.O(gen[2898]),
			.E(gen[2900]),

			.SO(gen[2958]),
			.S(gen[2959]),
			.SE(gen[2960]),

			.SELF(gen[2899]),
			.cell_state(gen[2899])
		); 

/******************* CELL 2900 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2900 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2839]),
			.N(gen[2840]),
			.NE(gen[2841]),

			.O(gen[2899]),
			.E(gen[2901]),

			.SO(gen[2959]),
			.S(gen[2960]),
			.SE(gen[2961]),

			.SELF(gen[2900]),
			.cell_state(gen[2900])
		); 

/******************* CELL 2901 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2901 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2840]),
			.N(gen[2841]),
			.NE(gen[2842]),

			.O(gen[2900]),
			.E(gen[2902]),

			.SO(gen[2960]),
			.S(gen[2961]),
			.SE(gen[2962]),

			.SELF(gen[2901]),
			.cell_state(gen[2901])
		); 

/******************* CELL 2902 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2902 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2841]),
			.N(gen[2842]),
			.NE(gen[2843]),

			.O(gen[2901]),
			.E(gen[2903]),

			.SO(gen[2961]),
			.S(gen[2962]),
			.SE(gen[2963]),

			.SELF(gen[2902]),
			.cell_state(gen[2902])
		); 

/******************* CELL 2903 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2903 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2842]),
			.N(gen[2843]),
			.NE(gen[2844]),

			.O(gen[2902]),
			.E(gen[2904]),

			.SO(gen[2962]),
			.S(gen[2963]),
			.SE(gen[2964]),

			.SELF(gen[2903]),
			.cell_state(gen[2903])
		); 

/******************* CELL 2904 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2904 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2843]),
			.N(gen[2844]),
			.NE(gen[2845]),

			.O(gen[2903]),
			.E(gen[2905]),

			.SO(gen[2963]),
			.S(gen[2964]),
			.SE(gen[2965]),

			.SELF(gen[2904]),
			.cell_state(gen[2904])
		); 

/******************* CELL 2905 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2905 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2844]),
			.N(gen[2845]),
			.NE(gen[2846]),

			.O(gen[2904]),
			.E(gen[2906]),

			.SO(gen[2964]),
			.S(gen[2965]),
			.SE(gen[2966]),

			.SELF(gen[2905]),
			.cell_state(gen[2905])
		); 

/******************* CELL 2906 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2906 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2845]),
			.N(gen[2846]),
			.NE(gen[2847]),

			.O(gen[2905]),
			.E(gen[2907]),

			.SO(gen[2965]),
			.S(gen[2966]),
			.SE(gen[2967]),

			.SELF(gen[2906]),
			.cell_state(gen[2906])
		); 

/******************* CELL 2907 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2907 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2846]),
			.N(gen[2847]),
			.NE(gen[2848]),

			.O(gen[2906]),
			.E(gen[2908]),

			.SO(gen[2966]),
			.S(gen[2967]),
			.SE(gen[2968]),

			.SELF(gen[2907]),
			.cell_state(gen[2907])
		); 

/******************* CELL 2908 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2908 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2847]),
			.N(gen[2848]),
			.NE(gen[2849]),

			.O(gen[2907]),
			.E(gen[2909]),

			.SO(gen[2967]),
			.S(gen[2968]),
			.SE(gen[2969]),

			.SELF(gen[2908]),
			.cell_state(gen[2908])
		); 

/******************* CELL 2909 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2909 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2848]),
			.N(gen[2849]),
			.NE(gen[2850]),

			.O(gen[2908]),
			.E(gen[2910]),

			.SO(gen[2968]),
			.S(gen[2969]),
			.SE(gen[2970]),

			.SELF(gen[2909]),
			.cell_state(gen[2909])
		); 

/******************* CELL 2910 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2910 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2849]),
			.N(gen[2850]),
			.NE(gen[2851]),

			.O(gen[2909]),
			.E(gen[2911]),

			.SO(gen[2969]),
			.S(gen[2970]),
			.SE(gen[2971]),

			.SELF(gen[2910]),
			.cell_state(gen[2910])
		); 

/******************* CELL 2911 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2911 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2850]),
			.N(gen[2851]),
			.NE(gen[2852]),

			.O(gen[2910]),
			.E(gen[2912]),

			.SO(gen[2970]),
			.S(gen[2971]),
			.SE(gen[2972]),

			.SELF(gen[2911]),
			.cell_state(gen[2911])
		); 

/******************* CELL 2912 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2912 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2851]),
			.N(gen[2852]),
			.NE(gen[2853]),

			.O(gen[2911]),
			.E(gen[2913]),

			.SO(gen[2971]),
			.S(gen[2972]),
			.SE(gen[2973]),

			.SELF(gen[2912]),
			.cell_state(gen[2912])
		); 

/******************* CELL 2913 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2913 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2852]),
			.N(gen[2853]),
			.NE(gen[2854]),

			.O(gen[2912]),
			.E(gen[2914]),

			.SO(gen[2972]),
			.S(gen[2973]),
			.SE(gen[2974]),

			.SELF(gen[2913]),
			.cell_state(gen[2913])
		); 

/******************* CELL 2914 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2914 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2853]),
			.N(gen[2854]),
			.NE(gen[2855]),

			.O(gen[2913]),
			.E(gen[2915]),

			.SO(gen[2973]),
			.S(gen[2974]),
			.SE(gen[2975]),

			.SELF(gen[2914]),
			.cell_state(gen[2914])
		); 

/******************* CELL 2915 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2915 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2854]),
			.N(gen[2855]),
			.NE(gen[2856]),

			.O(gen[2914]),
			.E(gen[2916]),

			.SO(gen[2974]),
			.S(gen[2975]),
			.SE(gen[2976]),

			.SELF(gen[2915]),
			.cell_state(gen[2915])
		); 

/******************* CELL 2916 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2916 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2855]),
			.N(gen[2856]),
			.NE(gen[2857]),

			.O(gen[2915]),
			.E(gen[2917]),

			.SO(gen[2975]),
			.S(gen[2976]),
			.SE(gen[2977]),

			.SELF(gen[2916]),
			.cell_state(gen[2916])
		); 

/******************* CELL 2917 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2917 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2856]),
			.N(gen[2857]),
			.NE(gen[2858]),

			.O(gen[2916]),
			.E(gen[2918]),

			.SO(gen[2976]),
			.S(gen[2977]),
			.SE(gen[2978]),

			.SELF(gen[2917]),
			.cell_state(gen[2917])
		); 

/******************* CELL 2918 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2918 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2857]),
			.N(gen[2858]),
			.NE(gen[2859]),

			.O(gen[2917]),
			.E(gen[2919]),

			.SO(gen[2977]),
			.S(gen[2978]),
			.SE(gen[2979]),

			.SELF(gen[2918]),
			.cell_state(gen[2918])
		); 

/******************* CELL 2919 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2919 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2858]),
			.N(gen[2859]),
			.NE(gen[2860]),

			.O(gen[2918]),
			.E(gen[2920]),

			.SO(gen[2978]),
			.S(gen[2979]),
			.SE(gen[2980]),

			.SELF(gen[2919]),
			.cell_state(gen[2919])
		); 

/******************* CELL 2920 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2920 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2859]),
			.N(gen[2860]),
			.NE(gen[2861]),

			.O(gen[2919]),
			.E(gen[2921]),

			.SO(gen[2979]),
			.S(gen[2980]),
			.SE(gen[2981]),

			.SELF(gen[2920]),
			.cell_state(gen[2920])
		); 

/******************* CELL 2921 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2921 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2860]),
			.N(gen[2861]),
			.NE(gen[2862]),

			.O(gen[2920]),
			.E(gen[2922]),

			.SO(gen[2980]),
			.S(gen[2981]),
			.SE(gen[2982]),

			.SELF(gen[2921]),
			.cell_state(gen[2921])
		); 

/******************* CELL 2922 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2922 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2861]),
			.N(gen[2862]),
			.NE(gen[2863]),

			.O(gen[2921]),
			.E(gen[2923]),

			.SO(gen[2981]),
			.S(gen[2982]),
			.SE(gen[2983]),

			.SELF(gen[2922]),
			.cell_state(gen[2922])
		); 

/******************* CELL 2923 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2923 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2862]),
			.N(gen[2863]),
			.NE(gen[2864]),

			.O(gen[2922]),
			.E(gen[2924]),

			.SO(gen[2982]),
			.S(gen[2983]),
			.SE(gen[2984]),

			.SELF(gen[2923]),
			.cell_state(gen[2923])
		); 

/******************* CELL 2924 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2924 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2863]),
			.N(gen[2864]),
			.NE(gen[2865]),

			.O(gen[2923]),
			.E(gen[2925]),

			.SO(gen[2983]),
			.S(gen[2984]),
			.SE(gen[2985]),

			.SELF(gen[2924]),
			.cell_state(gen[2924])
		); 

/******************* CELL 2925 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2925 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2864]),
			.N(gen[2865]),
			.NE(gen[2866]),

			.O(gen[2924]),
			.E(gen[2926]),

			.SO(gen[2984]),
			.S(gen[2985]),
			.SE(gen[2986]),

			.SELF(gen[2925]),
			.cell_state(gen[2925])
		); 

/******************* CELL 2926 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2926 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2865]),
			.N(gen[2866]),
			.NE(gen[2867]),

			.O(gen[2925]),
			.E(gen[2927]),

			.SO(gen[2985]),
			.S(gen[2986]),
			.SE(gen[2987]),

			.SELF(gen[2926]),
			.cell_state(gen[2926])
		); 

/******************* CELL 2927 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2927 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2866]),
			.N(gen[2867]),
			.NE(gen[2868]),

			.O(gen[2926]),
			.E(gen[2928]),

			.SO(gen[2986]),
			.S(gen[2987]),
			.SE(gen[2988]),

			.SELF(gen[2927]),
			.cell_state(gen[2927])
		); 

/******************* CELL 2928 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2928 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2867]),
			.N(gen[2868]),
			.NE(gen[2869]),

			.O(gen[2927]),
			.E(gen[2929]),

			.SO(gen[2987]),
			.S(gen[2988]),
			.SE(gen[2989]),

			.SELF(gen[2928]),
			.cell_state(gen[2928])
		); 

/******************* CELL 2929 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2929 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2868]),
			.N(gen[2869]),
			.NE(gen[2870]),

			.O(gen[2928]),
			.E(gen[2930]),

			.SO(gen[2988]),
			.S(gen[2989]),
			.SE(gen[2990]),

			.SELF(gen[2929]),
			.cell_state(gen[2929])
		); 

/******************* CELL 2930 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2930 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2869]),
			.N(gen[2870]),
			.NE(gen[2871]),

			.O(gen[2929]),
			.E(gen[2931]),

			.SO(gen[2989]),
			.S(gen[2990]),
			.SE(gen[2991]),

			.SELF(gen[2930]),
			.cell_state(gen[2930])
		); 

/******************* CELL 2931 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2931 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2870]),
			.N(gen[2871]),
			.NE(gen[2872]),

			.O(gen[2930]),
			.E(gen[2932]),

			.SO(gen[2990]),
			.S(gen[2991]),
			.SE(gen[2992]),

			.SELF(gen[2931]),
			.cell_state(gen[2931])
		); 

/******************* CELL 2932 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2932 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2871]),
			.N(gen[2872]),
			.NE(gen[2873]),

			.O(gen[2931]),
			.E(gen[2933]),

			.SO(gen[2991]),
			.S(gen[2992]),
			.SE(gen[2993]),

			.SELF(gen[2932]),
			.cell_state(gen[2932])
		); 

/******************* CELL 2933 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2933 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2872]),
			.N(gen[2873]),
			.NE(gen[2874]),

			.O(gen[2932]),
			.E(gen[2934]),

			.SO(gen[2992]),
			.S(gen[2993]),
			.SE(gen[2994]),

			.SELF(gen[2933]),
			.cell_state(gen[2933])
		); 

/******************* CELL 2934 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2934 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2873]),
			.N(gen[2874]),
			.NE(gen[2875]),

			.O(gen[2933]),
			.E(gen[2935]),

			.SO(gen[2993]),
			.S(gen[2994]),
			.SE(gen[2995]),

			.SELF(gen[2934]),
			.cell_state(gen[2934])
		); 

/******************* CELL 2935 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2935 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2874]),
			.N(gen[2875]),
			.NE(gen[2876]),

			.O(gen[2934]),
			.E(gen[2936]),

			.SO(gen[2994]),
			.S(gen[2995]),
			.SE(gen[2996]),

			.SELF(gen[2935]),
			.cell_state(gen[2935])
		); 

/******************* CELL 2936 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2936 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2875]),
			.N(gen[2876]),
			.NE(gen[2877]),

			.O(gen[2935]),
			.E(gen[2937]),

			.SO(gen[2995]),
			.S(gen[2996]),
			.SE(gen[2997]),

			.SELF(gen[2936]),
			.cell_state(gen[2936])
		); 

/******************* CELL 2937 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2937 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2876]),
			.N(gen[2877]),
			.NE(gen[2878]),

			.O(gen[2936]),
			.E(gen[2938]),

			.SO(gen[2996]),
			.S(gen[2997]),
			.SE(gen[2998]),

			.SELF(gen[2937]),
			.cell_state(gen[2937])
		); 

/******************* CELL 2938 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2938 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2877]),
			.N(gen[2878]),
			.NE(gen[2879]),

			.O(gen[2937]),
			.E(gen[2939]),

			.SO(gen[2997]),
			.S(gen[2998]),
			.SE(gen[2999]),

			.SELF(gen[2938]),
			.cell_state(gen[2938])
		); 

/******************* CELL 2939 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2939 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2878]),
			.N(gen[2879]),
			.NE(gen[2878]),

			.O(gen[2938]),
			.E(gen[2938]),

			.SO(gen[2998]),
			.S(gen[2999]),
			.SE(gen[2998]),

			.SELF(gen[2939]),
			.cell_state(gen[2939])
		); 

/******************* CELL 2940 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2940 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2881]),
			.N(gen[2880]),
			.NE(gen[2881]),

			.O(gen[2941]),
			.E(gen[2941]),

			.SO(gen[3001]),
			.S(gen[3000]),
			.SE(gen[3001]),

			.SELF(gen[2940]),
			.cell_state(gen[2940])
		); 

/******************* CELL 2941 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2941 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2880]),
			.N(gen[2881]),
			.NE(gen[2882]),

			.O(gen[2940]),
			.E(gen[2942]),

			.SO(gen[3000]),
			.S(gen[3001]),
			.SE(gen[3002]),

			.SELF(gen[2941]),
			.cell_state(gen[2941])
		); 

/******************* CELL 2942 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2942 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2881]),
			.N(gen[2882]),
			.NE(gen[2883]),

			.O(gen[2941]),
			.E(gen[2943]),

			.SO(gen[3001]),
			.S(gen[3002]),
			.SE(gen[3003]),

			.SELF(gen[2942]),
			.cell_state(gen[2942])
		); 

/******************* CELL 2943 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2943 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2882]),
			.N(gen[2883]),
			.NE(gen[2884]),

			.O(gen[2942]),
			.E(gen[2944]),

			.SO(gen[3002]),
			.S(gen[3003]),
			.SE(gen[3004]),

			.SELF(gen[2943]),
			.cell_state(gen[2943])
		); 

/******************* CELL 2944 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2944 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2883]),
			.N(gen[2884]),
			.NE(gen[2885]),

			.O(gen[2943]),
			.E(gen[2945]),

			.SO(gen[3003]),
			.S(gen[3004]),
			.SE(gen[3005]),

			.SELF(gen[2944]),
			.cell_state(gen[2944])
		); 

/******************* CELL 2945 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2945 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2884]),
			.N(gen[2885]),
			.NE(gen[2886]),

			.O(gen[2944]),
			.E(gen[2946]),

			.SO(gen[3004]),
			.S(gen[3005]),
			.SE(gen[3006]),

			.SELF(gen[2945]),
			.cell_state(gen[2945])
		); 

/******************* CELL 2946 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2946 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2885]),
			.N(gen[2886]),
			.NE(gen[2887]),

			.O(gen[2945]),
			.E(gen[2947]),

			.SO(gen[3005]),
			.S(gen[3006]),
			.SE(gen[3007]),

			.SELF(gen[2946]),
			.cell_state(gen[2946])
		); 

/******************* CELL 2947 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2947 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2886]),
			.N(gen[2887]),
			.NE(gen[2888]),

			.O(gen[2946]),
			.E(gen[2948]),

			.SO(gen[3006]),
			.S(gen[3007]),
			.SE(gen[3008]),

			.SELF(gen[2947]),
			.cell_state(gen[2947])
		); 

/******************* CELL 2948 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2948 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2887]),
			.N(gen[2888]),
			.NE(gen[2889]),

			.O(gen[2947]),
			.E(gen[2949]),

			.SO(gen[3007]),
			.S(gen[3008]),
			.SE(gen[3009]),

			.SELF(gen[2948]),
			.cell_state(gen[2948])
		); 

/******************* CELL 2949 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2949 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2888]),
			.N(gen[2889]),
			.NE(gen[2890]),

			.O(gen[2948]),
			.E(gen[2950]),

			.SO(gen[3008]),
			.S(gen[3009]),
			.SE(gen[3010]),

			.SELF(gen[2949]),
			.cell_state(gen[2949])
		); 

/******************* CELL 2950 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2950 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2889]),
			.N(gen[2890]),
			.NE(gen[2891]),

			.O(gen[2949]),
			.E(gen[2951]),

			.SO(gen[3009]),
			.S(gen[3010]),
			.SE(gen[3011]),

			.SELF(gen[2950]),
			.cell_state(gen[2950])
		); 

/******************* CELL 2951 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2951 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2890]),
			.N(gen[2891]),
			.NE(gen[2892]),

			.O(gen[2950]),
			.E(gen[2952]),

			.SO(gen[3010]),
			.S(gen[3011]),
			.SE(gen[3012]),

			.SELF(gen[2951]),
			.cell_state(gen[2951])
		); 

/******************* CELL 2952 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2952 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2891]),
			.N(gen[2892]),
			.NE(gen[2893]),

			.O(gen[2951]),
			.E(gen[2953]),

			.SO(gen[3011]),
			.S(gen[3012]),
			.SE(gen[3013]),

			.SELF(gen[2952]),
			.cell_state(gen[2952])
		); 

/******************* CELL 2953 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2953 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2892]),
			.N(gen[2893]),
			.NE(gen[2894]),

			.O(gen[2952]),
			.E(gen[2954]),

			.SO(gen[3012]),
			.S(gen[3013]),
			.SE(gen[3014]),

			.SELF(gen[2953]),
			.cell_state(gen[2953])
		); 

/******************* CELL 2954 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2954 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2893]),
			.N(gen[2894]),
			.NE(gen[2895]),

			.O(gen[2953]),
			.E(gen[2955]),

			.SO(gen[3013]),
			.S(gen[3014]),
			.SE(gen[3015]),

			.SELF(gen[2954]),
			.cell_state(gen[2954])
		); 

/******************* CELL 2955 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2955 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2894]),
			.N(gen[2895]),
			.NE(gen[2896]),

			.O(gen[2954]),
			.E(gen[2956]),

			.SO(gen[3014]),
			.S(gen[3015]),
			.SE(gen[3016]),

			.SELF(gen[2955]),
			.cell_state(gen[2955])
		); 

/******************* CELL 2956 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2956 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2895]),
			.N(gen[2896]),
			.NE(gen[2897]),

			.O(gen[2955]),
			.E(gen[2957]),

			.SO(gen[3015]),
			.S(gen[3016]),
			.SE(gen[3017]),

			.SELF(gen[2956]),
			.cell_state(gen[2956])
		); 

/******************* CELL 2957 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2957 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2896]),
			.N(gen[2897]),
			.NE(gen[2898]),

			.O(gen[2956]),
			.E(gen[2958]),

			.SO(gen[3016]),
			.S(gen[3017]),
			.SE(gen[3018]),

			.SELF(gen[2957]),
			.cell_state(gen[2957])
		); 

/******************* CELL 2958 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2958 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2897]),
			.N(gen[2898]),
			.NE(gen[2899]),

			.O(gen[2957]),
			.E(gen[2959]),

			.SO(gen[3017]),
			.S(gen[3018]),
			.SE(gen[3019]),

			.SELF(gen[2958]),
			.cell_state(gen[2958])
		); 

/******************* CELL 2959 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2959 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2898]),
			.N(gen[2899]),
			.NE(gen[2900]),

			.O(gen[2958]),
			.E(gen[2960]),

			.SO(gen[3018]),
			.S(gen[3019]),
			.SE(gen[3020]),

			.SELF(gen[2959]),
			.cell_state(gen[2959])
		); 

/******************* CELL 2960 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2960 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2899]),
			.N(gen[2900]),
			.NE(gen[2901]),

			.O(gen[2959]),
			.E(gen[2961]),

			.SO(gen[3019]),
			.S(gen[3020]),
			.SE(gen[3021]),

			.SELF(gen[2960]),
			.cell_state(gen[2960])
		); 

/******************* CELL 2961 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2961 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2900]),
			.N(gen[2901]),
			.NE(gen[2902]),

			.O(gen[2960]),
			.E(gen[2962]),

			.SO(gen[3020]),
			.S(gen[3021]),
			.SE(gen[3022]),

			.SELF(gen[2961]),
			.cell_state(gen[2961])
		); 

/******************* CELL 2962 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2962 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2901]),
			.N(gen[2902]),
			.NE(gen[2903]),

			.O(gen[2961]),
			.E(gen[2963]),

			.SO(gen[3021]),
			.S(gen[3022]),
			.SE(gen[3023]),

			.SELF(gen[2962]),
			.cell_state(gen[2962])
		); 

/******************* CELL 2963 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2963 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2902]),
			.N(gen[2903]),
			.NE(gen[2904]),

			.O(gen[2962]),
			.E(gen[2964]),

			.SO(gen[3022]),
			.S(gen[3023]),
			.SE(gen[3024]),

			.SELF(gen[2963]),
			.cell_state(gen[2963])
		); 

/******************* CELL 2964 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2964 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2903]),
			.N(gen[2904]),
			.NE(gen[2905]),

			.O(gen[2963]),
			.E(gen[2965]),

			.SO(gen[3023]),
			.S(gen[3024]),
			.SE(gen[3025]),

			.SELF(gen[2964]),
			.cell_state(gen[2964])
		); 

/******************* CELL 2965 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2965 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2904]),
			.N(gen[2905]),
			.NE(gen[2906]),

			.O(gen[2964]),
			.E(gen[2966]),

			.SO(gen[3024]),
			.S(gen[3025]),
			.SE(gen[3026]),

			.SELF(gen[2965]),
			.cell_state(gen[2965])
		); 

/******************* CELL 2966 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2966 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2905]),
			.N(gen[2906]),
			.NE(gen[2907]),

			.O(gen[2965]),
			.E(gen[2967]),

			.SO(gen[3025]),
			.S(gen[3026]),
			.SE(gen[3027]),

			.SELF(gen[2966]),
			.cell_state(gen[2966])
		); 

/******************* CELL 2967 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2967 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2906]),
			.N(gen[2907]),
			.NE(gen[2908]),

			.O(gen[2966]),
			.E(gen[2968]),

			.SO(gen[3026]),
			.S(gen[3027]),
			.SE(gen[3028]),

			.SELF(gen[2967]),
			.cell_state(gen[2967])
		); 

/******************* CELL 2968 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2968 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2907]),
			.N(gen[2908]),
			.NE(gen[2909]),

			.O(gen[2967]),
			.E(gen[2969]),

			.SO(gen[3027]),
			.S(gen[3028]),
			.SE(gen[3029]),

			.SELF(gen[2968]),
			.cell_state(gen[2968])
		); 

/******************* CELL 2969 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2969 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2908]),
			.N(gen[2909]),
			.NE(gen[2910]),

			.O(gen[2968]),
			.E(gen[2970]),

			.SO(gen[3028]),
			.S(gen[3029]),
			.SE(gen[3030]),

			.SELF(gen[2969]),
			.cell_state(gen[2969])
		); 

/******************* CELL 2970 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2970 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2909]),
			.N(gen[2910]),
			.NE(gen[2911]),

			.O(gen[2969]),
			.E(gen[2971]),

			.SO(gen[3029]),
			.S(gen[3030]),
			.SE(gen[3031]),

			.SELF(gen[2970]),
			.cell_state(gen[2970])
		); 

/******************* CELL 2971 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2971 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2910]),
			.N(gen[2911]),
			.NE(gen[2912]),

			.O(gen[2970]),
			.E(gen[2972]),

			.SO(gen[3030]),
			.S(gen[3031]),
			.SE(gen[3032]),

			.SELF(gen[2971]),
			.cell_state(gen[2971])
		); 

/******************* CELL 2972 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2972 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2911]),
			.N(gen[2912]),
			.NE(gen[2913]),

			.O(gen[2971]),
			.E(gen[2973]),

			.SO(gen[3031]),
			.S(gen[3032]),
			.SE(gen[3033]),

			.SELF(gen[2972]),
			.cell_state(gen[2972])
		); 

/******************* CELL 2973 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2973 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2912]),
			.N(gen[2913]),
			.NE(gen[2914]),

			.O(gen[2972]),
			.E(gen[2974]),

			.SO(gen[3032]),
			.S(gen[3033]),
			.SE(gen[3034]),

			.SELF(gen[2973]),
			.cell_state(gen[2973])
		); 

/******************* CELL 2974 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2974 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2913]),
			.N(gen[2914]),
			.NE(gen[2915]),

			.O(gen[2973]),
			.E(gen[2975]),

			.SO(gen[3033]),
			.S(gen[3034]),
			.SE(gen[3035]),

			.SELF(gen[2974]),
			.cell_state(gen[2974])
		); 

/******************* CELL 2975 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2975 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2914]),
			.N(gen[2915]),
			.NE(gen[2916]),

			.O(gen[2974]),
			.E(gen[2976]),

			.SO(gen[3034]),
			.S(gen[3035]),
			.SE(gen[3036]),

			.SELF(gen[2975]),
			.cell_state(gen[2975])
		); 

/******************* CELL 2976 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2976 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2915]),
			.N(gen[2916]),
			.NE(gen[2917]),

			.O(gen[2975]),
			.E(gen[2977]),

			.SO(gen[3035]),
			.S(gen[3036]),
			.SE(gen[3037]),

			.SELF(gen[2976]),
			.cell_state(gen[2976])
		); 

/******************* CELL 2977 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2977 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2916]),
			.N(gen[2917]),
			.NE(gen[2918]),

			.O(gen[2976]),
			.E(gen[2978]),

			.SO(gen[3036]),
			.S(gen[3037]),
			.SE(gen[3038]),

			.SELF(gen[2977]),
			.cell_state(gen[2977])
		); 

/******************* CELL 2978 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2978 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2917]),
			.N(gen[2918]),
			.NE(gen[2919]),

			.O(gen[2977]),
			.E(gen[2979]),

			.SO(gen[3037]),
			.S(gen[3038]),
			.SE(gen[3039]),

			.SELF(gen[2978]),
			.cell_state(gen[2978])
		); 

/******************* CELL 2979 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2979 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2918]),
			.N(gen[2919]),
			.NE(gen[2920]),

			.O(gen[2978]),
			.E(gen[2980]),

			.SO(gen[3038]),
			.S(gen[3039]),
			.SE(gen[3040]),

			.SELF(gen[2979]),
			.cell_state(gen[2979])
		); 

/******************* CELL 2980 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2980 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2919]),
			.N(gen[2920]),
			.NE(gen[2921]),

			.O(gen[2979]),
			.E(gen[2981]),

			.SO(gen[3039]),
			.S(gen[3040]),
			.SE(gen[3041]),

			.SELF(gen[2980]),
			.cell_state(gen[2980])
		); 

/******************* CELL 2981 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2981 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2920]),
			.N(gen[2921]),
			.NE(gen[2922]),

			.O(gen[2980]),
			.E(gen[2982]),

			.SO(gen[3040]),
			.S(gen[3041]),
			.SE(gen[3042]),

			.SELF(gen[2981]),
			.cell_state(gen[2981])
		); 

/******************* CELL 2982 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2982 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2921]),
			.N(gen[2922]),
			.NE(gen[2923]),

			.O(gen[2981]),
			.E(gen[2983]),

			.SO(gen[3041]),
			.S(gen[3042]),
			.SE(gen[3043]),

			.SELF(gen[2982]),
			.cell_state(gen[2982])
		); 

/******************* CELL 2983 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2983 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2922]),
			.N(gen[2923]),
			.NE(gen[2924]),

			.O(gen[2982]),
			.E(gen[2984]),

			.SO(gen[3042]),
			.S(gen[3043]),
			.SE(gen[3044]),

			.SELF(gen[2983]),
			.cell_state(gen[2983])
		); 

/******************* CELL 2984 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2984 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2923]),
			.N(gen[2924]),
			.NE(gen[2925]),

			.O(gen[2983]),
			.E(gen[2985]),

			.SO(gen[3043]),
			.S(gen[3044]),
			.SE(gen[3045]),

			.SELF(gen[2984]),
			.cell_state(gen[2984])
		); 

/******************* CELL 2985 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2985 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2924]),
			.N(gen[2925]),
			.NE(gen[2926]),

			.O(gen[2984]),
			.E(gen[2986]),

			.SO(gen[3044]),
			.S(gen[3045]),
			.SE(gen[3046]),

			.SELF(gen[2985]),
			.cell_state(gen[2985])
		); 

/******************* CELL 2986 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2986 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2925]),
			.N(gen[2926]),
			.NE(gen[2927]),

			.O(gen[2985]),
			.E(gen[2987]),

			.SO(gen[3045]),
			.S(gen[3046]),
			.SE(gen[3047]),

			.SELF(gen[2986]),
			.cell_state(gen[2986])
		); 

/******************* CELL 2987 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2987 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2926]),
			.N(gen[2927]),
			.NE(gen[2928]),

			.O(gen[2986]),
			.E(gen[2988]),

			.SO(gen[3046]),
			.S(gen[3047]),
			.SE(gen[3048]),

			.SELF(gen[2987]),
			.cell_state(gen[2987])
		); 

/******************* CELL 2988 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2988 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2927]),
			.N(gen[2928]),
			.NE(gen[2929]),

			.O(gen[2987]),
			.E(gen[2989]),

			.SO(gen[3047]),
			.S(gen[3048]),
			.SE(gen[3049]),

			.SELF(gen[2988]),
			.cell_state(gen[2988])
		); 

/******************* CELL 2989 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2989 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2928]),
			.N(gen[2929]),
			.NE(gen[2930]),

			.O(gen[2988]),
			.E(gen[2990]),

			.SO(gen[3048]),
			.S(gen[3049]),
			.SE(gen[3050]),

			.SELF(gen[2989]),
			.cell_state(gen[2989])
		); 

/******************* CELL 2990 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2990 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2929]),
			.N(gen[2930]),
			.NE(gen[2931]),

			.O(gen[2989]),
			.E(gen[2991]),

			.SO(gen[3049]),
			.S(gen[3050]),
			.SE(gen[3051]),

			.SELF(gen[2990]),
			.cell_state(gen[2990])
		); 

/******************* CELL 2991 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2991 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2930]),
			.N(gen[2931]),
			.NE(gen[2932]),

			.O(gen[2990]),
			.E(gen[2992]),

			.SO(gen[3050]),
			.S(gen[3051]),
			.SE(gen[3052]),

			.SELF(gen[2991]),
			.cell_state(gen[2991])
		); 

/******************* CELL 2992 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2992 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2931]),
			.N(gen[2932]),
			.NE(gen[2933]),

			.O(gen[2991]),
			.E(gen[2993]),

			.SO(gen[3051]),
			.S(gen[3052]),
			.SE(gen[3053]),

			.SELF(gen[2992]),
			.cell_state(gen[2992])
		); 

/******************* CELL 2993 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2993 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2932]),
			.N(gen[2933]),
			.NE(gen[2934]),

			.O(gen[2992]),
			.E(gen[2994]),

			.SO(gen[3052]),
			.S(gen[3053]),
			.SE(gen[3054]),

			.SELF(gen[2993]),
			.cell_state(gen[2993])
		); 

/******************* CELL 2994 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2994 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2933]),
			.N(gen[2934]),
			.NE(gen[2935]),

			.O(gen[2993]),
			.E(gen[2995]),

			.SO(gen[3053]),
			.S(gen[3054]),
			.SE(gen[3055]),

			.SELF(gen[2994]),
			.cell_state(gen[2994])
		); 

/******************* CELL 2995 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2995 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2934]),
			.N(gen[2935]),
			.NE(gen[2936]),

			.O(gen[2994]),
			.E(gen[2996]),

			.SO(gen[3054]),
			.S(gen[3055]),
			.SE(gen[3056]),

			.SELF(gen[2995]),
			.cell_state(gen[2995])
		); 

/******************* CELL 2996 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2996 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2935]),
			.N(gen[2936]),
			.NE(gen[2937]),

			.O(gen[2995]),
			.E(gen[2997]),

			.SO(gen[3055]),
			.S(gen[3056]),
			.SE(gen[3057]),

			.SELF(gen[2996]),
			.cell_state(gen[2996])
		); 

/******************* CELL 2997 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2997 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2936]),
			.N(gen[2937]),
			.NE(gen[2938]),

			.O(gen[2996]),
			.E(gen[2998]),

			.SO(gen[3056]),
			.S(gen[3057]),
			.SE(gen[3058]),

			.SELF(gen[2997]),
			.cell_state(gen[2997])
		); 

/******************* CELL 2998 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2998 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2937]),
			.N(gen[2938]),
			.NE(gen[2939]),

			.O(gen[2997]),
			.E(gen[2999]),

			.SO(gen[3057]),
			.S(gen[3058]),
			.SE(gen[3059]),

			.SELF(gen[2998]),
			.cell_state(gen[2998])
		); 

/******************* CELL 2999 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell2999 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2938]),
			.N(gen[2939]),
			.NE(gen[2938]),

			.O(gen[2998]),
			.E(gen[2998]),

			.SO(gen[3058]),
			.S(gen[3059]),
			.SE(gen[3058]),

			.SELF(gen[2999]),
			.cell_state(gen[2999])
		); 

/******************* CELL 3000 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3000 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2941]),
			.N(gen[2940]),
			.NE(gen[2941]),

			.O(gen[3001]),
			.E(gen[3001]),

			.SO(gen[3061]),
			.S(gen[3060]),
			.SE(gen[3061]),

			.SELF(gen[3000]),
			.cell_state(gen[3000])
		); 

/******************* CELL 3001 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3001 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2940]),
			.N(gen[2941]),
			.NE(gen[2942]),

			.O(gen[3000]),
			.E(gen[3002]),

			.SO(gen[3060]),
			.S(gen[3061]),
			.SE(gen[3062]),

			.SELF(gen[3001]),
			.cell_state(gen[3001])
		); 

/******************* CELL 3002 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3002 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2941]),
			.N(gen[2942]),
			.NE(gen[2943]),

			.O(gen[3001]),
			.E(gen[3003]),

			.SO(gen[3061]),
			.S(gen[3062]),
			.SE(gen[3063]),

			.SELF(gen[3002]),
			.cell_state(gen[3002])
		); 

/******************* CELL 3003 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3003 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2942]),
			.N(gen[2943]),
			.NE(gen[2944]),

			.O(gen[3002]),
			.E(gen[3004]),

			.SO(gen[3062]),
			.S(gen[3063]),
			.SE(gen[3064]),

			.SELF(gen[3003]),
			.cell_state(gen[3003])
		); 

/******************* CELL 3004 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3004 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2943]),
			.N(gen[2944]),
			.NE(gen[2945]),

			.O(gen[3003]),
			.E(gen[3005]),

			.SO(gen[3063]),
			.S(gen[3064]),
			.SE(gen[3065]),

			.SELF(gen[3004]),
			.cell_state(gen[3004])
		); 

/******************* CELL 3005 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3005 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2944]),
			.N(gen[2945]),
			.NE(gen[2946]),

			.O(gen[3004]),
			.E(gen[3006]),

			.SO(gen[3064]),
			.S(gen[3065]),
			.SE(gen[3066]),

			.SELF(gen[3005]),
			.cell_state(gen[3005])
		); 

/******************* CELL 3006 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3006 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2945]),
			.N(gen[2946]),
			.NE(gen[2947]),

			.O(gen[3005]),
			.E(gen[3007]),

			.SO(gen[3065]),
			.S(gen[3066]),
			.SE(gen[3067]),

			.SELF(gen[3006]),
			.cell_state(gen[3006])
		); 

/******************* CELL 3007 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3007 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2946]),
			.N(gen[2947]),
			.NE(gen[2948]),

			.O(gen[3006]),
			.E(gen[3008]),

			.SO(gen[3066]),
			.S(gen[3067]),
			.SE(gen[3068]),

			.SELF(gen[3007]),
			.cell_state(gen[3007])
		); 

/******************* CELL 3008 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3008 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2947]),
			.N(gen[2948]),
			.NE(gen[2949]),

			.O(gen[3007]),
			.E(gen[3009]),

			.SO(gen[3067]),
			.S(gen[3068]),
			.SE(gen[3069]),

			.SELF(gen[3008]),
			.cell_state(gen[3008])
		); 

/******************* CELL 3009 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3009 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2948]),
			.N(gen[2949]),
			.NE(gen[2950]),

			.O(gen[3008]),
			.E(gen[3010]),

			.SO(gen[3068]),
			.S(gen[3069]),
			.SE(gen[3070]),

			.SELF(gen[3009]),
			.cell_state(gen[3009])
		); 

/******************* CELL 3010 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3010 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2949]),
			.N(gen[2950]),
			.NE(gen[2951]),

			.O(gen[3009]),
			.E(gen[3011]),

			.SO(gen[3069]),
			.S(gen[3070]),
			.SE(gen[3071]),

			.SELF(gen[3010]),
			.cell_state(gen[3010])
		); 

/******************* CELL 3011 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3011 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2950]),
			.N(gen[2951]),
			.NE(gen[2952]),

			.O(gen[3010]),
			.E(gen[3012]),

			.SO(gen[3070]),
			.S(gen[3071]),
			.SE(gen[3072]),

			.SELF(gen[3011]),
			.cell_state(gen[3011])
		); 

/******************* CELL 3012 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3012 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2951]),
			.N(gen[2952]),
			.NE(gen[2953]),

			.O(gen[3011]),
			.E(gen[3013]),

			.SO(gen[3071]),
			.S(gen[3072]),
			.SE(gen[3073]),

			.SELF(gen[3012]),
			.cell_state(gen[3012])
		); 

/******************* CELL 3013 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3013 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2952]),
			.N(gen[2953]),
			.NE(gen[2954]),

			.O(gen[3012]),
			.E(gen[3014]),

			.SO(gen[3072]),
			.S(gen[3073]),
			.SE(gen[3074]),

			.SELF(gen[3013]),
			.cell_state(gen[3013])
		); 

/******************* CELL 3014 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3014 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2953]),
			.N(gen[2954]),
			.NE(gen[2955]),

			.O(gen[3013]),
			.E(gen[3015]),

			.SO(gen[3073]),
			.S(gen[3074]),
			.SE(gen[3075]),

			.SELF(gen[3014]),
			.cell_state(gen[3014])
		); 

/******************* CELL 3015 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3015 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2954]),
			.N(gen[2955]),
			.NE(gen[2956]),

			.O(gen[3014]),
			.E(gen[3016]),

			.SO(gen[3074]),
			.S(gen[3075]),
			.SE(gen[3076]),

			.SELF(gen[3015]),
			.cell_state(gen[3015])
		); 

/******************* CELL 3016 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3016 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2955]),
			.N(gen[2956]),
			.NE(gen[2957]),

			.O(gen[3015]),
			.E(gen[3017]),

			.SO(gen[3075]),
			.S(gen[3076]),
			.SE(gen[3077]),

			.SELF(gen[3016]),
			.cell_state(gen[3016])
		); 

/******************* CELL 3017 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3017 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2956]),
			.N(gen[2957]),
			.NE(gen[2958]),

			.O(gen[3016]),
			.E(gen[3018]),

			.SO(gen[3076]),
			.S(gen[3077]),
			.SE(gen[3078]),

			.SELF(gen[3017]),
			.cell_state(gen[3017])
		); 

/******************* CELL 3018 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3018 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2957]),
			.N(gen[2958]),
			.NE(gen[2959]),

			.O(gen[3017]),
			.E(gen[3019]),

			.SO(gen[3077]),
			.S(gen[3078]),
			.SE(gen[3079]),

			.SELF(gen[3018]),
			.cell_state(gen[3018])
		); 

/******************* CELL 3019 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3019 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2958]),
			.N(gen[2959]),
			.NE(gen[2960]),

			.O(gen[3018]),
			.E(gen[3020]),

			.SO(gen[3078]),
			.S(gen[3079]),
			.SE(gen[3080]),

			.SELF(gen[3019]),
			.cell_state(gen[3019])
		); 

/******************* CELL 3020 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3020 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2959]),
			.N(gen[2960]),
			.NE(gen[2961]),

			.O(gen[3019]),
			.E(gen[3021]),

			.SO(gen[3079]),
			.S(gen[3080]),
			.SE(gen[3081]),

			.SELF(gen[3020]),
			.cell_state(gen[3020])
		); 

/******************* CELL 3021 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3021 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2960]),
			.N(gen[2961]),
			.NE(gen[2962]),

			.O(gen[3020]),
			.E(gen[3022]),

			.SO(gen[3080]),
			.S(gen[3081]),
			.SE(gen[3082]),

			.SELF(gen[3021]),
			.cell_state(gen[3021])
		); 

/******************* CELL 3022 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3022 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2961]),
			.N(gen[2962]),
			.NE(gen[2963]),

			.O(gen[3021]),
			.E(gen[3023]),

			.SO(gen[3081]),
			.S(gen[3082]),
			.SE(gen[3083]),

			.SELF(gen[3022]),
			.cell_state(gen[3022])
		); 

/******************* CELL 3023 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3023 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2962]),
			.N(gen[2963]),
			.NE(gen[2964]),

			.O(gen[3022]),
			.E(gen[3024]),

			.SO(gen[3082]),
			.S(gen[3083]),
			.SE(gen[3084]),

			.SELF(gen[3023]),
			.cell_state(gen[3023])
		); 

/******************* CELL 3024 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3024 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2963]),
			.N(gen[2964]),
			.NE(gen[2965]),

			.O(gen[3023]),
			.E(gen[3025]),

			.SO(gen[3083]),
			.S(gen[3084]),
			.SE(gen[3085]),

			.SELF(gen[3024]),
			.cell_state(gen[3024])
		); 

/******************* CELL 3025 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3025 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2964]),
			.N(gen[2965]),
			.NE(gen[2966]),

			.O(gen[3024]),
			.E(gen[3026]),

			.SO(gen[3084]),
			.S(gen[3085]),
			.SE(gen[3086]),

			.SELF(gen[3025]),
			.cell_state(gen[3025])
		); 

/******************* CELL 3026 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3026 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2965]),
			.N(gen[2966]),
			.NE(gen[2967]),

			.O(gen[3025]),
			.E(gen[3027]),

			.SO(gen[3085]),
			.S(gen[3086]),
			.SE(gen[3087]),

			.SELF(gen[3026]),
			.cell_state(gen[3026])
		); 

/******************* CELL 3027 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3027 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2966]),
			.N(gen[2967]),
			.NE(gen[2968]),

			.O(gen[3026]),
			.E(gen[3028]),

			.SO(gen[3086]),
			.S(gen[3087]),
			.SE(gen[3088]),

			.SELF(gen[3027]),
			.cell_state(gen[3027])
		); 

/******************* CELL 3028 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3028 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2967]),
			.N(gen[2968]),
			.NE(gen[2969]),

			.O(gen[3027]),
			.E(gen[3029]),

			.SO(gen[3087]),
			.S(gen[3088]),
			.SE(gen[3089]),

			.SELF(gen[3028]),
			.cell_state(gen[3028])
		); 

/******************* CELL 3029 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3029 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2968]),
			.N(gen[2969]),
			.NE(gen[2970]),

			.O(gen[3028]),
			.E(gen[3030]),

			.SO(gen[3088]),
			.S(gen[3089]),
			.SE(gen[3090]),

			.SELF(gen[3029]),
			.cell_state(gen[3029])
		); 

/******************* CELL 3030 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3030 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2969]),
			.N(gen[2970]),
			.NE(gen[2971]),

			.O(gen[3029]),
			.E(gen[3031]),

			.SO(gen[3089]),
			.S(gen[3090]),
			.SE(gen[3091]),

			.SELF(gen[3030]),
			.cell_state(gen[3030])
		); 

/******************* CELL 3031 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3031 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2970]),
			.N(gen[2971]),
			.NE(gen[2972]),

			.O(gen[3030]),
			.E(gen[3032]),

			.SO(gen[3090]),
			.S(gen[3091]),
			.SE(gen[3092]),

			.SELF(gen[3031]),
			.cell_state(gen[3031])
		); 

/******************* CELL 3032 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3032 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2971]),
			.N(gen[2972]),
			.NE(gen[2973]),

			.O(gen[3031]),
			.E(gen[3033]),

			.SO(gen[3091]),
			.S(gen[3092]),
			.SE(gen[3093]),

			.SELF(gen[3032]),
			.cell_state(gen[3032])
		); 

/******************* CELL 3033 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3033 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2972]),
			.N(gen[2973]),
			.NE(gen[2974]),

			.O(gen[3032]),
			.E(gen[3034]),

			.SO(gen[3092]),
			.S(gen[3093]),
			.SE(gen[3094]),

			.SELF(gen[3033]),
			.cell_state(gen[3033])
		); 

/******************* CELL 3034 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3034 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2973]),
			.N(gen[2974]),
			.NE(gen[2975]),

			.O(gen[3033]),
			.E(gen[3035]),

			.SO(gen[3093]),
			.S(gen[3094]),
			.SE(gen[3095]),

			.SELF(gen[3034]),
			.cell_state(gen[3034])
		); 

/******************* CELL 3035 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3035 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2974]),
			.N(gen[2975]),
			.NE(gen[2976]),

			.O(gen[3034]),
			.E(gen[3036]),

			.SO(gen[3094]),
			.S(gen[3095]),
			.SE(gen[3096]),

			.SELF(gen[3035]),
			.cell_state(gen[3035])
		); 

/******************* CELL 3036 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3036 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2975]),
			.N(gen[2976]),
			.NE(gen[2977]),

			.O(gen[3035]),
			.E(gen[3037]),

			.SO(gen[3095]),
			.S(gen[3096]),
			.SE(gen[3097]),

			.SELF(gen[3036]),
			.cell_state(gen[3036])
		); 

/******************* CELL 3037 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3037 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2976]),
			.N(gen[2977]),
			.NE(gen[2978]),

			.O(gen[3036]),
			.E(gen[3038]),

			.SO(gen[3096]),
			.S(gen[3097]),
			.SE(gen[3098]),

			.SELF(gen[3037]),
			.cell_state(gen[3037])
		); 

/******************* CELL 3038 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3038 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2977]),
			.N(gen[2978]),
			.NE(gen[2979]),

			.O(gen[3037]),
			.E(gen[3039]),

			.SO(gen[3097]),
			.S(gen[3098]),
			.SE(gen[3099]),

			.SELF(gen[3038]),
			.cell_state(gen[3038])
		); 

/******************* CELL 3039 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3039 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2978]),
			.N(gen[2979]),
			.NE(gen[2980]),

			.O(gen[3038]),
			.E(gen[3040]),

			.SO(gen[3098]),
			.S(gen[3099]),
			.SE(gen[3100]),

			.SELF(gen[3039]),
			.cell_state(gen[3039])
		); 

/******************* CELL 3040 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3040 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2979]),
			.N(gen[2980]),
			.NE(gen[2981]),

			.O(gen[3039]),
			.E(gen[3041]),

			.SO(gen[3099]),
			.S(gen[3100]),
			.SE(gen[3101]),

			.SELF(gen[3040]),
			.cell_state(gen[3040])
		); 

/******************* CELL 3041 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3041 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2980]),
			.N(gen[2981]),
			.NE(gen[2982]),

			.O(gen[3040]),
			.E(gen[3042]),

			.SO(gen[3100]),
			.S(gen[3101]),
			.SE(gen[3102]),

			.SELF(gen[3041]),
			.cell_state(gen[3041])
		); 

/******************* CELL 3042 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3042 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2981]),
			.N(gen[2982]),
			.NE(gen[2983]),

			.O(gen[3041]),
			.E(gen[3043]),

			.SO(gen[3101]),
			.S(gen[3102]),
			.SE(gen[3103]),

			.SELF(gen[3042]),
			.cell_state(gen[3042])
		); 

/******************* CELL 3043 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3043 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2982]),
			.N(gen[2983]),
			.NE(gen[2984]),

			.O(gen[3042]),
			.E(gen[3044]),

			.SO(gen[3102]),
			.S(gen[3103]),
			.SE(gen[3104]),

			.SELF(gen[3043]),
			.cell_state(gen[3043])
		); 

/******************* CELL 3044 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3044 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2983]),
			.N(gen[2984]),
			.NE(gen[2985]),

			.O(gen[3043]),
			.E(gen[3045]),

			.SO(gen[3103]),
			.S(gen[3104]),
			.SE(gen[3105]),

			.SELF(gen[3044]),
			.cell_state(gen[3044])
		); 

/******************* CELL 3045 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3045 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2984]),
			.N(gen[2985]),
			.NE(gen[2986]),

			.O(gen[3044]),
			.E(gen[3046]),

			.SO(gen[3104]),
			.S(gen[3105]),
			.SE(gen[3106]),

			.SELF(gen[3045]),
			.cell_state(gen[3045])
		); 

/******************* CELL 3046 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3046 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2985]),
			.N(gen[2986]),
			.NE(gen[2987]),

			.O(gen[3045]),
			.E(gen[3047]),

			.SO(gen[3105]),
			.S(gen[3106]),
			.SE(gen[3107]),

			.SELF(gen[3046]),
			.cell_state(gen[3046])
		); 

/******************* CELL 3047 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3047 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2986]),
			.N(gen[2987]),
			.NE(gen[2988]),

			.O(gen[3046]),
			.E(gen[3048]),

			.SO(gen[3106]),
			.S(gen[3107]),
			.SE(gen[3108]),

			.SELF(gen[3047]),
			.cell_state(gen[3047])
		); 

/******************* CELL 3048 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3048 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2987]),
			.N(gen[2988]),
			.NE(gen[2989]),

			.O(gen[3047]),
			.E(gen[3049]),

			.SO(gen[3107]),
			.S(gen[3108]),
			.SE(gen[3109]),

			.SELF(gen[3048]),
			.cell_state(gen[3048])
		); 

/******************* CELL 3049 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3049 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2988]),
			.N(gen[2989]),
			.NE(gen[2990]),

			.O(gen[3048]),
			.E(gen[3050]),

			.SO(gen[3108]),
			.S(gen[3109]),
			.SE(gen[3110]),

			.SELF(gen[3049]),
			.cell_state(gen[3049])
		); 

/******************* CELL 3050 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3050 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2989]),
			.N(gen[2990]),
			.NE(gen[2991]),

			.O(gen[3049]),
			.E(gen[3051]),

			.SO(gen[3109]),
			.S(gen[3110]),
			.SE(gen[3111]),

			.SELF(gen[3050]),
			.cell_state(gen[3050])
		); 

/******************* CELL 3051 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3051 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2990]),
			.N(gen[2991]),
			.NE(gen[2992]),

			.O(gen[3050]),
			.E(gen[3052]),

			.SO(gen[3110]),
			.S(gen[3111]),
			.SE(gen[3112]),

			.SELF(gen[3051]),
			.cell_state(gen[3051])
		); 

/******************* CELL 3052 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3052 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2991]),
			.N(gen[2992]),
			.NE(gen[2993]),

			.O(gen[3051]),
			.E(gen[3053]),

			.SO(gen[3111]),
			.S(gen[3112]),
			.SE(gen[3113]),

			.SELF(gen[3052]),
			.cell_state(gen[3052])
		); 

/******************* CELL 3053 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3053 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2992]),
			.N(gen[2993]),
			.NE(gen[2994]),

			.O(gen[3052]),
			.E(gen[3054]),

			.SO(gen[3112]),
			.S(gen[3113]),
			.SE(gen[3114]),

			.SELF(gen[3053]),
			.cell_state(gen[3053])
		); 

/******************* CELL 3054 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3054 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2993]),
			.N(gen[2994]),
			.NE(gen[2995]),

			.O(gen[3053]),
			.E(gen[3055]),

			.SO(gen[3113]),
			.S(gen[3114]),
			.SE(gen[3115]),

			.SELF(gen[3054]),
			.cell_state(gen[3054])
		); 

/******************* CELL 3055 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3055 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2994]),
			.N(gen[2995]),
			.NE(gen[2996]),

			.O(gen[3054]),
			.E(gen[3056]),

			.SO(gen[3114]),
			.S(gen[3115]),
			.SE(gen[3116]),

			.SELF(gen[3055]),
			.cell_state(gen[3055])
		); 

/******************* CELL 3056 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3056 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2995]),
			.N(gen[2996]),
			.NE(gen[2997]),

			.O(gen[3055]),
			.E(gen[3057]),

			.SO(gen[3115]),
			.S(gen[3116]),
			.SE(gen[3117]),

			.SELF(gen[3056]),
			.cell_state(gen[3056])
		); 

/******************* CELL 3057 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3057 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2996]),
			.N(gen[2997]),
			.NE(gen[2998]),

			.O(gen[3056]),
			.E(gen[3058]),

			.SO(gen[3116]),
			.S(gen[3117]),
			.SE(gen[3118]),

			.SELF(gen[3057]),
			.cell_state(gen[3057])
		); 

/******************* CELL 3058 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3058 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2997]),
			.N(gen[2998]),
			.NE(gen[2999]),

			.O(gen[3057]),
			.E(gen[3059]),

			.SO(gen[3117]),
			.S(gen[3118]),
			.SE(gen[3119]),

			.SELF(gen[3058]),
			.cell_state(gen[3058])
		); 

/******************* CELL 3059 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3059 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[2998]),
			.N(gen[2999]),
			.NE(gen[2998]),

			.O(gen[3058]),
			.E(gen[3058]),

			.SO(gen[3118]),
			.S(gen[3119]),
			.SE(gen[3118]),

			.SELF(gen[3059]),
			.cell_state(gen[3059])
		); 

/******************* CELL 3060 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3060 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3001]),
			.N(gen[3000]),
			.NE(gen[3001]),

			.O(gen[3061]),
			.E(gen[3061]),

			.SO(gen[3121]),
			.S(gen[3120]),
			.SE(gen[3121]),

			.SELF(gen[3060]),
			.cell_state(gen[3060])
		); 

/******************* CELL 3061 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3061 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3000]),
			.N(gen[3001]),
			.NE(gen[3002]),

			.O(gen[3060]),
			.E(gen[3062]),

			.SO(gen[3120]),
			.S(gen[3121]),
			.SE(gen[3122]),

			.SELF(gen[3061]),
			.cell_state(gen[3061])
		); 

/******************* CELL 3062 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3062 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3001]),
			.N(gen[3002]),
			.NE(gen[3003]),

			.O(gen[3061]),
			.E(gen[3063]),

			.SO(gen[3121]),
			.S(gen[3122]),
			.SE(gen[3123]),

			.SELF(gen[3062]),
			.cell_state(gen[3062])
		); 

/******************* CELL 3063 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3063 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3002]),
			.N(gen[3003]),
			.NE(gen[3004]),

			.O(gen[3062]),
			.E(gen[3064]),

			.SO(gen[3122]),
			.S(gen[3123]),
			.SE(gen[3124]),

			.SELF(gen[3063]),
			.cell_state(gen[3063])
		); 

/******************* CELL 3064 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3064 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3003]),
			.N(gen[3004]),
			.NE(gen[3005]),

			.O(gen[3063]),
			.E(gen[3065]),

			.SO(gen[3123]),
			.S(gen[3124]),
			.SE(gen[3125]),

			.SELF(gen[3064]),
			.cell_state(gen[3064])
		); 

/******************* CELL 3065 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3065 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3004]),
			.N(gen[3005]),
			.NE(gen[3006]),

			.O(gen[3064]),
			.E(gen[3066]),

			.SO(gen[3124]),
			.S(gen[3125]),
			.SE(gen[3126]),

			.SELF(gen[3065]),
			.cell_state(gen[3065])
		); 

/******************* CELL 3066 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3066 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3005]),
			.N(gen[3006]),
			.NE(gen[3007]),

			.O(gen[3065]),
			.E(gen[3067]),

			.SO(gen[3125]),
			.S(gen[3126]),
			.SE(gen[3127]),

			.SELF(gen[3066]),
			.cell_state(gen[3066])
		); 

/******************* CELL 3067 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3067 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3006]),
			.N(gen[3007]),
			.NE(gen[3008]),

			.O(gen[3066]),
			.E(gen[3068]),

			.SO(gen[3126]),
			.S(gen[3127]),
			.SE(gen[3128]),

			.SELF(gen[3067]),
			.cell_state(gen[3067])
		); 

/******************* CELL 3068 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3068 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3007]),
			.N(gen[3008]),
			.NE(gen[3009]),

			.O(gen[3067]),
			.E(gen[3069]),

			.SO(gen[3127]),
			.S(gen[3128]),
			.SE(gen[3129]),

			.SELF(gen[3068]),
			.cell_state(gen[3068])
		); 

/******************* CELL 3069 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3069 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3008]),
			.N(gen[3009]),
			.NE(gen[3010]),

			.O(gen[3068]),
			.E(gen[3070]),

			.SO(gen[3128]),
			.S(gen[3129]),
			.SE(gen[3130]),

			.SELF(gen[3069]),
			.cell_state(gen[3069])
		); 

/******************* CELL 3070 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3070 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3009]),
			.N(gen[3010]),
			.NE(gen[3011]),

			.O(gen[3069]),
			.E(gen[3071]),

			.SO(gen[3129]),
			.S(gen[3130]),
			.SE(gen[3131]),

			.SELF(gen[3070]),
			.cell_state(gen[3070])
		); 

/******************* CELL 3071 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3071 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3010]),
			.N(gen[3011]),
			.NE(gen[3012]),

			.O(gen[3070]),
			.E(gen[3072]),

			.SO(gen[3130]),
			.S(gen[3131]),
			.SE(gen[3132]),

			.SELF(gen[3071]),
			.cell_state(gen[3071])
		); 

/******************* CELL 3072 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3072 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3011]),
			.N(gen[3012]),
			.NE(gen[3013]),

			.O(gen[3071]),
			.E(gen[3073]),

			.SO(gen[3131]),
			.S(gen[3132]),
			.SE(gen[3133]),

			.SELF(gen[3072]),
			.cell_state(gen[3072])
		); 

/******************* CELL 3073 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3073 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3012]),
			.N(gen[3013]),
			.NE(gen[3014]),

			.O(gen[3072]),
			.E(gen[3074]),

			.SO(gen[3132]),
			.S(gen[3133]),
			.SE(gen[3134]),

			.SELF(gen[3073]),
			.cell_state(gen[3073])
		); 

/******************* CELL 3074 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3074 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3013]),
			.N(gen[3014]),
			.NE(gen[3015]),

			.O(gen[3073]),
			.E(gen[3075]),

			.SO(gen[3133]),
			.S(gen[3134]),
			.SE(gen[3135]),

			.SELF(gen[3074]),
			.cell_state(gen[3074])
		); 

/******************* CELL 3075 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3075 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3014]),
			.N(gen[3015]),
			.NE(gen[3016]),

			.O(gen[3074]),
			.E(gen[3076]),

			.SO(gen[3134]),
			.S(gen[3135]),
			.SE(gen[3136]),

			.SELF(gen[3075]),
			.cell_state(gen[3075])
		); 

/******************* CELL 3076 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3076 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3015]),
			.N(gen[3016]),
			.NE(gen[3017]),

			.O(gen[3075]),
			.E(gen[3077]),

			.SO(gen[3135]),
			.S(gen[3136]),
			.SE(gen[3137]),

			.SELF(gen[3076]),
			.cell_state(gen[3076])
		); 

/******************* CELL 3077 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3077 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3016]),
			.N(gen[3017]),
			.NE(gen[3018]),

			.O(gen[3076]),
			.E(gen[3078]),

			.SO(gen[3136]),
			.S(gen[3137]),
			.SE(gen[3138]),

			.SELF(gen[3077]),
			.cell_state(gen[3077])
		); 

/******************* CELL 3078 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3078 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3017]),
			.N(gen[3018]),
			.NE(gen[3019]),

			.O(gen[3077]),
			.E(gen[3079]),

			.SO(gen[3137]),
			.S(gen[3138]),
			.SE(gen[3139]),

			.SELF(gen[3078]),
			.cell_state(gen[3078])
		); 

/******************* CELL 3079 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3079 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3018]),
			.N(gen[3019]),
			.NE(gen[3020]),

			.O(gen[3078]),
			.E(gen[3080]),

			.SO(gen[3138]),
			.S(gen[3139]),
			.SE(gen[3140]),

			.SELF(gen[3079]),
			.cell_state(gen[3079])
		); 

/******************* CELL 3080 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3080 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3019]),
			.N(gen[3020]),
			.NE(gen[3021]),

			.O(gen[3079]),
			.E(gen[3081]),

			.SO(gen[3139]),
			.S(gen[3140]),
			.SE(gen[3141]),

			.SELF(gen[3080]),
			.cell_state(gen[3080])
		); 

/******************* CELL 3081 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3081 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3020]),
			.N(gen[3021]),
			.NE(gen[3022]),

			.O(gen[3080]),
			.E(gen[3082]),

			.SO(gen[3140]),
			.S(gen[3141]),
			.SE(gen[3142]),

			.SELF(gen[3081]),
			.cell_state(gen[3081])
		); 

/******************* CELL 3082 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3082 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3021]),
			.N(gen[3022]),
			.NE(gen[3023]),

			.O(gen[3081]),
			.E(gen[3083]),

			.SO(gen[3141]),
			.S(gen[3142]),
			.SE(gen[3143]),

			.SELF(gen[3082]),
			.cell_state(gen[3082])
		); 

/******************* CELL 3083 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3083 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3022]),
			.N(gen[3023]),
			.NE(gen[3024]),

			.O(gen[3082]),
			.E(gen[3084]),

			.SO(gen[3142]),
			.S(gen[3143]),
			.SE(gen[3144]),

			.SELF(gen[3083]),
			.cell_state(gen[3083])
		); 

/******************* CELL 3084 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3084 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3023]),
			.N(gen[3024]),
			.NE(gen[3025]),

			.O(gen[3083]),
			.E(gen[3085]),

			.SO(gen[3143]),
			.S(gen[3144]),
			.SE(gen[3145]),

			.SELF(gen[3084]),
			.cell_state(gen[3084])
		); 

/******************* CELL 3085 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3085 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3024]),
			.N(gen[3025]),
			.NE(gen[3026]),

			.O(gen[3084]),
			.E(gen[3086]),

			.SO(gen[3144]),
			.S(gen[3145]),
			.SE(gen[3146]),

			.SELF(gen[3085]),
			.cell_state(gen[3085])
		); 

/******************* CELL 3086 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3086 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3025]),
			.N(gen[3026]),
			.NE(gen[3027]),

			.O(gen[3085]),
			.E(gen[3087]),

			.SO(gen[3145]),
			.S(gen[3146]),
			.SE(gen[3147]),

			.SELF(gen[3086]),
			.cell_state(gen[3086])
		); 

/******************* CELL 3087 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3087 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3026]),
			.N(gen[3027]),
			.NE(gen[3028]),

			.O(gen[3086]),
			.E(gen[3088]),

			.SO(gen[3146]),
			.S(gen[3147]),
			.SE(gen[3148]),

			.SELF(gen[3087]),
			.cell_state(gen[3087])
		); 

/******************* CELL 3088 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3088 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3027]),
			.N(gen[3028]),
			.NE(gen[3029]),

			.O(gen[3087]),
			.E(gen[3089]),

			.SO(gen[3147]),
			.S(gen[3148]),
			.SE(gen[3149]),

			.SELF(gen[3088]),
			.cell_state(gen[3088])
		); 

/******************* CELL 3089 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3089 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3028]),
			.N(gen[3029]),
			.NE(gen[3030]),

			.O(gen[3088]),
			.E(gen[3090]),

			.SO(gen[3148]),
			.S(gen[3149]),
			.SE(gen[3150]),

			.SELF(gen[3089]),
			.cell_state(gen[3089])
		); 

/******************* CELL 3090 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3090 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3029]),
			.N(gen[3030]),
			.NE(gen[3031]),

			.O(gen[3089]),
			.E(gen[3091]),

			.SO(gen[3149]),
			.S(gen[3150]),
			.SE(gen[3151]),

			.SELF(gen[3090]),
			.cell_state(gen[3090])
		); 

/******************* CELL 3091 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3091 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3030]),
			.N(gen[3031]),
			.NE(gen[3032]),

			.O(gen[3090]),
			.E(gen[3092]),

			.SO(gen[3150]),
			.S(gen[3151]),
			.SE(gen[3152]),

			.SELF(gen[3091]),
			.cell_state(gen[3091])
		); 

/******************* CELL 3092 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3092 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3031]),
			.N(gen[3032]),
			.NE(gen[3033]),

			.O(gen[3091]),
			.E(gen[3093]),

			.SO(gen[3151]),
			.S(gen[3152]),
			.SE(gen[3153]),

			.SELF(gen[3092]),
			.cell_state(gen[3092])
		); 

/******************* CELL 3093 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3093 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3032]),
			.N(gen[3033]),
			.NE(gen[3034]),

			.O(gen[3092]),
			.E(gen[3094]),

			.SO(gen[3152]),
			.S(gen[3153]),
			.SE(gen[3154]),

			.SELF(gen[3093]),
			.cell_state(gen[3093])
		); 

/******************* CELL 3094 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3094 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3033]),
			.N(gen[3034]),
			.NE(gen[3035]),

			.O(gen[3093]),
			.E(gen[3095]),

			.SO(gen[3153]),
			.S(gen[3154]),
			.SE(gen[3155]),

			.SELF(gen[3094]),
			.cell_state(gen[3094])
		); 

/******************* CELL 3095 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3095 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3034]),
			.N(gen[3035]),
			.NE(gen[3036]),

			.O(gen[3094]),
			.E(gen[3096]),

			.SO(gen[3154]),
			.S(gen[3155]),
			.SE(gen[3156]),

			.SELF(gen[3095]),
			.cell_state(gen[3095])
		); 

/******************* CELL 3096 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3096 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3035]),
			.N(gen[3036]),
			.NE(gen[3037]),

			.O(gen[3095]),
			.E(gen[3097]),

			.SO(gen[3155]),
			.S(gen[3156]),
			.SE(gen[3157]),

			.SELF(gen[3096]),
			.cell_state(gen[3096])
		); 

/******************* CELL 3097 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3097 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3036]),
			.N(gen[3037]),
			.NE(gen[3038]),

			.O(gen[3096]),
			.E(gen[3098]),

			.SO(gen[3156]),
			.S(gen[3157]),
			.SE(gen[3158]),

			.SELF(gen[3097]),
			.cell_state(gen[3097])
		); 

/******************* CELL 3098 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3098 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3037]),
			.N(gen[3038]),
			.NE(gen[3039]),

			.O(gen[3097]),
			.E(gen[3099]),

			.SO(gen[3157]),
			.S(gen[3158]),
			.SE(gen[3159]),

			.SELF(gen[3098]),
			.cell_state(gen[3098])
		); 

/******************* CELL 3099 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3099 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3038]),
			.N(gen[3039]),
			.NE(gen[3040]),

			.O(gen[3098]),
			.E(gen[3100]),

			.SO(gen[3158]),
			.S(gen[3159]),
			.SE(gen[3160]),

			.SELF(gen[3099]),
			.cell_state(gen[3099])
		); 

/******************* CELL 3100 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3100 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3039]),
			.N(gen[3040]),
			.NE(gen[3041]),

			.O(gen[3099]),
			.E(gen[3101]),

			.SO(gen[3159]),
			.S(gen[3160]),
			.SE(gen[3161]),

			.SELF(gen[3100]),
			.cell_state(gen[3100])
		); 

/******************* CELL 3101 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3101 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3040]),
			.N(gen[3041]),
			.NE(gen[3042]),

			.O(gen[3100]),
			.E(gen[3102]),

			.SO(gen[3160]),
			.S(gen[3161]),
			.SE(gen[3162]),

			.SELF(gen[3101]),
			.cell_state(gen[3101])
		); 

/******************* CELL 3102 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3102 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3041]),
			.N(gen[3042]),
			.NE(gen[3043]),

			.O(gen[3101]),
			.E(gen[3103]),

			.SO(gen[3161]),
			.S(gen[3162]),
			.SE(gen[3163]),

			.SELF(gen[3102]),
			.cell_state(gen[3102])
		); 

/******************* CELL 3103 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3103 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3042]),
			.N(gen[3043]),
			.NE(gen[3044]),

			.O(gen[3102]),
			.E(gen[3104]),

			.SO(gen[3162]),
			.S(gen[3163]),
			.SE(gen[3164]),

			.SELF(gen[3103]),
			.cell_state(gen[3103])
		); 

/******************* CELL 3104 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3104 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3043]),
			.N(gen[3044]),
			.NE(gen[3045]),

			.O(gen[3103]),
			.E(gen[3105]),

			.SO(gen[3163]),
			.S(gen[3164]),
			.SE(gen[3165]),

			.SELF(gen[3104]),
			.cell_state(gen[3104])
		); 

/******************* CELL 3105 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3105 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3044]),
			.N(gen[3045]),
			.NE(gen[3046]),

			.O(gen[3104]),
			.E(gen[3106]),

			.SO(gen[3164]),
			.S(gen[3165]),
			.SE(gen[3166]),

			.SELF(gen[3105]),
			.cell_state(gen[3105])
		); 

/******************* CELL 3106 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3106 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3045]),
			.N(gen[3046]),
			.NE(gen[3047]),

			.O(gen[3105]),
			.E(gen[3107]),

			.SO(gen[3165]),
			.S(gen[3166]),
			.SE(gen[3167]),

			.SELF(gen[3106]),
			.cell_state(gen[3106])
		); 

/******************* CELL 3107 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3107 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3046]),
			.N(gen[3047]),
			.NE(gen[3048]),

			.O(gen[3106]),
			.E(gen[3108]),

			.SO(gen[3166]),
			.S(gen[3167]),
			.SE(gen[3168]),

			.SELF(gen[3107]),
			.cell_state(gen[3107])
		); 

/******************* CELL 3108 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3108 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3047]),
			.N(gen[3048]),
			.NE(gen[3049]),

			.O(gen[3107]),
			.E(gen[3109]),

			.SO(gen[3167]),
			.S(gen[3168]),
			.SE(gen[3169]),

			.SELF(gen[3108]),
			.cell_state(gen[3108])
		); 

/******************* CELL 3109 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3109 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3048]),
			.N(gen[3049]),
			.NE(gen[3050]),

			.O(gen[3108]),
			.E(gen[3110]),

			.SO(gen[3168]),
			.S(gen[3169]),
			.SE(gen[3170]),

			.SELF(gen[3109]),
			.cell_state(gen[3109])
		); 

/******************* CELL 3110 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3110 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3049]),
			.N(gen[3050]),
			.NE(gen[3051]),

			.O(gen[3109]),
			.E(gen[3111]),

			.SO(gen[3169]),
			.S(gen[3170]),
			.SE(gen[3171]),

			.SELF(gen[3110]),
			.cell_state(gen[3110])
		); 

/******************* CELL 3111 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3111 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3050]),
			.N(gen[3051]),
			.NE(gen[3052]),

			.O(gen[3110]),
			.E(gen[3112]),

			.SO(gen[3170]),
			.S(gen[3171]),
			.SE(gen[3172]),

			.SELF(gen[3111]),
			.cell_state(gen[3111])
		); 

/******************* CELL 3112 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3112 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3051]),
			.N(gen[3052]),
			.NE(gen[3053]),

			.O(gen[3111]),
			.E(gen[3113]),

			.SO(gen[3171]),
			.S(gen[3172]),
			.SE(gen[3173]),

			.SELF(gen[3112]),
			.cell_state(gen[3112])
		); 

/******************* CELL 3113 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3113 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3052]),
			.N(gen[3053]),
			.NE(gen[3054]),

			.O(gen[3112]),
			.E(gen[3114]),

			.SO(gen[3172]),
			.S(gen[3173]),
			.SE(gen[3174]),

			.SELF(gen[3113]),
			.cell_state(gen[3113])
		); 

/******************* CELL 3114 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3114 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3053]),
			.N(gen[3054]),
			.NE(gen[3055]),

			.O(gen[3113]),
			.E(gen[3115]),

			.SO(gen[3173]),
			.S(gen[3174]),
			.SE(gen[3175]),

			.SELF(gen[3114]),
			.cell_state(gen[3114])
		); 

/******************* CELL 3115 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3115 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3054]),
			.N(gen[3055]),
			.NE(gen[3056]),

			.O(gen[3114]),
			.E(gen[3116]),

			.SO(gen[3174]),
			.S(gen[3175]),
			.SE(gen[3176]),

			.SELF(gen[3115]),
			.cell_state(gen[3115])
		); 

/******************* CELL 3116 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3116 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3055]),
			.N(gen[3056]),
			.NE(gen[3057]),

			.O(gen[3115]),
			.E(gen[3117]),

			.SO(gen[3175]),
			.S(gen[3176]),
			.SE(gen[3177]),

			.SELF(gen[3116]),
			.cell_state(gen[3116])
		); 

/******************* CELL 3117 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3117 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3056]),
			.N(gen[3057]),
			.NE(gen[3058]),

			.O(gen[3116]),
			.E(gen[3118]),

			.SO(gen[3176]),
			.S(gen[3177]),
			.SE(gen[3178]),

			.SELF(gen[3117]),
			.cell_state(gen[3117])
		); 

/******************* CELL 3118 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3118 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3057]),
			.N(gen[3058]),
			.NE(gen[3059]),

			.O(gen[3117]),
			.E(gen[3119]),

			.SO(gen[3177]),
			.S(gen[3178]),
			.SE(gen[3179]),

			.SELF(gen[3118]),
			.cell_state(gen[3118])
		); 

/******************* CELL 3119 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3119 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3058]),
			.N(gen[3059]),
			.NE(gen[3058]),

			.O(gen[3118]),
			.E(gen[3118]),

			.SO(gen[3178]),
			.S(gen[3179]),
			.SE(gen[3178]),

			.SELF(gen[3119]),
			.cell_state(gen[3119])
		); 

/******************* CELL 3120 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3120 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3061]),
			.N(gen[3060]),
			.NE(gen[3061]),

			.O(gen[3121]),
			.E(gen[3121]),

			.SO(gen[3181]),
			.S(gen[3180]),
			.SE(gen[3181]),

			.SELF(gen[3120]),
			.cell_state(gen[3120])
		); 

/******************* CELL 3121 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3121 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3060]),
			.N(gen[3061]),
			.NE(gen[3062]),

			.O(gen[3120]),
			.E(gen[3122]),

			.SO(gen[3180]),
			.S(gen[3181]),
			.SE(gen[3182]),

			.SELF(gen[3121]),
			.cell_state(gen[3121])
		); 

/******************* CELL 3122 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3122 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3061]),
			.N(gen[3062]),
			.NE(gen[3063]),

			.O(gen[3121]),
			.E(gen[3123]),

			.SO(gen[3181]),
			.S(gen[3182]),
			.SE(gen[3183]),

			.SELF(gen[3122]),
			.cell_state(gen[3122])
		); 

/******************* CELL 3123 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3123 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3062]),
			.N(gen[3063]),
			.NE(gen[3064]),

			.O(gen[3122]),
			.E(gen[3124]),

			.SO(gen[3182]),
			.S(gen[3183]),
			.SE(gen[3184]),

			.SELF(gen[3123]),
			.cell_state(gen[3123])
		); 

/******************* CELL 3124 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3124 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3063]),
			.N(gen[3064]),
			.NE(gen[3065]),

			.O(gen[3123]),
			.E(gen[3125]),

			.SO(gen[3183]),
			.S(gen[3184]),
			.SE(gen[3185]),

			.SELF(gen[3124]),
			.cell_state(gen[3124])
		); 

/******************* CELL 3125 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3125 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3064]),
			.N(gen[3065]),
			.NE(gen[3066]),

			.O(gen[3124]),
			.E(gen[3126]),

			.SO(gen[3184]),
			.S(gen[3185]),
			.SE(gen[3186]),

			.SELF(gen[3125]),
			.cell_state(gen[3125])
		); 

/******************* CELL 3126 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3126 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3065]),
			.N(gen[3066]),
			.NE(gen[3067]),

			.O(gen[3125]),
			.E(gen[3127]),

			.SO(gen[3185]),
			.S(gen[3186]),
			.SE(gen[3187]),

			.SELF(gen[3126]),
			.cell_state(gen[3126])
		); 

/******************* CELL 3127 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3127 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3066]),
			.N(gen[3067]),
			.NE(gen[3068]),

			.O(gen[3126]),
			.E(gen[3128]),

			.SO(gen[3186]),
			.S(gen[3187]),
			.SE(gen[3188]),

			.SELF(gen[3127]),
			.cell_state(gen[3127])
		); 

/******************* CELL 3128 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3128 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3067]),
			.N(gen[3068]),
			.NE(gen[3069]),

			.O(gen[3127]),
			.E(gen[3129]),

			.SO(gen[3187]),
			.S(gen[3188]),
			.SE(gen[3189]),

			.SELF(gen[3128]),
			.cell_state(gen[3128])
		); 

/******************* CELL 3129 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3129 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3068]),
			.N(gen[3069]),
			.NE(gen[3070]),

			.O(gen[3128]),
			.E(gen[3130]),

			.SO(gen[3188]),
			.S(gen[3189]),
			.SE(gen[3190]),

			.SELF(gen[3129]),
			.cell_state(gen[3129])
		); 

/******************* CELL 3130 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3130 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3069]),
			.N(gen[3070]),
			.NE(gen[3071]),

			.O(gen[3129]),
			.E(gen[3131]),

			.SO(gen[3189]),
			.S(gen[3190]),
			.SE(gen[3191]),

			.SELF(gen[3130]),
			.cell_state(gen[3130])
		); 

/******************* CELL 3131 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3131 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3070]),
			.N(gen[3071]),
			.NE(gen[3072]),

			.O(gen[3130]),
			.E(gen[3132]),

			.SO(gen[3190]),
			.S(gen[3191]),
			.SE(gen[3192]),

			.SELF(gen[3131]),
			.cell_state(gen[3131])
		); 

/******************* CELL 3132 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3132 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3071]),
			.N(gen[3072]),
			.NE(gen[3073]),

			.O(gen[3131]),
			.E(gen[3133]),

			.SO(gen[3191]),
			.S(gen[3192]),
			.SE(gen[3193]),

			.SELF(gen[3132]),
			.cell_state(gen[3132])
		); 

/******************* CELL 3133 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3133 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3072]),
			.N(gen[3073]),
			.NE(gen[3074]),

			.O(gen[3132]),
			.E(gen[3134]),

			.SO(gen[3192]),
			.S(gen[3193]),
			.SE(gen[3194]),

			.SELF(gen[3133]),
			.cell_state(gen[3133])
		); 

/******************* CELL 3134 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3134 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3073]),
			.N(gen[3074]),
			.NE(gen[3075]),

			.O(gen[3133]),
			.E(gen[3135]),

			.SO(gen[3193]),
			.S(gen[3194]),
			.SE(gen[3195]),

			.SELF(gen[3134]),
			.cell_state(gen[3134])
		); 

/******************* CELL 3135 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3135 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3074]),
			.N(gen[3075]),
			.NE(gen[3076]),

			.O(gen[3134]),
			.E(gen[3136]),

			.SO(gen[3194]),
			.S(gen[3195]),
			.SE(gen[3196]),

			.SELF(gen[3135]),
			.cell_state(gen[3135])
		); 

/******************* CELL 3136 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3136 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3075]),
			.N(gen[3076]),
			.NE(gen[3077]),

			.O(gen[3135]),
			.E(gen[3137]),

			.SO(gen[3195]),
			.S(gen[3196]),
			.SE(gen[3197]),

			.SELF(gen[3136]),
			.cell_state(gen[3136])
		); 

/******************* CELL 3137 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3137 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3076]),
			.N(gen[3077]),
			.NE(gen[3078]),

			.O(gen[3136]),
			.E(gen[3138]),

			.SO(gen[3196]),
			.S(gen[3197]),
			.SE(gen[3198]),

			.SELF(gen[3137]),
			.cell_state(gen[3137])
		); 

/******************* CELL 3138 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3138 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3077]),
			.N(gen[3078]),
			.NE(gen[3079]),

			.O(gen[3137]),
			.E(gen[3139]),

			.SO(gen[3197]),
			.S(gen[3198]),
			.SE(gen[3199]),

			.SELF(gen[3138]),
			.cell_state(gen[3138])
		); 

/******************* CELL 3139 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3139 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3078]),
			.N(gen[3079]),
			.NE(gen[3080]),

			.O(gen[3138]),
			.E(gen[3140]),

			.SO(gen[3198]),
			.S(gen[3199]),
			.SE(gen[3200]),

			.SELF(gen[3139]),
			.cell_state(gen[3139])
		); 

/******************* CELL 3140 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3140 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3079]),
			.N(gen[3080]),
			.NE(gen[3081]),

			.O(gen[3139]),
			.E(gen[3141]),

			.SO(gen[3199]),
			.S(gen[3200]),
			.SE(gen[3201]),

			.SELF(gen[3140]),
			.cell_state(gen[3140])
		); 

/******************* CELL 3141 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3141 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3080]),
			.N(gen[3081]),
			.NE(gen[3082]),

			.O(gen[3140]),
			.E(gen[3142]),

			.SO(gen[3200]),
			.S(gen[3201]),
			.SE(gen[3202]),

			.SELF(gen[3141]),
			.cell_state(gen[3141])
		); 

/******************* CELL 3142 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3142 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3081]),
			.N(gen[3082]),
			.NE(gen[3083]),

			.O(gen[3141]),
			.E(gen[3143]),

			.SO(gen[3201]),
			.S(gen[3202]),
			.SE(gen[3203]),

			.SELF(gen[3142]),
			.cell_state(gen[3142])
		); 

/******************* CELL 3143 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3143 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3082]),
			.N(gen[3083]),
			.NE(gen[3084]),

			.O(gen[3142]),
			.E(gen[3144]),

			.SO(gen[3202]),
			.S(gen[3203]),
			.SE(gen[3204]),

			.SELF(gen[3143]),
			.cell_state(gen[3143])
		); 

/******************* CELL 3144 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3144 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3083]),
			.N(gen[3084]),
			.NE(gen[3085]),

			.O(gen[3143]),
			.E(gen[3145]),

			.SO(gen[3203]),
			.S(gen[3204]),
			.SE(gen[3205]),

			.SELF(gen[3144]),
			.cell_state(gen[3144])
		); 

/******************* CELL 3145 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3145 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3084]),
			.N(gen[3085]),
			.NE(gen[3086]),

			.O(gen[3144]),
			.E(gen[3146]),

			.SO(gen[3204]),
			.S(gen[3205]),
			.SE(gen[3206]),

			.SELF(gen[3145]),
			.cell_state(gen[3145])
		); 

/******************* CELL 3146 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3146 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3085]),
			.N(gen[3086]),
			.NE(gen[3087]),

			.O(gen[3145]),
			.E(gen[3147]),

			.SO(gen[3205]),
			.S(gen[3206]),
			.SE(gen[3207]),

			.SELF(gen[3146]),
			.cell_state(gen[3146])
		); 

/******************* CELL 3147 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3147 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3086]),
			.N(gen[3087]),
			.NE(gen[3088]),

			.O(gen[3146]),
			.E(gen[3148]),

			.SO(gen[3206]),
			.S(gen[3207]),
			.SE(gen[3208]),

			.SELF(gen[3147]),
			.cell_state(gen[3147])
		); 

/******************* CELL 3148 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3148 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3087]),
			.N(gen[3088]),
			.NE(gen[3089]),

			.O(gen[3147]),
			.E(gen[3149]),

			.SO(gen[3207]),
			.S(gen[3208]),
			.SE(gen[3209]),

			.SELF(gen[3148]),
			.cell_state(gen[3148])
		); 

/******************* CELL 3149 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3149 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3088]),
			.N(gen[3089]),
			.NE(gen[3090]),

			.O(gen[3148]),
			.E(gen[3150]),

			.SO(gen[3208]),
			.S(gen[3209]),
			.SE(gen[3210]),

			.SELF(gen[3149]),
			.cell_state(gen[3149])
		); 

/******************* CELL 3150 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3150 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3089]),
			.N(gen[3090]),
			.NE(gen[3091]),

			.O(gen[3149]),
			.E(gen[3151]),

			.SO(gen[3209]),
			.S(gen[3210]),
			.SE(gen[3211]),

			.SELF(gen[3150]),
			.cell_state(gen[3150])
		); 

/******************* CELL 3151 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3151 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3090]),
			.N(gen[3091]),
			.NE(gen[3092]),

			.O(gen[3150]),
			.E(gen[3152]),

			.SO(gen[3210]),
			.S(gen[3211]),
			.SE(gen[3212]),

			.SELF(gen[3151]),
			.cell_state(gen[3151])
		); 

/******************* CELL 3152 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3152 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3091]),
			.N(gen[3092]),
			.NE(gen[3093]),

			.O(gen[3151]),
			.E(gen[3153]),

			.SO(gen[3211]),
			.S(gen[3212]),
			.SE(gen[3213]),

			.SELF(gen[3152]),
			.cell_state(gen[3152])
		); 

/******************* CELL 3153 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3153 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3092]),
			.N(gen[3093]),
			.NE(gen[3094]),

			.O(gen[3152]),
			.E(gen[3154]),

			.SO(gen[3212]),
			.S(gen[3213]),
			.SE(gen[3214]),

			.SELF(gen[3153]),
			.cell_state(gen[3153])
		); 

/******************* CELL 3154 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3154 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3093]),
			.N(gen[3094]),
			.NE(gen[3095]),

			.O(gen[3153]),
			.E(gen[3155]),

			.SO(gen[3213]),
			.S(gen[3214]),
			.SE(gen[3215]),

			.SELF(gen[3154]),
			.cell_state(gen[3154])
		); 

/******************* CELL 3155 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3155 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3094]),
			.N(gen[3095]),
			.NE(gen[3096]),

			.O(gen[3154]),
			.E(gen[3156]),

			.SO(gen[3214]),
			.S(gen[3215]),
			.SE(gen[3216]),

			.SELF(gen[3155]),
			.cell_state(gen[3155])
		); 

/******************* CELL 3156 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3156 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3095]),
			.N(gen[3096]),
			.NE(gen[3097]),

			.O(gen[3155]),
			.E(gen[3157]),

			.SO(gen[3215]),
			.S(gen[3216]),
			.SE(gen[3217]),

			.SELF(gen[3156]),
			.cell_state(gen[3156])
		); 

/******************* CELL 3157 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3157 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3096]),
			.N(gen[3097]),
			.NE(gen[3098]),

			.O(gen[3156]),
			.E(gen[3158]),

			.SO(gen[3216]),
			.S(gen[3217]),
			.SE(gen[3218]),

			.SELF(gen[3157]),
			.cell_state(gen[3157])
		); 

/******************* CELL 3158 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3158 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3097]),
			.N(gen[3098]),
			.NE(gen[3099]),

			.O(gen[3157]),
			.E(gen[3159]),

			.SO(gen[3217]),
			.S(gen[3218]),
			.SE(gen[3219]),

			.SELF(gen[3158]),
			.cell_state(gen[3158])
		); 

/******************* CELL 3159 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3159 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3098]),
			.N(gen[3099]),
			.NE(gen[3100]),

			.O(gen[3158]),
			.E(gen[3160]),

			.SO(gen[3218]),
			.S(gen[3219]),
			.SE(gen[3220]),

			.SELF(gen[3159]),
			.cell_state(gen[3159])
		); 

/******************* CELL 3160 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3160 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3099]),
			.N(gen[3100]),
			.NE(gen[3101]),

			.O(gen[3159]),
			.E(gen[3161]),

			.SO(gen[3219]),
			.S(gen[3220]),
			.SE(gen[3221]),

			.SELF(gen[3160]),
			.cell_state(gen[3160])
		); 

/******************* CELL 3161 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3161 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3100]),
			.N(gen[3101]),
			.NE(gen[3102]),

			.O(gen[3160]),
			.E(gen[3162]),

			.SO(gen[3220]),
			.S(gen[3221]),
			.SE(gen[3222]),

			.SELF(gen[3161]),
			.cell_state(gen[3161])
		); 

/******************* CELL 3162 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3162 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3101]),
			.N(gen[3102]),
			.NE(gen[3103]),

			.O(gen[3161]),
			.E(gen[3163]),

			.SO(gen[3221]),
			.S(gen[3222]),
			.SE(gen[3223]),

			.SELF(gen[3162]),
			.cell_state(gen[3162])
		); 

/******************* CELL 3163 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3163 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3102]),
			.N(gen[3103]),
			.NE(gen[3104]),

			.O(gen[3162]),
			.E(gen[3164]),

			.SO(gen[3222]),
			.S(gen[3223]),
			.SE(gen[3224]),

			.SELF(gen[3163]),
			.cell_state(gen[3163])
		); 

/******************* CELL 3164 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3164 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3103]),
			.N(gen[3104]),
			.NE(gen[3105]),

			.O(gen[3163]),
			.E(gen[3165]),

			.SO(gen[3223]),
			.S(gen[3224]),
			.SE(gen[3225]),

			.SELF(gen[3164]),
			.cell_state(gen[3164])
		); 

/******************* CELL 3165 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3165 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3104]),
			.N(gen[3105]),
			.NE(gen[3106]),

			.O(gen[3164]),
			.E(gen[3166]),

			.SO(gen[3224]),
			.S(gen[3225]),
			.SE(gen[3226]),

			.SELF(gen[3165]),
			.cell_state(gen[3165])
		); 

/******************* CELL 3166 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3166 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3105]),
			.N(gen[3106]),
			.NE(gen[3107]),

			.O(gen[3165]),
			.E(gen[3167]),

			.SO(gen[3225]),
			.S(gen[3226]),
			.SE(gen[3227]),

			.SELF(gen[3166]),
			.cell_state(gen[3166])
		); 

/******************* CELL 3167 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3167 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3106]),
			.N(gen[3107]),
			.NE(gen[3108]),

			.O(gen[3166]),
			.E(gen[3168]),

			.SO(gen[3226]),
			.S(gen[3227]),
			.SE(gen[3228]),

			.SELF(gen[3167]),
			.cell_state(gen[3167])
		); 

/******************* CELL 3168 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3168 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3107]),
			.N(gen[3108]),
			.NE(gen[3109]),

			.O(gen[3167]),
			.E(gen[3169]),

			.SO(gen[3227]),
			.S(gen[3228]),
			.SE(gen[3229]),

			.SELF(gen[3168]),
			.cell_state(gen[3168])
		); 

/******************* CELL 3169 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3169 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3108]),
			.N(gen[3109]),
			.NE(gen[3110]),

			.O(gen[3168]),
			.E(gen[3170]),

			.SO(gen[3228]),
			.S(gen[3229]),
			.SE(gen[3230]),

			.SELF(gen[3169]),
			.cell_state(gen[3169])
		); 

/******************* CELL 3170 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3170 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3109]),
			.N(gen[3110]),
			.NE(gen[3111]),

			.O(gen[3169]),
			.E(gen[3171]),

			.SO(gen[3229]),
			.S(gen[3230]),
			.SE(gen[3231]),

			.SELF(gen[3170]),
			.cell_state(gen[3170])
		); 

/******************* CELL 3171 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3171 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3110]),
			.N(gen[3111]),
			.NE(gen[3112]),

			.O(gen[3170]),
			.E(gen[3172]),

			.SO(gen[3230]),
			.S(gen[3231]),
			.SE(gen[3232]),

			.SELF(gen[3171]),
			.cell_state(gen[3171])
		); 

/******************* CELL 3172 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3172 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3111]),
			.N(gen[3112]),
			.NE(gen[3113]),

			.O(gen[3171]),
			.E(gen[3173]),

			.SO(gen[3231]),
			.S(gen[3232]),
			.SE(gen[3233]),

			.SELF(gen[3172]),
			.cell_state(gen[3172])
		); 

/******************* CELL 3173 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3173 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3112]),
			.N(gen[3113]),
			.NE(gen[3114]),

			.O(gen[3172]),
			.E(gen[3174]),

			.SO(gen[3232]),
			.S(gen[3233]),
			.SE(gen[3234]),

			.SELF(gen[3173]),
			.cell_state(gen[3173])
		); 

/******************* CELL 3174 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3174 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3113]),
			.N(gen[3114]),
			.NE(gen[3115]),

			.O(gen[3173]),
			.E(gen[3175]),

			.SO(gen[3233]),
			.S(gen[3234]),
			.SE(gen[3235]),

			.SELF(gen[3174]),
			.cell_state(gen[3174])
		); 

/******************* CELL 3175 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3175 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3114]),
			.N(gen[3115]),
			.NE(gen[3116]),

			.O(gen[3174]),
			.E(gen[3176]),

			.SO(gen[3234]),
			.S(gen[3235]),
			.SE(gen[3236]),

			.SELF(gen[3175]),
			.cell_state(gen[3175])
		); 

/******************* CELL 3176 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3176 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3115]),
			.N(gen[3116]),
			.NE(gen[3117]),

			.O(gen[3175]),
			.E(gen[3177]),

			.SO(gen[3235]),
			.S(gen[3236]),
			.SE(gen[3237]),

			.SELF(gen[3176]),
			.cell_state(gen[3176])
		); 

/******************* CELL 3177 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3177 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3116]),
			.N(gen[3117]),
			.NE(gen[3118]),

			.O(gen[3176]),
			.E(gen[3178]),

			.SO(gen[3236]),
			.S(gen[3237]),
			.SE(gen[3238]),

			.SELF(gen[3177]),
			.cell_state(gen[3177])
		); 

/******************* CELL 3178 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3178 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3117]),
			.N(gen[3118]),
			.NE(gen[3119]),

			.O(gen[3177]),
			.E(gen[3179]),

			.SO(gen[3237]),
			.S(gen[3238]),
			.SE(gen[3239]),

			.SELF(gen[3178]),
			.cell_state(gen[3178])
		); 

/******************* CELL 3179 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3179 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3118]),
			.N(gen[3119]),
			.NE(gen[3118]),

			.O(gen[3178]),
			.E(gen[3178]),

			.SO(gen[3238]),
			.S(gen[3239]),
			.SE(gen[3238]),

			.SELF(gen[3179]),
			.cell_state(gen[3179])
		); 

/******************* CELL 3180 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3180 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3121]),
			.N(gen[3120]),
			.NE(gen[3121]),

			.O(gen[3181]),
			.E(gen[3181]),

			.SO(gen[3241]),
			.S(gen[3240]),
			.SE(gen[3241]),

			.SELF(gen[3180]),
			.cell_state(gen[3180])
		); 

/******************* CELL 3181 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3181 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3120]),
			.N(gen[3121]),
			.NE(gen[3122]),

			.O(gen[3180]),
			.E(gen[3182]),

			.SO(gen[3240]),
			.S(gen[3241]),
			.SE(gen[3242]),

			.SELF(gen[3181]),
			.cell_state(gen[3181])
		); 

/******************* CELL 3182 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3182 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3121]),
			.N(gen[3122]),
			.NE(gen[3123]),

			.O(gen[3181]),
			.E(gen[3183]),

			.SO(gen[3241]),
			.S(gen[3242]),
			.SE(gen[3243]),

			.SELF(gen[3182]),
			.cell_state(gen[3182])
		); 

/******************* CELL 3183 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3183 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3122]),
			.N(gen[3123]),
			.NE(gen[3124]),

			.O(gen[3182]),
			.E(gen[3184]),

			.SO(gen[3242]),
			.S(gen[3243]),
			.SE(gen[3244]),

			.SELF(gen[3183]),
			.cell_state(gen[3183])
		); 

/******************* CELL 3184 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3184 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3123]),
			.N(gen[3124]),
			.NE(gen[3125]),

			.O(gen[3183]),
			.E(gen[3185]),

			.SO(gen[3243]),
			.S(gen[3244]),
			.SE(gen[3245]),

			.SELF(gen[3184]),
			.cell_state(gen[3184])
		); 

/******************* CELL 3185 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3185 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3124]),
			.N(gen[3125]),
			.NE(gen[3126]),

			.O(gen[3184]),
			.E(gen[3186]),

			.SO(gen[3244]),
			.S(gen[3245]),
			.SE(gen[3246]),

			.SELF(gen[3185]),
			.cell_state(gen[3185])
		); 

/******************* CELL 3186 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3186 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3125]),
			.N(gen[3126]),
			.NE(gen[3127]),

			.O(gen[3185]),
			.E(gen[3187]),

			.SO(gen[3245]),
			.S(gen[3246]),
			.SE(gen[3247]),

			.SELF(gen[3186]),
			.cell_state(gen[3186])
		); 

/******************* CELL 3187 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3187 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3126]),
			.N(gen[3127]),
			.NE(gen[3128]),

			.O(gen[3186]),
			.E(gen[3188]),

			.SO(gen[3246]),
			.S(gen[3247]),
			.SE(gen[3248]),

			.SELF(gen[3187]),
			.cell_state(gen[3187])
		); 

/******************* CELL 3188 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3188 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3127]),
			.N(gen[3128]),
			.NE(gen[3129]),

			.O(gen[3187]),
			.E(gen[3189]),

			.SO(gen[3247]),
			.S(gen[3248]),
			.SE(gen[3249]),

			.SELF(gen[3188]),
			.cell_state(gen[3188])
		); 

/******************* CELL 3189 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3189 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3128]),
			.N(gen[3129]),
			.NE(gen[3130]),

			.O(gen[3188]),
			.E(gen[3190]),

			.SO(gen[3248]),
			.S(gen[3249]),
			.SE(gen[3250]),

			.SELF(gen[3189]),
			.cell_state(gen[3189])
		); 

/******************* CELL 3190 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3190 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3129]),
			.N(gen[3130]),
			.NE(gen[3131]),

			.O(gen[3189]),
			.E(gen[3191]),

			.SO(gen[3249]),
			.S(gen[3250]),
			.SE(gen[3251]),

			.SELF(gen[3190]),
			.cell_state(gen[3190])
		); 

/******************* CELL 3191 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3191 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3130]),
			.N(gen[3131]),
			.NE(gen[3132]),

			.O(gen[3190]),
			.E(gen[3192]),

			.SO(gen[3250]),
			.S(gen[3251]),
			.SE(gen[3252]),

			.SELF(gen[3191]),
			.cell_state(gen[3191])
		); 

/******************* CELL 3192 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3192 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3131]),
			.N(gen[3132]),
			.NE(gen[3133]),

			.O(gen[3191]),
			.E(gen[3193]),

			.SO(gen[3251]),
			.S(gen[3252]),
			.SE(gen[3253]),

			.SELF(gen[3192]),
			.cell_state(gen[3192])
		); 

/******************* CELL 3193 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3193 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3132]),
			.N(gen[3133]),
			.NE(gen[3134]),

			.O(gen[3192]),
			.E(gen[3194]),

			.SO(gen[3252]),
			.S(gen[3253]),
			.SE(gen[3254]),

			.SELF(gen[3193]),
			.cell_state(gen[3193])
		); 

/******************* CELL 3194 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3194 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3133]),
			.N(gen[3134]),
			.NE(gen[3135]),

			.O(gen[3193]),
			.E(gen[3195]),

			.SO(gen[3253]),
			.S(gen[3254]),
			.SE(gen[3255]),

			.SELF(gen[3194]),
			.cell_state(gen[3194])
		); 

/******************* CELL 3195 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3195 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3134]),
			.N(gen[3135]),
			.NE(gen[3136]),

			.O(gen[3194]),
			.E(gen[3196]),

			.SO(gen[3254]),
			.S(gen[3255]),
			.SE(gen[3256]),

			.SELF(gen[3195]),
			.cell_state(gen[3195])
		); 

/******************* CELL 3196 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3196 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3135]),
			.N(gen[3136]),
			.NE(gen[3137]),

			.O(gen[3195]),
			.E(gen[3197]),

			.SO(gen[3255]),
			.S(gen[3256]),
			.SE(gen[3257]),

			.SELF(gen[3196]),
			.cell_state(gen[3196])
		); 

/******************* CELL 3197 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3197 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3136]),
			.N(gen[3137]),
			.NE(gen[3138]),

			.O(gen[3196]),
			.E(gen[3198]),

			.SO(gen[3256]),
			.S(gen[3257]),
			.SE(gen[3258]),

			.SELF(gen[3197]),
			.cell_state(gen[3197])
		); 

/******************* CELL 3198 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3198 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3137]),
			.N(gen[3138]),
			.NE(gen[3139]),

			.O(gen[3197]),
			.E(gen[3199]),

			.SO(gen[3257]),
			.S(gen[3258]),
			.SE(gen[3259]),

			.SELF(gen[3198]),
			.cell_state(gen[3198])
		); 

/******************* CELL 3199 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3199 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3138]),
			.N(gen[3139]),
			.NE(gen[3140]),

			.O(gen[3198]),
			.E(gen[3200]),

			.SO(gen[3258]),
			.S(gen[3259]),
			.SE(gen[3260]),

			.SELF(gen[3199]),
			.cell_state(gen[3199])
		); 

/******************* CELL 3200 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3200 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3139]),
			.N(gen[3140]),
			.NE(gen[3141]),

			.O(gen[3199]),
			.E(gen[3201]),

			.SO(gen[3259]),
			.S(gen[3260]),
			.SE(gen[3261]),

			.SELF(gen[3200]),
			.cell_state(gen[3200])
		); 

/******************* CELL 3201 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3201 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3140]),
			.N(gen[3141]),
			.NE(gen[3142]),

			.O(gen[3200]),
			.E(gen[3202]),

			.SO(gen[3260]),
			.S(gen[3261]),
			.SE(gen[3262]),

			.SELF(gen[3201]),
			.cell_state(gen[3201])
		); 

/******************* CELL 3202 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3202 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3141]),
			.N(gen[3142]),
			.NE(gen[3143]),

			.O(gen[3201]),
			.E(gen[3203]),

			.SO(gen[3261]),
			.S(gen[3262]),
			.SE(gen[3263]),

			.SELF(gen[3202]),
			.cell_state(gen[3202])
		); 

/******************* CELL 3203 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3203 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3142]),
			.N(gen[3143]),
			.NE(gen[3144]),

			.O(gen[3202]),
			.E(gen[3204]),

			.SO(gen[3262]),
			.S(gen[3263]),
			.SE(gen[3264]),

			.SELF(gen[3203]),
			.cell_state(gen[3203])
		); 

/******************* CELL 3204 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3204 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3143]),
			.N(gen[3144]),
			.NE(gen[3145]),

			.O(gen[3203]),
			.E(gen[3205]),

			.SO(gen[3263]),
			.S(gen[3264]),
			.SE(gen[3265]),

			.SELF(gen[3204]),
			.cell_state(gen[3204])
		); 

/******************* CELL 3205 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3205 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3144]),
			.N(gen[3145]),
			.NE(gen[3146]),

			.O(gen[3204]),
			.E(gen[3206]),

			.SO(gen[3264]),
			.S(gen[3265]),
			.SE(gen[3266]),

			.SELF(gen[3205]),
			.cell_state(gen[3205])
		); 

/******************* CELL 3206 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3206 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3145]),
			.N(gen[3146]),
			.NE(gen[3147]),

			.O(gen[3205]),
			.E(gen[3207]),

			.SO(gen[3265]),
			.S(gen[3266]),
			.SE(gen[3267]),

			.SELF(gen[3206]),
			.cell_state(gen[3206])
		); 

/******************* CELL 3207 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3207 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3146]),
			.N(gen[3147]),
			.NE(gen[3148]),

			.O(gen[3206]),
			.E(gen[3208]),

			.SO(gen[3266]),
			.S(gen[3267]),
			.SE(gen[3268]),

			.SELF(gen[3207]),
			.cell_state(gen[3207])
		); 

/******************* CELL 3208 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3208 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3147]),
			.N(gen[3148]),
			.NE(gen[3149]),

			.O(gen[3207]),
			.E(gen[3209]),

			.SO(gen[3267]),
			.S(gen[3268]),
			.SE(gen[3269]),

			.SELF(gen[3208]),
			.cell_state(gen[3208])
		); 

/******************* CELL 3209 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3209 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3148]),
			.N(gen[3149]),
			.NE(gen[3150]),

			.O(gen[3208]),
			.E(gen[3210]),

			.SO(gen[3268]),
			.S(gen[3269]),
			.SE(gen[3270]),

			.SELF(gen[3209]),
			.cell_state(gen[3209])
		); 

/******************* CELL 3210 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3210 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3149]),
			.N(gen[3150]),
			.NE(gen[3151]),

			.O(gen[3209]),
			.E(gen[3211]),

			.SO(gen[3269]),
			.S(gen[3270]),
			.SE(gen[3271]),

			.SELF(gen[3210]),
			.cell_state(gen[3210])
		); 

/******************* CELL 3211 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3211 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3150]),
			.N(gen[3151]),
			.NE(gen[3152]),

			.O(gen[3210]),
			.E(gen[3212]),

			.SO(gen[3270]),
			.S(gen[3271]),
			.SE(gen[3272]),

			.SELF(gen[3211]),
			.cell_state(gen[3211])
		); 

/******************* CELL 3212 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3212 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3151]),
			.N(gen[3152]),
			.NE(gen[3153]),

			.O(gen[3211]),
			.E(gen[3213]),

			.SO(gen[3271]),
			.S(gen[3272]),
			.SE(gen[3273]),

			.SELF(gen[3212]),
			.cell_state(gen[3212])
		); 

/******************* CELL 3213 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3213 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3152]),
			.N(gen[3153]),
			.NE(gen[3154]),

			.O(gen[3212]),
			.E(gen[3214]),

			.SO(gen[3272]),
			.S(gen[3273]),
			.SE(gen[3274]),

			.SELF(gen[3213]),
			.cell_state(gen[3213])
		); 

/******************* CELL 3214 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3214 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3153]),
			.N(gen[3154]),
			.NE(gen[3155]),

			.O(gen[3213]),
			.E(gen[3215]),

			.SO(gen[3273]),
			.S(gen[3274]),
			.SE(gen[3275]),

			.SELF(gen[3214]),
			.cell_state(gen[3214])
		); 

/******************* CELL 3215 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3215 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3154]),
			.N(gen[3155]),
			.NE(gen[3156]),

			.O(gen[3214]),
			.E(gen[3216]),

			.SO(gen[3274]),
			.S(gen[3275]),
			.SE(gen[3276]),

			.SELF(gen[3215]),
			.cell_state(gen[3215])
		); 

/******************* CELL 3216 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3216 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3155]),
			.N(gen[3156]),
			.NE(gen[3157]),

			.O(gen[3215]),
			.E(gen[3217]),

			.SO(gen[3275]),
			.S(gen[3276]),
			.SE(gen[3277]),

			.SELF(gen[3216]),
			.cell_state(gen[3216])
		); 

/******************* CELL 3217 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3217 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3156]),
			.N(gen[3157]),
			.NE(gen[3158]),

			.O(gen[3216]),
			.E(gen[3218]),

			.SO(gen[3276]),
			.S(gen[3277]),
			.SE(gen[3278]),

			.SELF(gen[3217]),
			.cell_state(gen[3217])
		); 

/******************* CELL 3218 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3218 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3157]),
			.N(gen[3158]),
			.NE(gen[3159]),

			.O(gen[3217]),
			.E(gen[3219]),

			.SO(gen[3277]),
			.S(gen[3278]),
			.SE(gen[3279]),

			.SELF(gen[3218]),
			.cell_state(gen[3218])
		); 

/******************* CELL 3219 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3219 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3158]),
			.N(gen[3159]),
			.NE(gen[3160]),

			.O(gen[3218]),
			.E(gen[3220]),

			.SO(gen[3278]),
			.S(gen[3279]),
			.SE(gen[3280]),

			.SELF(gen[3219]),
			.cell_state(gen[3219])
		); 

/******************* CELL 3220 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3220 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3159]),
			.N(gen[3160]),
			.NE(gen[3161]),

			.O(gen[3219]),
			.E(gen[3221]),

			.SO(gen[3279]),
			.S(gen[3280]),
			.SE(gen[3281]),

			.SELF(gen[3220]),
			.cell_state(gen[3220])
		); 

/******************* CELL 3221 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3221 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3160]),
			.N(gen[3161]),
			.NE(gen[3162]),

			.O(gen[3220]),
			.E(gen[3222]),

			.SO(gen[3280]),
			.S(gen[3281]),
			.SE(gen[3282]),

			.SELF(gen[3221]),
			.cell_state(gen[3221])
		); 

/******************* CELL 3222 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3222 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3161]),
			.N(gen[3162]),
			.NE(gen[3163]),

			.O(gen[3221]),
			.E(gen[3223]),

			.SO(gen[3281]),
			.S(gen[3282]),
			.SE(gen[3283]),

			.SELF(gen[3222]),
			.cell_state(gen[3222])
		); 

/******************* CELL 3223 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3223 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3162]),
			.N(gen[3163]),
			.NE(gen[3164]),

			.O(gen[3222]),
			.E(gen[3224]),

			.SO(gen[3282]),
			.S(gen[3283]),
			.SE(gen[3284]),

			.SELF(gen[3223]),
			.cell_state(gen[3223])
		); 

/******************* CELL 3224 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3224 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3163]),
			.N(gen[3164]),
			.NE(gen[3165]),

			.O(gen[3223]),
			.E(gen[3225]),

			.SO(gen[3283]),
			.S(gen[3284]),
			.SE(gen[3285]),

			.SELF(gen[3224]),
			.cell_state(gen[3224])
		); 

/******************* CELL 3225 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3225 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3164]),
			.N(gen[3165]),
			.NE(gen[3166]),

			.O(gen[3224]),
			.E(gen[3226]),

			.SO(gen[3284]),
			.S(gen[3285]),
			.SE(gen[3286]),

			.SELF(gen[3225]),
			.cell_state(gen[3225])
		); 

/******************* CELL 3226 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3226 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3165]),
			.N(gen[3166]),
			.NE(gen[3167]),

			.O(gen[3225]),
			.E(gen[3227]),

			.SO(gen[3285]),
			.S(gen[3286]),
			.SE(gen[3287]),

			.SELF(gen[3226]),
			.cell_state(gen[3226])
		); 

/******************* CELL 3227 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3227 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3166]),
			.N(gen[3167]),
			.NE(gen[3168]),

			.O(gen[3226]),
			.E(gen[3228]),

			.SO(gen[3286]),
			.S(gen[3287]),
			.SE(gen[3288]),

			.SELF(gen[3227]),
			.cell_state(gen[3227])
		); 

/******************* CELL 3228 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3228 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3167]),
			.N(gen[3168]),
			.NE(gen[3169]),

			.O(gen[3227]),
			.E(gen[3229]),

			.SO(gen[3287]),
			.S(gen[3288]),
			.SE(gen[3289]),

			.SELF(gen[3228]),
			.cell_state(gen[3228])
		); 

/******************* CELL 3229 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3229 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3168]),
			.N(gen[3169]),
			.NE(gen[3170]),

			.O(gen[3228]),
			.E(gen[3230]),

			.SO(gen[3288]),
			.S(gen[3289]),
			.SE(gen[3290]),

			.SELF(gen[3229]),
			.cell_state(gen[3229])
		); 

/******************* CELL 3230 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3230 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3169]),
			.N(gen[3170]),
			.NE(gen[3171]),

			.O(gen[3229]),
			.E(gen[3231]),

			.SO(gen[3289]),
			.S(gen[3290]),
			.SE(gen[3291]),

			.SELF(gen[3230]),
			.cell_state(gen[3230])
		); 

/******************* CELL 3231 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3231 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3170]),
			.N(gen[3171]),
			.NE(gen[3172]),

			.O(gen[3230]),
			.E(gen[3232]),

			.SO(gen[3290]),
			.S(gen[3291]),
			.SE(gen[3292]),

			.SELF(gen[3231]),
			.cell_state(gen[3231])
		); 

/******************* CELL 3232 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3232 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3171]),
			.N(gen[3172]),
			.NE(gen[3173]),

			.O(gen[3231]),
			.E(gen[3233]),

			.SO(gen[3291]),
			.S(gen[3292]),
			.SE(gen[3293]),

			.SELF(gen[3232]),
			.cell_state(gen[3232])
		); 

/******************* CELL 3233 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3233 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3172]),
			.N(gen[3173]),
			.NE(gen[3174]),

			.O(gen[3232]),
			.E(gen[3234]),

			.SO(gen[3292]),
			.S(gen[3293]),
			.SE(gen[3294]),

			.SELF(gen[3233]),
			.cell_state(gen[3233])
		); 

/******************* CELL 3234 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3234 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3173]),
			.N(gen[3174]),
			.NE(gen[3175]),

			.O(gen[3233]),
			.E(gen[3235]),

			.SO(gen[3293]),
			.S(gen[3294]),
			.SE(gen[3295]),

			.SELF(gen[3234]),
			.cell_state(gen[3234])
		); 

/******************* CELL 3235 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3235 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3174]),
			.N(gen[3175]),
			.NE(gen[3176]),

			.O(gen[3234]),
			.E(gen[3236]),

			.SO(gen[3294]),
			.S(gen[3295]),
			.SE(gen[3296]),

			.SELF(gen[3235]),
			.cell_state(gen[3235])
		); 

/******************* CELL 3236 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3236 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3175]),
			.N(gen[3176]),
			.NE(gen[3177]),

			.O(gen[3235]),
			.E(gen[3237]),

			.SO(gen[3295]),
			.S(gen[3296]),
			.SE(gen[3297]),

			.SELF(gen[3236]),
			.cell_state(gen[3236])
		); 

/******************* CELL 3237 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3237 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3176]),
			.N(gen[3177]),
			.NE(gen[3178]),

			.O(gen[3236]),
			.E(gen[3238]),

			.SO(gen[3296]),
			.S(gen[3297]),
			.SE(gen[3298]),

			.SELF(gen[3237]),
			.cell_state(gen[3237])
		); 

/******************* CELL 3238 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3238 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3177]),
			.N(gen[3178]),
			.NE(gen[3179]),

			.O(gen[3237]),
			.E(gen[3239]),

			.SO(gen[3297]),
			.S(gen[3298]),
			.SE(gen[3299]),

			.SELF(gen[3238]),
			.cell_state(gen[3238])
		); 

/******************* CELL 3239 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3239 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3178]),
			.N(gen[3179]),
			.NE(gen[3178]),

			.O(gen[3238]),
			.E(gen[3238]),

			.SO(gen[3298]),
			.S(gen[3299]),
			.SE(gen[3298]),

			.SELF(gen[3239]),
			.cell_state(gen[3239])
		); 

/******************* CELL 3240 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3240 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3181]),
			.N(gen[3180]),
			.NE(gen[3181]),

			.O(gen[3241]),
			.E(gen[3241]),

			.SO(gen[3301]),
			.S(gen[3300]),
			.SE(gen[3301]),

			.SELF(gen[3240]),
			.cell_state(gen[3240])
		); 

/******************* CELL 3241 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3241 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3180]),
			.N(gen[3181]),
			.NE(gen[3182]),

			.O(gen[3240]),
			.E(gen[3242]),

			.SO(gen[3300]),
			.S(gen[3301]),
			.SE(gen[3302]),

			.SELF(gen[3241]),
			.cell_state(gen[3241])
		); 

/******************* CELL 3242 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3242 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3181]),
			.N(gen[3182]),
			.NE(gen[3183]),

			.O(gen[3241]),
			.E(gen[3243]),

			.SO(gen[3301]),
			.S(gen[3302]),
			.SE(gen[3303]),

			.SELF(gen[3242]),
			.cell_state(gen[3242])
		); 

/******************* CELL 3243 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3243 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3182]),
			.N(gen[3183]),
			.NE(gen[3184]),

			.O(gen[3242]),
			.E(gen[3244]),

			.SO(gen[3302]),
			.S(gen[3303]),
			.SE(gen[3304]),

			.SELF(gen[3243]),
			.cell_state(gen[3243])
		); 

/******************* CELL 3244 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3244 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3183]),
			.N(gen[3184]),
			.NE(gen[3185]),

			.O(gen[3243]),
			.E(gen[3245]),

			.SO(gen[3303]),
			.S(gen[3304]),
			.SE(gen[3305]),

			.SELF(gen[3244]),
			.cell_state(gen[3244])
		); 

/******************* CELL 3245 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3245 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3184]),
			.N(gen[3185]),
			.NE(gen[3186]),

			.O(gen[3244]),
			.E(gen[3246]),

			.SO(gen[3304]),
			.S(gen[3305]),
			.SE(gen[3306]),

			.SELF(gen[3245]),
			.cell_state(gen[3245])
		); 

/******************* CELL 3246 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3246 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3185]),
			.N(gen[3186]),
			.NE(gen[3187]),

			.O(gen[3245]),
			.E(gen[3247]),

			.SO(gen[3305]),
			.S(gen[3306]),
			.SE(gen[3307]),

			.SELF(gen[3246]),
			.cell_state(gen[3246])
		); 

/******************* CELL 3247 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3247 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3186]),
			.N(gen[3187]),
			.NE(gen[3188]),

			.O(gen[3246]),
			.E(gen[3248]),

			.SO(gen[3306]),
			.S(gen[3307]),
			.SE(gen[3308]),

			.SELF(gen[3247]),
			.cell_state(gen[3247])
		); 

/******************* CELL 3248 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3248 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3187]),
			.N(gen[3188]),
			.NE(gen[3189]),

			.O(gen[3247]),
			.E(gen[3249]),

			.SO(gen[3307]),
			.S(gen[3308]),
			.SE(gen[3309]),

			.SELF(gen[3248]),
			.cell_state(gen[3248])
		); 

/******************* CELL 3249 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3249 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3188]),
			.N(gen[3189]),
			.NE(gen[3190]),

			.O(gen[3248]),
			.E(gen[3250]),

			.SO(gen[3308]),
			.S(gen[3309]),
			.SE(gen[3310]),

			.SELF(gen[3249]),
			.cell_state(gen[3249])
		); 

/******************* CELL 3250 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3250 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3189]),
			.N(gen[3190]),
			.NE(gen[3191]),

			.O(gen[3249]),
			.E(gen[3251]),

			.SO(gen[3309]),
			.S(gen[3310]),
			.SE(gen[3311]),

			.SELF(gen[3250]),
			.cell_state(gen[3250])
		); 

/******************* CELL 3251 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3251 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3190]),
			.N(gen[3191]),
			.NE(gen[3192]),

			.O(gen[3250]),
			.E(gen[3252]),

			.SO(gen[3310]),
			.S(gen[3311]),
			.SE(gen[3312]),

			.SELF(gen[3251]),
			.cell_state(gen[3251])
		); 

/******************* CELL 3252 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3252 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3191]),
			.N(gen[3192]),
			.NE(gen[3193]),

			.O(gen[3251]),
			.E(gen[3253]),

			.SO(gen[3311]),
			.S(gen[3312]),
			.SE(gen[3313]),

			.SELF(gen[3252]),
			.cell_state(gen[3252])
		); 

/******************* CELL 3253 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3253 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3192]),
			.N(gen[3193]),
			.NE(gen[3194]),

			.O(gen[3252]),
			.E(gen[3254]),

			.SO(gen[3312]),
			.S(gen[3313]),
			.SE(gen[3314]),

			.SELF(gen[3253]),
			.cell_state(gen[3253])
		); 

/******************* CELL 3254 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3254 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3193]),
			.N(gen[3194]),
			.NE(gen[3195]),

			.O(gen[3253]),
			.E(gen[3255]),

			.SO(gen[3313]),
			.S(gen[3314]),
			.SE(gen[3315]),

			.SELF(gen[3254]),
			.cell_state(gen[3254])
		); 

/******************* CELL 3255 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3255 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3194]),
			.N(gen[3195]),
			.NE(gen[3196]),

			.O(gen[3254]),
			.E(gen[3256]),

			.SO(gen[3314]),
			.S(gen[3315]),
			.SE(gen[3316]),

			.SELF(gen[3255]),
			.cell_state(gen[3255])
		); 

/******************* CELL 3256 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3256 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3195]),
			.N(gen[3196]),
			.NE(gen[3197]),

			.O(gen[3255]),
			.E(gen[3257]),

			.SO(gen[3315]),
			.S(gen[3316]),
			.SE(gen[3317]),

			.SELF(gen[3256]),
			.cell_state(gen[3256])
		); 

/******************* CELL 3257 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3257 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3196]),
			.N(gen[3197]),
			.NE(gen[3198]),

			.O(gen[3256]),
			.E(gen[3258]),

			.SO(gen[3316]),
			.S(gen[3317]),
			.SE(gen[3318]),

			.SELF(gen[3257]),
			.cell_state(gen[3257])
		); 

/******************* CELL 3258 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3258 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3197]),
			.N(gen[3198]),
			.NE(gen[3199]),

			.O(gen[3257]),
			.E(gen[3259]),

			.SO(gen[3317]),
			.S(gen[3318]),
			.SE(gen[3319]),

			.SELF(gen[3258]),
			.cell_state(gen[3258])
		); 

/******************* CELL 3259 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3259 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3198]),
			.N(gen[3199]),
			.NE(gen[3200]),

			.O(gen[3258]),
			.E(gen[3260]),

			.SO(gen[3318]),
			.S(gen[3319]),
			.SE(gen[3320]),

			.SELF(gen[3259]),
			.cell_state(gen[3259])
		); 

/******************* CELL 3260 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3260 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3199]),
			.N(gen[3200]),
			.NE(gen[3201]),

			.O(gen[3259]),
			.E(gen[3261]),

			.SO(gen[3319]),
			.S(gen[3320]),
			.SE(gen[3321]),

			.SELF(gen[3260]),
			.cell_state(gen[3260])
		); 

/******************* CELL 3261 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3261 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3200]),
			.N(gen[3201]),
			.NE(gen[3202]),

			.O(gen[3260]),
			.E(gen[3262]),

			.SO(gen[3320]),
			.S(gen[3321]),
			.SE(gen[3322]),

			.SELF(gen[3261]),
			.cell_state(gen[3261])
		); 

/******************* CELL 3262 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3262 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3201]),
			.N(gen[3202]),
			.NE(gen[3203]),

			.O(gen[3261]),
			.E(gen[3263]),

			.SO(gen[3321]),
			.S(gen[3322]),
			.SE(gen[3323]),

			.SELF(gen[3262]),
			.cell_state(gen[3262])
		); 

/******************* CELL 3263 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3263 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3202]),
			.N(gen[3203]),
			.NE(gen[3204]),

			.O(gen[3262]),
			.E(gen[3264]),

			.SO(gen[3322]),
			.S(gen[3323]),
			.SE(gen[3324]),

			.SELF(gen[3263]),
			.cell_state(gen[3263])
		); 

/******************* CELL 3264 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3264 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3203]),
			.N(gen[3204]),
			.NE(gen[3205]),

			.O(gen[3263]),
			.E(gen[3265]),

			.SO(gen[3323]),
			.S(gen[3324]),
			.SE(gen[3325]),

			.SELF(gen[3264]),
			.cell_state(gen[3264])
		); 

/******************* CELL 3265 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3265 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3204]),
			.N(gen[3205]),
			.NE(gen[3206]),

			.O(gen[3264]),
			.E(gen[3266]),

			.SO(gen[3324]),
			.S(gen[3325]),
			.SE(gen[3326]),

			.SELF(gen[3265]),
			.cell_state(gen[3265])
		); 

/******************* CELL 3266 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3266 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3205]),
			.N(gen[3206]),
			.NE(gen[3207]),

			.O(gen[3265]),
			.E(gen[3267]),

			.SO(gen[3325]),
			.S(gen[3326]),
			.SE(gen[3327]),

			.SELF(gen[3266]),
			.cell_state(gen[3266])
		); 

/******************* CELL 3267 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3267 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3206]),
			.N(gen[3207]),
			.NE(gen[3208]),

			.O(gen[3266]),
			.E(gen[3268]),

			.SO(gen[3326]),
			.S(gen[3327]),
			.SE(gen[3328]),

			.SELF(gen[3267]),
			.cell_state(gen[3267])
		); 

/******************* CELL 3268 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3268 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3207]),
			.N(gen[3208]),
			.NE(gen[3209]),

			.O(gen[3267]),
			.E(gen[3269]),

			.SO(gen[3327]),
			.S(gen[3328]),
			.SE(gen[3329]),

			.SELF(gen[3268]),
			.cell_state(gen[3268])
		); 

/******************* CELL 3269 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3269 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3208]),
			.N(gen[3209]),
			.NE(gen[3210]),

			.O(gen[3268]),
			.E(gen[3270]),

			.SO(gen[3328]),
			.S(gen[3329]),
			.SE(gen[3330]),

			.SELF(gen[3269]),
			.cell_state(gen[3269])
		); 

/******************* CELL 3270 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3270 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3209]),
			.N(gen[3210]),
			.NE(gen[3211]),

			.O(gen[3269]),
			.E(gen[3271]),

			.SO(gen[3329]),
			.S(gen[3330]),
			.SE(gen[3331]),

			.SELF(gen[3270]),
			.cell_state(gen[3270])
		); 

/******************* CELL 3271 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3271 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3210]),
			.N(gen[3211]),
			.NE(gen[3212]),

			.O(gen[3270]),
			.E(gen[3272]),

			.SO(gen[3330]),
			.S(gen[3331]),
			.SE(gen[3332]),

			.SELF(gen[3271]),
			.cell_state(gen[3271])
		); 

/******************* CELL 3272 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3272 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3211]),
			.N(gen[3212]),
			.NE(gen[3213]),

			.O(gen[3271]),
			.E(gen[3273]),

			.SO(gen[3331]),
			.S(gen[3332]),
			.SE(gen[3333]),

			.SELF(gen[3272]),
			.cell_state(gen[3272])
		); 

/******************* CELL 3273 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3273 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3212]),
			.N(gen[3213]),
			.NE(gen[3214]),

			.O(gen[3272]),
			.E(gen[3274]),

			.SO(gen[3332]),
			.S(gen[3333]),
			.SE(gen[3334]),

			.SELF(gen[3273]),
			.cell_state(gen[3273])
		); 

/******************* CELL 3274 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3274 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3213]),
			.N(gen[3214]),
			.NE(gen[3215]),

			.O(gen[3273]),
			.E(gen[3275]),

			.SO(gen[3333]),
			.S(gen[3334]),
			.SE(gen[3335]),

			.SELF(gen[3274]),
			.cell_state(gen[3274])
		); 

/******************* CELL 3275 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3275 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3214]),
			.N(gen[3215]),
			.NE(gen[3216]),

			.O(gen[3274]),
			.E(gen[3276]),

			.SO(gen[3334]),
			.S(gen[3335]),
			.SE(gen[3336]),

			.SELF(gen[3275]),
			.cell_state(gen[3275])
		); 

/******************* CELL 3276 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3276 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3215]),
			.N(gen[3216]),
			.NE(gen[3217]),

			.O(gen[3275]),
			.E(gen[3277]),

			.SO(gen[3335]),
			.S(gen[3336]),
			.SE(gen[3337]),

			.SELF(gen[3276]),
			.cell_state(gen[3276])
		); 

/******************* CELL 3277 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3277 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3216]),
			.N(gen[3217]),
			.NE(gen[3218]),

			.O(gen[3276]),
			.E(gen[3278]),

			.SO(gen[3336]),
			.S(gen[3337]),
			.SE(gen[3338]),

			.SELF(gen[3277]),
			.cell_state(gen[3277])
		); 

/******************* CELL 3278 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3278 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3217]),
			.N(gen[3218]),
			.NE(gen[3219]),

			.O(gen[3277]),
			.E(gen[3279]),

			.SO(gen[3337]),
			.S(gen[3338]),
			.SE(gen[3339]),

			.SELF(gen[3278]),
			.cell_state(gen[3278])
		); 

/******************* CELL 3279 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3279 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3218]),
			.N(gen[3219]),
			.NE(gen[3220]),

			.O(gen[3278]),
			.E(gen[3280]),

			.SO(gen[3338]),
			.S(gen[3339]),
			.SE(gen[3340]),

			.SELF(gen[3279]),
			.cell_state(gen[3279])
		); 

/******************* CELL 3280 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3280 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3219]),
			.N(gen[3220]),
			.NE(gen[3221]),

			.O(gen[3279]),
			.E(gen[3281]),

			.SO(gen[3339]),
			.S(gen[3340]),
			.SE(gen[3341]),

			.SELF(gen[3280]),
			.cell_state(gen[3280])
		); 

/******************* CELL 3281 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3281 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3220]),
			.N(gen[3221]),
			.NE(gen[3222]),

			.O(gen[3280]),
			.E(gen[3282]),

			.SO(gen[3340]),
			.S(gen[3341]),
			.SE(gen[3342]),

			.SELF(gen[3281]),
			.cell_state(gen[3281])
		); 

/******************* CELL 3282 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3282 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3221]),
			.N(gen[3222]),
			.NE(gen[3223]),

			.O(gen[3281]),
			.E(gen[3283]),

			.SO(gen[3341]),
			.S(gen[3342]),
			.SE(gen[3343]),

			.SELF(gen[3282]),
			.cell_state(gen[3282])
		); 

/******************* CELL 3283 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3283 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3222]),
			.N(gen[3223]),
			.NE(gen[3224]),

			.O(gen[3282]),
			.E(gen[3284]),

			.SO(gen[3342]),
			.S(gen[3343]),
			.SE(gen[3344]),

			.SELF(gen[3283]),
			.cell_state(gen[3283])
		); 

/******************* CELL 3284 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3284 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3223]),
			.N(gen[3224]),
			.NE(gen[3225]),

			.O(gen[3283]),
			.E(gen[3285]),

			.SO(gen[3343]),
			.S(gen[3344]),
			.SE(gen[3345]),

			.SELF(gen[3284]),
			.cell_state(gen[3284])
		); 

/******************* CELL 3285 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3285 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3224]),
			.N(gen[3225]),
			.NE(gen[3226]),

			.O(gen[3284]),
			.E(gen[3286]),

			.SO(gen[3344]),
			.S(gen[3345]),
			.SE(gen[3346]),

			.SELF(gen[3285]),
			.cell_state(gen[3285])
		); 

/******************* CELL 3286 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3286 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3225]),
			.N(gen[3226]),
			.NE(gen[3227]),

			.O(gen[3285]),
			.E(gen[3287]),

			.SO(gen[3345]),
			.S(gen[3346]),
			.SE(gen[3347]),

			.SELF(gen[3286]),
			.cell_state(gen[3286])
		); 

/******************* CELL 3287 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3287 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3226]),
			.N(gen[3227]),
			.NE(gen[3228]),

			.O(gen[3286]),
			.E(gen[3288]),

			.SO(gen[3346]),
			.S(gen[3347]),
			.SE(gen[3348]),

			.SELF(gen[3287]),
			.cell_state(gen[3287])
		); 

/******************* CELL 3288 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3288 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3227]),
			.N(gen[3228]),
			.NE(gen[3229]),

			.O(gen[3287]),
			.E(gen[3289]),

			.SO(gen[3347]),
			.S(gen[3348]),
			.SE(gen[3349]),

			.SELF(gen[3288]),
			.cell_state(gen[3288])
		); 

/******************* CELL 3289 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3289 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3228]),
			.N(gen[3229]),
			.NE(gen[3230]),

			.O(gen[3288]),
			.E(gen[3290]),

			.SO(gen[3348]),
			.S(gen[3349]),
			.SE(gen[3350]),

			.SELF(gen[3289]),
			.cell_state(gen[3289])
		); 

/******************* CELL 3290 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3290 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3229]),
			.N(gen[3230]),
			.NE(gen[3231]),

			.O(gen[3289]),
			.E(gen[3291]),

			.SO(gen[3349]),
			.S(gen[3350]),
			.SE(gen[3351]),

			.SELF(gen[3290]),
			.cell_state(gen[3290])
		); 

/******************* CELL 3291 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3291 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3230]),
			.N(gen[3231]),
			.NE(gen[3232]),

			.O(gen[3290]),
			.E(gen[3292]),

			.SO(gen[3350]),
			.S(gen[3351]),
			.SE(gen[3352]),

			.SELF(gen[3291]),
			.cell_state(gen[3291])
		); 

/******************* CELL 3292 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3292 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3231]),
			.N(gen[3232]),
			.NE(gen[3233]),

			.O(gen[3291]),
			.E(gen[3293]),

			.SO(gen[3351]),
			.S(gen[3352]),
			.SE(gen[3353]),

			.SELF(gen[3292]),
			.cell_state(gen[3292])
		); 

/******************* CELL 3293 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3293 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3232]),
			.N(gen[3233]),
			.NE(gen[3234]),

			.O(gen[3292]),
			.E(gen[3294]),

			.SO(gen[3352]),
			.S(gen[3353]),
			.SE(gen[3354]),

			.SELF(gen[3293]),
			.cell_state(gen[3293])
		); 

/******************* CELL 3294 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3294 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3233]),
			.N(gen[3234]),
			.NE(gen[3235]),

			.O(gen[3293]),
			.E(gen[3295]),

			.SO(gen[3353]),
			.S(gen[3354]),
			.SE(gen[3355]),

			.SELF(gen[3294]),
			.cell_state(gen[3294])
		); 

/******************* CELL 3295 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3295 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3234]),
			.N(gen[3235]),
			.NE(gen[3236]),

			.O(gen[3294]),
			.E(gen[3296]),

			.SO(gen[3354]),
			.S(gen[3355]),
			.SE(gen[3356]),

			.SELF(gen[3295]),
			.cell_state(gen[3295])
		); 

/******************* CELL 3296 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3296 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3235]),
			.N(gen[3236]),
			.NE(gen[3237]),

			.O(gen[3295]),
			.E(gen[3297]),

			.SO(gen[3355]),
			.S(gen[3356]),
			.SE(gen[3357]),

			.SELF(gen[3296]),
			.cell_state(gen[3296])
		); 

/******************* CELL 3297 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3297 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3236]),
			.N(gen[3237]),
			.NE(gen[3238]),

			.O(gen[3296]),
			.E(gen[3298]),

			.SO(gen[3356]),
			.S(gen[3357]),
			.SE(gen[3358]),

			.SELF(gen[3297]),
			.cell_state(gen[3297])
		); 

/******************* CELL 3298 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3298 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3237]),
			.N(gen[3238]),
			.NE(gen[3239]),

			.O(gen[3297]),
			.E(gen[3299]),

			.SO(gen[3357]),
			.S(gen[3358]),
			.SE(gen[3359]),

			.SELF(gen[3298]),
			.cell_state(gen[3298])
		); 

/******************* CELL 3299 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3299 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3238]),
			.N(gen[3239]),
			.NE(gen[3238]),

			.O(gen[3298]),
			.E(gen[3298]),

			.SO(gen[3358]),
			.S(gen[3359]),
			.SE(gen[3358]),

			.SELF(gen[3299]),
			.cell_state(gen[3299])
		); 

/******************* CELL 3300 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3300 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3241]),
			.N(gen[3240]),
			.NE(gen[3241]),

			.O(gen[3301]),
			.E(gen[3301]),

			.SO(gen[3361]),
			.S(gen[3360]),
			.SE(gen[3361]),

			.SELF(gen[3300]),
			.cell_state(gen[3300])
		); 

/******************* CELL 3301 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3301 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3240]),
			.N(gen[3241]),
			.NE(gen[3242]),

			.O(gen[3300]),
			.E(gen[3302]),

			.SO(gen[3360]),
			.S(gen[3361]),
			.SE(gen[3362]),

			.SELF(gen[3301]),
			.cell_state(gen[3301])
		); 

/******************* CELL 3302 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3302 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3241]),
			.N(gen[3242]),
			.NE(gen[3243]),

			.O(gen[3301]),
			.E(gen[3303]),

			.SO(gen[3361]),
			.S(gen[3362]),
			.SE(gen[3363]),

			.SELF(gen[3302]),
			.cell_state(gen[3302])
		); 

/******************* CELL 3303 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3303 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3242]),
			.N(gen[3243]),
			.NE(gen[3244]),

			.O(gen[3302]),
			.E(gen[3304]),

			.SO(gen[3362]),
			.S(gen[3363]),
			.SE(gen[3364]),

			.SELF(gen[3303]),
			.cell_state(gen[3303])
		); 

/******************* CELL 3304 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3304 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3243]),
			.N(gen[3244]),
			.NE(gen[3245]),

			.O(gen[3303]),
			.E(gen[3305]),

			.SO(gen[3363]),
			.S(gen[3364]),
			.SE(gen[3365]),

			.SELF(gen[3304]),
			.cell_state(gen[3304])
		); 

/******************* CELL 3305 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3305 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3244]),
			.N(gen[3245]),
			.NE(gen[3246]),

			.O(gen[3304]),
			.E(gen[3306]),

			.SO(gen[3364]),
			.S(gen[3365]),
			.SE(gen[3366]),

			.SELF(gen[3305]),
			.cell_state(gen[3305])
		); 

/******************* CELL 3306 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3306 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3245]),
			.N(gen[3246]),
			.NE(gen[3247]),

			.O(gen[3305]),
			.E(gen[3307]),

			.SO(gen[3365]),
			.S(gen[3366]),
			.SE(gen[3367]),

			.SELF(gen[3306]),
			.cell_state(gen[3306])
		); 

/******************* CELL 3307 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3307 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3246]),
			.N(gen[3247]),
			.NE(gen[3248]),

			.O(gen[3306]),
			.E(gen[3308]),

			.SO(gen[3366]),
			.S(gen[3367]),
			.SE(gen[3368]),

			.SELF(gen[3307]),
			.cell_state(gen[3307])
		); 

/******************* CELL 3308 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3308 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3247]),
			.N(gen[3248]),
			.NE(gen[3249]),

			.O(gen[3307]),
			.E(gen[3309]),

			.SO(gen[3367]),
			.S(gen[3368]),
			.SE(gen[3369]),

			.SELF(gen[3308]),
			.cell_state(gen[3308])
		); 

/******************* CELL 3309 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3309 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3248]),
			.N(gen[3249]),
			.NE(gen[3250]),

			.O(gen[3308]),
			.E(gen[3310]),

			.SO(gen[3368]),
			.S(gen[3369]),
			.SE(gen[3370]),

			.SELF(gen[3309]),
			.cell_state(gen[3309])
		); 

/******************* CELL 3310 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3310 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3249]),
			.N(gen[3250]),
			.NE(gen[3251]),

			.O(gen[3309]),
			.E(gen[3311]),

			.SO(gen[3369]),
			.S(gen[3370]),
			.SE(gen[3371]),

			.SELF(gen[3310]),
			.cell_state(gen[3310])
		); 

/******************* CELL 3311 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3311 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3250]),
			.N(gen[3251]),
			.NE(gen[3252]),

			.O(gen[3310]),
			.E(gen[3312]),

			.SO(gen[3370]),
			.S(gen[3371]),
			.SE(gen[3372]),

			.SELF(gen[3311]),
			.cell_state(gen[3311])
		); 

/******************* CELL 3312 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3312 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3251]),
			.N(gen[3252]),
			.NE(gen[3253]),

			.O(gen[3311]),
			.E(gen[3313]),

			.SO(gen[3371]),
			.S(gen[3372]),
			.SE(gen[3373]),

			.SELF(gen[3312]),
			.cell_state(gen[3312])
		); 

/******************* CELL 3313 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3313 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3252]),
			.N(gen[3253]),
			.NE(gen[3254]),

			.O(gen[3312]),
			.E(gen[3314]),

			.SO(gen[3372]),
			.S(gen[3373]),
			.SE(gen[3374]),

			.SELF(gen[3313]),
			.cell_state(gen[3313])
		); 

/******************* CELL 3314 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3314 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3253]),
			.N(gen[3254]),
			.NE(gen[3255]),

			.O(gen[3313]),
			.E(gen[3315]),

			.SO(gen[3373]),
			.S(gen[3374]),
			.SE(gen[3375]),

			.SELF(gen[3314]),
			.cell_state(gen[3314])
		); 

/******************* CELL 3315 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3315 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3254]),
			.N(gen[3255]),
			.NE(gen[3256]),

			.O(gen[3314]),
			.E(gen[3316]),

			.SO(gen[3374]),
			.S(gen[3375]),
			.SE(gen[3376]),

			.SELF(gen[3315]),
			.cell_state(gen[3315])
		); 

/******************* CELL 3316 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3316 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3255]),
			.N(gen[3256]),
			.NE(gen[3257]),

			.O(gen[3315]),
			.E(gen[3317]),

			.SO(gen[3375]),
			.S(gen[3376]),
			.SE(gen[3377]),

			.SELF(gen[3316]),
			.cell_state(gen[3316])
		); 

/******************* CELL 3317 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3317 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3256]),
			.N(gen[3257]),
			.NE(gen[3258]),

			.O(gen[3316]),
			.E(gen[3318]),

			.SO(gen[3376]),
			.S(gen[3377]),
			.SE(gen[3378]),

			.SELF(gen[3317]),
			.cell_state(gen[3317])
		); 

/******************* CELL 3318 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3318 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3257]),
			.N(gen[3258]),
			.NE(gen[3259]),

			.O(gen[3317]),
			.E(gen[3319]),

			.SO(gen[3377]),
			.S(gen[3378]),
			.SE(gen[3379]),

			.SELF(gen[3318]),
			.cell_state(gen[3318])
		); 

/******************* CELL 3319 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3319 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3258]),
			.N(gen[3259]),
			.NE(gen[3260]),

			.O(gen[3318]),
			.E(gen[3320]),

			.SO(gen[3378]),
			.S(gen[3379]),
			.SE(gen[3380]),

			.SELF(gen[3319]),
			.cell_state(gen[3319])
		); 

/******************* CELL 3320 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3320 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3259]),
			.N(gen[3260]),
			.NE(gen[3261]),

			.O(gen[3319]),
			.E(gen[3321]),

			.SO(gen[3379]),
			.S(gen[3380]),
			.SE(gen[3381]),

			.SELF(gen[3320]),
			.cell_state(gen[3320])
		); 

/******************* CELL 3321 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3321 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3260]),
			.N(gen[3261]),
			.NE(gen[3262]),

			.O(gen[3320]),
			.E(gen[3322]),

			.SO(gen[3380]),
			.S(gen[3381]),
			.SE(gen[3382]),

			.SELF(gen[3321]),
			.cell_state(gen[3321])
		); 

/******************* CELL 3322 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3322 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3261]),
			.N(gen[3262]),
			.NE(gen[3263]),

			.O(gen[3321]),
			.E(gen[3323]),

			.SO(gen[3381]),
			.S(gen[3382]),
			.SE(gen[3383]),

			.SELF(gen[3322]),
			.cell_state(gen[3322])
		); 

/******************* CELL 3323 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3323 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3262]),
			.N(gen[3263]),
			.NE(gen[3264]),

			.O(gen[3322]),
			.E(gen[3324]),

			.SO(gen[3382]),
			.S(gen[3383]),
			.SE(gen[3384]),

			.SELF(gen[3323]),
			.cell_state(gen[3323])
		); 

/******************* CELL 3324 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3324 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3263]),
			.N(gen[3264]),
			.NE(gen[3265]),

			.O(gen[3323]),
			.E(gen[3325]),

			.SO(gen[3383]),
			.S(gen[3384]),
			.SE(gen[3385]),

			.SELF(gen[3324]),
			.cell_state(gen[3324])
		); 

/******************* CELL 3325 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3325 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3264]),
			.N(gen[3265]),
			.NE(gen[3266]),

			.O(gen[3324]),
			.E(gen[3326]),

			.SO(gen[3384]),
			.S(gen[3385]),
			.SE(gen[3386]),

			.SELF(gen[3325]),
			.cell_state(gen[3325])
		); 

/******************* CELL 3326 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3326 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3265]),
			.N(gen[3266]),
			.NE(gen[3267]),

			.O(gen[3325]),
			.E(gen[3327]),

			.SO(gen[3385]),
			.S(gen[3386]),
			.SE(gen[3387]),

			.SELF(gen[3326]),
			.cell_state(gen[3326])
		); 

/******************* CELL 3327 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3327 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3266]),
			.N(gen[3267]),
			.NE(gen[3268]),

			.O(gen[3326]),
			.E(gen[3328]),

			.SO(gen[3386]),
			.S(gen[3387]),
			.SE(gen[3388]),

			.SELF(gen[3327]),
			.cell_state(gen[3327])
		); 

/******************* CELL 3328 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3328 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3267]),
			.N(gen[3268]),
			.NE(gen[3269]),

			.O(gen[3327]),
			.E(gen[3329]),

			.SO(gen[3387]),
			.S(gen[3388]),
			.SE(gen[3389]),

			.SELF(gen[3328]),
			.cell_state(gen[3328])
		); 

/******************* CELL 3329 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3329 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3268]),
			.N(gen[3269]),
			.NE(gen[3270]),

			.O(gen[3328]),
			.E(gen[3330]),

			.SO(gen[3388]),
			.S(gen[3389]),
			.SE(gen[3390]),

			.SELF(gen[3329]),
			.cell_state(gen[3329])
		); 

/******************* CELL 3330 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3330 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3269]),
			.N(gen[3270]),
			.NE(gen[3271]),

			.O(gen[3329]),
			.E(gen[3331]),

			.SO(gen[3389]),
			.S(gen[3390]),
			.SE(gen[3391]),

			.SELF(gen[3330]),
			.cell_state(gen[3330])
		); 

/******************* CELL 3331 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3331 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3270]),
			.N(gen[3271]),
			.NE(gen[3272]),

			.O(gen[3330]),
			.E(gen[3332]),

			.SO(gen[3390]),
			.S(gen[3391]),
			.SE(gen[3392]),

			.SELF(gen[3331]),
			.cell_state(gen[3331])
		); 

/******************* CELL 3332 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3332 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3271]),
			.N(gen[3272]),
			.NE(gen[3273]),

			.O(gen[3331]),
			.E(gen[3333]),

			.SO(gen[3391]),
			.S(gen[3392]),
			.SE(gen[3393]),

			.SELF(gen[3332]),
			.cell_state(gen[3332])
		); 

/******************* CELL 3333 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3333 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3272]),
			.N(gen[3273]),
			.NE(gen[3274]),

			.O(gen[3332]),
			.E(gen[3334]),

			.SO(gen[3392]),
			.S(gen[3393]),
			.SE(gen[3394]),

			.SELF(gen[3333]),
			.cell_state(gen[3333])
		); 

/******************* CELL 3334 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3334 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3273]),
			.N(gen[3274]),
			.NE(gen[3275]),

			.O(gen[3333]),
			.E(gen[3335]),

			.SO(gen[3393]),
			.S(gen[3394]),
			.SE(gen[3395]),

			.SELF(gen[3334]),
			.cell_state(gen[3334])
		); 

/******************* CELL 3335 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3335 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3274]),
			.N(gen[3275]),
			.NE(gen[3276]),

			.O(gen[3334]),
			.E(gen[3336]),

			.SO(gen[3394]),
			.S(gen[3395]),
			.SE(gen[3396]),

			.SELF(gen[3335]),
			.cell_state(gen[3335])
		); 

/******************* CELL 3336 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3336 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3275]),
			.N(gen[3276]),
			.NE(gen[3277]),

			.O(gen[3335]),
			.E(gen[3337]),

			.SO(gen[3395]),
			.S(gen[3396]),
			.SE(gen[3397]),

			.SELF(gen[3336]),
			.cell_state(gen[3336])
		); 

/******************* CELL 3337 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3337 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3276]),
			.N(gen[3277]),
			.NE(gen[3278]),

			.O(gen[3336]),
			.E(gen[3338]),

			.SO(gen[3396]),
			.S(gen[3397]),
			.SE(gen[3398]),

			.SELF(gen[3337]),
			.cell_state(gen[3337])
		); 

/******************* CELL 3338 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3338 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3277]),
			.N(gen[3278]),
			.NE(gen[3279]),

			.O(gen[3337]),
			.E(gen[3339]),

			.SO(gen[3397]),
			.S(gen[3398]),
			.SE(gen[3399]),

			.SELF(gen[3338]),
			.cell_state(gen[3338])
		); 

/******************* CELL 3339 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3339 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3278]),
			.N(gen[3279]),
			.NE(gen[3280]),

			.O(gen[3338]),
			.E(gen[3340]),

			.SO(gen[3398]),
			.S(gen[3399]),
			.SE(gen[3400]),

			.SELF(gen[3339]),
			.cell_state(gen[3339])
		); 

/******************* CELL 3340 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3340 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3279]),
			.N(gen[3280]),
			.NE(gen[3281]),

			.O(gen[3339]),
			.E(gen[3341]),

			.SO(gen[3399]),
			.S(gen[3400]),
			.SE(gen[3401]),

			.SELF(gen[3340]),
			.cell_state(gen[3340])
		); 

/******************* CELL 3341 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3341 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3280]),
			.N(gen[3281]),
			.NE(gen[3282]),

			.O(gen[3340]),
			.E(gen[3342]),

			.SO(gen[3400]),
			.S(gen[3401]),
			.SE(gen[3402]),

			.SELF(gen[3341]),
			.cell_state(gen[3341])
		); 

/******************* CELL 3342 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3342 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3281]),
			.N(gen[3282]),
			.NE(gen[3283]),

			.O(gen[3341]),
			.E(gen[3343]),

			.SO(gen[3401]),
			.S(gen[3402]),
			.SE(gen[3403]),

			.SELF(gen[3342]),
			.cell_state(gen[3342])
		); 

/******************* CELL 3343 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3343 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3282]),
			.N(gen[3283]),
			.NE(gen[3284]),

			.O(gen[3342]),
			.E(gen[3344]),

			.SO(gen[3402]),
			.S(gen[3403]),
			.SE(gen[3404]),

			.SELF(gen[3343]),
			.cell_state(gen[3343])
		); 

/******************* CELL 3344 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3344 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3283]),
			.N(gen[3284]),
			.NE(gen[3285]),

			.O(gen[3343]),
			.E(gen[3345]),

			.SO(gen[3403]),
			.S(gen[3404]),
			.SE(gen[3405]),

			.SELF(gen[3344]),
			.cell_state(gen[3344])
		); 

/******************* CELL 3345 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3345 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3284]),
			.N(gen[3285]),
			.NE(gen[3286]),

			.O(gen[3344]),
			.E(gen[3346]),

			.SO(gen[3404]),
			.S(gen[3405]),
			.SE(gen[3406]),

			.SELF(gen[3345]),
			.cell_state(gen[3345])
		); 

/******************* CELL 3346 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3346 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3285]),
			.N(gen[3286]),
			.NE(gen[3287]),

			.O(gen[3345]),
			.E(gen[3347]),

			.SO(gen[3405]),
			.S(gen[3406]),
			.SE(gen[3407]),

			.SELF(gen[3346]),
			.cell_state(gen[3346])
		); 

/******************* CELL 3347 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3347 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3286]),
			.N(gen[3287]),
			.NE(gen[3288]),

			.O(gen[3346]),
			.E(gen[3348]),

			.SO(gen[3406]),
			.S(gen[3407]),
			.SE(gen[3408]),

			.SELF(gen[3347]),
			.cell_state(gen[3347])
		); 

/******************* CELL 3348 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3348 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3287]),
			.N(gen[3288]),
			.NE(gen[3289]),

			.O(gen[3347]),
			.E(gen[3349]),

			.SO(gen[3407]),
			.S(gen[3408]),
			.SE(gen[3409]),

			.SELF(gen[3348]),
			.cell_state(gen[3348])
		); 

/******************* CELL 3349 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3349 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3288]),
			.N(gen[3289]),
			.NE(gen[3290]),

			.O(gen[3348]),
			.E(gen[3350]),

			.SO(gen[3408]),
			.S(gen[3409]),
			.SE(gen[3410]),

			.SELF(gen[3349]),
			.cell_state(gen[3349])
		); 

/******************* CELL 3350 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3350 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3289]),
			.N(gen[3290]),
			.NE(gen[3291]),

			.O(gen[3349]),
			.E(gen[3351]),

			.SO(gen[3409]),
			.S(gen[3410]),
			.SE(gen[3411]),

			.SELF(gen[3350]),
			.cell_state(gen[3350])
		); 

/******************* CELL 3351 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3351 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3290]),
			.N(gen[3291]),
			.NE(gen[3292]),

			.O(gen[3350]),
			.E(gen[3352]),

			.SO(gen[3410]),
			.S(gen[3411]),
			.SE(gen[3412]),

			.SELF(gen[3351]),
			.cell_state(gen[3351])
		); 

/******************* CELL 3352 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3352 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3291]),
			.N(gen[3292]),
			.NE(gen[3293]),

			.O(gen[3351]),
			.E(gen[3353]),

			.SO(gen[3411]),
			.S(gen[3412]),
			.SE(gen[3413]),

			.SELF(gen[3352]),
			.cell_state(gen[3352])
		); 

/******************* CELL 3353 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3353 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3292]),
			.N(gen[3293]),
			.NE(gen[3294]),

			.O(gen[3352]),
			.E(gen[3354]),

			.SO(gen[3412]),
			.S(gen[3413]),
			.SE(gen[3414]),

			.SELF(gen[3353]),
			.cell_state(gen[3353])
		); 

/******************* CELL 3354 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3354 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3293]),
			.N(gen[3294]),
			.NE(gen[3295]),

			.O(gen[3353]),
			.E(gen[3355]),

			.SO(gen[3413]),
			.S(gen[3414]),
			.SE(gen[3415]),

			.SELF(gen[3354]),
			.cell_state(gen[3354])
		); 

/******************* CELL 3355 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3355 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3294]),
			.N(gen[3295]),
			.NE(gen[3296]),

			.O(gen[3354]),
			.E(gen[3356]),

			.SO(gen[3414]),
			.S(gen[3415]),
			.SE(gen[3416]),

			.SELF(gen[3355]),
			.cell_state(gen[3355])
		); 

/******************* CELL 3356 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3356 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3295]),
			.N(gen[3296]),
			.NE(gen[3297]),

			.O(gen[3355]),
			.E(gen[3357]),

			.SO(gen[3415]),
			.S(gen[3416]),
			.SE(gen[3417]),

			.SELF(gen[3356]),
			.cell_state(gen[3356])
		); 

/******************* CELL 3357 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3357 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3296]),
			.N(gen[3297]),
			.NE(gen[3298]),

			.O(gen[3356]),
			.E(gen[3358]),

			.SO(gen[3416]),
			.S(gen[3417]),
			.SE(gen[3418]),

			.SELF(gen[3357]),
			.cell_state(gen[3357])
		); 

/******************* CELL 3358 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3358 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3297]),
			.N(gen[3298]),
			.NE(gen[3299]),

			.O(gen[3357]),
			.E(gen[3359]),

			.SO(gen[3417]),
			.S(gen[3418]),
			.SE(gen[3419]),

			.SELF(gen[3358]),
			.cell_state(gen[3358])
		); 

/******************* CELL 3359 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3359 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3298]),
			.N(gen[3299]),
			.NE(gen[3298]),

			.O(gen[3358]),
			.E(gen[3358]),

			.SO(gen[3418]),
			.S(gen[3419]),
			.SE(gen[3418]),

			.SELF(gen[3359]),
			.cell_state(gen[3359])
		); 

/******************* CELL 3360 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3360 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3301]),
			.N(gen[3300]),
			.NE(gen[3301]),

			.O(gen[3361]),
			.E(gen[3361]),

			.SO(gen[3421]),
			.S(gen[3420]),
			.SE(gen[3421]),

			.SELF(gen[3360]),
			.cell_state(gen[3360])
		); 

/******************* CELL 3361 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3361 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3300]),
			.N(gen[3301]),
			.NE(gen[3302]),

			.O(gen[3360]),
			.E(gen[3362]),

			.SO(gen[3420]),
			.S(gen[3421]),
			.SE(gen[3422]),

			.SELF(gen[3361]),
			.cell_state(gen[3361])
		); 

/******************* CELL 3362 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3362 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3301]),
			.N(gen[3302]),
			.NE(gen[3303]),

			.O(gen[3361]),
			.E(gen[3363]),

			.SO(gen[3421]),
			.S(gen[3422]),
			.SE(gen[3423]),

			.SELF(gen[3362]),
			.cell_state(gen[3362])
		); 

/******************* CELL 3363 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3363 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3302]),
			.N(gen[3303]),
			.NE(gen[3304]),

			.O(gen[3362]),
			.E(gen[3364]),

			.SO(gen[3422]),
			.S(gen[3423]),
			.SE(gen[3424]),

			.SELF(gen[3363]),
			.cell_state(gen[3363])
		); 

/******************* CELL 3364 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3364 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3303]),
			.N(gen[3304]),
			.NE(gen[3305]),

			.O(gen[3363]),
			.E(gen[3365]),

			.SO(gen[3423]),
			.S(gen[3424]),
			.SE(gen[3425]),

			.SELF(gen[3364]),
			.cell_state(gen[3364])
		); 

/******************* CELL 3365 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3365 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3304]),
			.N(gen[3305]),
			.NE(gen[3306]),

			.O(gen[3364]),
			.E(gen[3366]),

			.SO(gen[3424]),
			.S(gen[3425]),
			.SE(gen[3426]),

			.SELF(gen[3365]),
			.cell_state(gen[3365])
		); 

/******************* CELL 3366 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3366 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3305]),
			.N(gen[3306]),
			.NE(gen[3307]),

			.O(gen[3365]),
			.E(gen[3367]),

			.SO(gen[3425]),
			.S(gen[3426]),
			.SE(gen[3427]),

			.SELF(gen[3366]),
			.cell_state(gen[3366])
		); 

/******************* CELL 3367 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3367 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3306]),
			.N(gen[3307]),
			.NE(gen[3308]),

			.O(gen[3366]),
			.E(gen[3368]),

			.SO(gen[3426]),
			.S(gen[3427]),
			.SE(gen[3428]),

			.SELF(gen[3367]),
			.cell_state(gen[3367])
		); 

/******************* CELL 3368 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3368 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3307]),
			.N(gen[3308]),
			.NE(gen[3309]),

			.O(gen[3367]),
			.E(gen[3369]),

			.SO(gen[3427]),
			.S(gen[3428]),
			.SE(gen[3429]),

			.SELF(gen[3368]),
			.cell_state(gen[3368])
		); 

/******************* CELL 3369 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3369 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3308]),
			.N(gen[3309]),
			.NE(gen[3310]),

			.O(gen[3368]),
			.E(gen[3370]),

			.SO(gen[3428]),
			.S(gen[3429]),
			.SE(gen[3430]),

			.SELF(gen[3369]),
			.cell_state(gen[3369])
		); 

/******************* CELL 3370 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3370 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3309]),
			.N(gen[3310]),
			.NE(gen[3311]),

			.O(gen[3369]),
			.E(gen[3371]),

			.SO(gen[3429]),
			.S(gen[3430]),
			.SE(gen[3431]),

			.SELF(gen[3370]),
			.cell_state(gen[3370])
		); 

/******************* CELL 3371 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3371 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3310]),
			.N(gen[3311]),
			.NE(gen[3312]),

			.O(gen[3370]),
			.E(gen[3372]),

			.SO(gen[3430]),
			.S(gen[3431]),
			.SE(gen[3432]),

			.SELF(gen[3371]),
			.cell_state(gen[3371])
		); 

/******************* CELL 3372 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3372 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3311]),
			.N(gen[3312]),
			.NE(gen[3313]),

			.O(gen[3371]),
			.E(gen[3373]),

			.SO(gen[3431]),
			.S(gen[3432]),
			.SE(gen[3433]),

			.SELF(gen[3372]),
			.cell_state(gen[3372])
		); 

/******************* CELL 3373 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3373 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3312]),
			.N(gen[3313]),
			.NE(gen[3314]),

			.O(gen[3372]),
			.E(gen[3374]),

			.SO(gen[3432]),
			.S(gen[3433]),
			.SE(gen[3434]),

			.SELF(gen[3373]),
			.cell_state(gen[3373])
		); 

/******************* CELL 3374 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3374 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3313]),
			.N(gen[3314]),
			.NE(gen[3315]),

			.O(gen[3373]),
			.E(gen[3375]),

			.SO(gen[3433]),
			.S(gen[3434]),
			.SE(gen[3435]),

			.SELF(gen[3374]),
			.cell_state(gen[3374])
		); 

/******************* CELL 3375 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3375 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3314]),
			.N(gen[3315]),
			.NE(gen[3316]),

			.O(gen[3374]),
			.E(gen[3376]),

			.SO(gen[3434]),
			.S(gen[3435]),
			.SE(gen[3436]),

			.SELF(gen[3375]),
			.cell_state(gen[3375])
		); 

/******************* CELL 3376 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3376 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3315]),
			.N(gen[3316]),
			.NE(gen[3317]),

			.O(gen[3375]),
			.E(gen[3377]),

			.SO(gen[3435]),
			.S(gen[3436]),
			.SE(gen[3437]),

			.SELF(gen[3376]),
			.cell_state(gen[3376])
		); 

/******************* CELL 3377 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3377 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3316]),
			.N(gen[3317]),
			.NE(gen[3318]),

			.O(gen[3376]),
			.E(gen[3378]),

			.SO(gen[3436]),
			.S(gen[3437]),
			.SE(gen[3438]),

			.SELF(gen[3377]),
			.cell_state(gen[3377])
		); 

/******************* CELL 3378 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3378 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3317]),
			.N(gen[3318]),
			.NE(gen[3319]),

			.O(gen[3377]),
			.E(gen[3379]),

			.SO(gen[3437]),
			.S(gen[3438]),
			.SE(gen[3439]),

			.SELF(gen[3378]),
			.cell_state(gen[3378])
		); 

/******************* CELL 3379 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3379 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3318]),
			.N(gen[3319]),
			.NE(gen[3320]),

			.O(gen[3378]),
			.E(gen[3380]),

			.SO(gen[3438]),
			.S(gen[3439]),
			.SE(gen[3440]),

			.SELF(gen[3379]),
			.cell_state(gen[3379])
		); 

/******************* CELL 3380 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3380 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3319]),
			.N(gen[3320]),
			.NE(gen[3321]),

			.O(gen[3379]),
			.E(gen[3381]),

			.SO(gen[3439]),
			.S(gen[3440]),
			.SE(gen[3441]),

			.SELF(gen[3380]),
			.cell_state(gen[3380])
		); 

/******************* CELL 3381 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3381 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3320]),
			.N(gen[3321]),
			.NE(gen[3322]),

			.O(gen[3380]),
			.E(gen[3382]),

			.SO(gen[3440]),
			.S(gen[3441]),
			.SE(gen[3442]),

			.SELF(gen[3381]),
			.cell_state(gen[3381])
		); 

/******************* CELL 3382 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3382 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3321]),
			.N(gen[3322]),
			.NE(gen[3323]),

			.O(gen[3381]),
			.E(gen[3383]),

			.SO(gen[3441]),
			.S(gen[3442]),
			.SE(gen[3443]),

			.SELF(gen[3382]),
			.cell_state(gen[3382])
		); 

/******************* CELL 3383 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3383 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3322]),
			.N(gen[3323]),
			.NE(gen[3324]),

			.O(gen[3382]),
			.E(gen[3384]),

			.SO(gen[3442]),
			.S(gen[3443]),
			.SE(gen[3444]),

			.SELF(gen[3383]),
			.cell_state(gen[3383])
		); 

/******************* CELL 3384 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3384 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3323]),
			.N(gen[3324]),
			.NE(gen[3325]),

			.O(gen[3383]),
			.E(gen[3385]),

			.SO(gen[3443]),
			.S(gen[3444]),
			.SE(gen[3445]),

			.SELF(gen[3384]),
			.cell_state(gen[3384])
		); 

/******************* CELL 3385 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3385 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3324]),
			.N(gen[3325]),
			.NE(gen[3326]),

			.O(gen[3384]),
			.E(gen[3386]),

			.SO(gen[3444]),
			.S(gen[3445]),
			.SE(gen[3446]),

			.SELF(gen[3385]),
			.cell_state(gen[3385])
		); 

/******************* CELL 3386 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3386 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3325]),
			.N(gen[3326]),
			.NE(gen[3327]),

			.O(gen[3385]),
			.E(gen[3387]),

			.SO(gen[3445]),
			.S(gen[3446]),
			.SE(gen[3447]),

			.SELF(gen[3386]),
			.cell_state(gen[3386])
		); 

/******************* CELL 3387 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3387 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3326]),
			.N(gen[3327]),
			.NE(gen[3328]),

			.O(gen[3386]),
			.E(gen[3388]),

			.SO(gen[3446]),
			.S(gen[3447]),
			.SE(gen[3448]),

			.SELF(gen[3387]),
			.cell_state(gen[3387])
		); 

/******************* CELL 3388 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3388 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3327]),
			.N(gen[3328]),
			.NE(gen[3329]),

			.O(gen[3387]),
			.E(gen[3389]),

			.SO(gen[3447]),
			.S(gen[3448]),
			.SE(gen[3449]),

			.SELF(gen[3388]),
			.cell_state(gen[3388])
		); 

/******************* CELL 3389 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3389 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3328]),
			.N(gen[3329]),
			.NE(gen[3330]),

			.O(gen[3388]),
			.E(gen[3390]),

			.SO(gen[3448]),
			.S(gen[3449]),
			.SE(gen[3450]),

			.SELF(gen[3389]),
			.cell_state(gen[3389])
		); 

/******************* CELL 3390 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3390 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3329]),
			.N(gen[3330]),
			.NE(gen[3331]),

			.O(gen[3389]),
			.E(gen[3391]),

			.SO(gen[3449]),
			.S(gen[3450]),
			.SE(gen[3451]),

			.SELF(gen[3390]),
			.cell_state(gen[3390])
		); 

/******************* CELL 3391 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3391 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3330]),
			.N(gen[3331]),
			.NE(gen[3332]),

			.O(gen[3390]),
			.E(gen[3392]),

			.SO(gen[3450]),
			.S(gen[3451]),
			.SE(gen[3452]),

			.SELF(gen[3391]),
			.cell_state(gen[3391])
		); 

/******************* CELL 3392 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3392 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3331]),
			.N(gen[3332]),
			.NE(gen[3333]),

			.O(gen[3391]),
			.E(gen[3393]),

			.SO(gen[3451]),
			.S(gen[3452]),
			.SE(gen[3453]),

			.SELF(gen[3392]),
			.cell_state(gen[3392])
		); 

/******************* CELL 3393 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3393 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3332]),
			.N(gen[3333]),
			.NE(gen[3334]),

			.O(gen[3392]),
			.E(gen[3394]),

			.SO(gen[3452]),
			.S(gen[3453]),
			.SE(gen[3454]),

			.SELF(gen[3393]),
			.cell_state(gen[3393])
		); 

/******************* CELL 3394 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3394 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3333]),
			.N(gen[3334]),
			.NE(gen[3335]),

			.O(gen[3393]),
			.E(gen[3395]),

			.SO(gen[3453]),
			.S(gen[3454]),
			.SE(gen[3455]),

			.SELF(gen[3394]),
			.cell_state(gen[3394])
		); 

/******************* CELL 3395 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3395 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3334]),
			.N(gen[3335]),
			.NE(gen[3336]),

			.O(gen[3394]),
			.E(gen[3396]),

			.SO(gen[3454]),
			.S(gen[3455]),
			.SE(gen[3456]),

			.SELF(gen[3395]),
			.cell_state(gen[3395])
		); 

/******************* CELL 3396 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3396 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3335]),
			.N(gen[3336]),
			.NE(gen[3337]),

			.O(gen[3395]),
			.E(gen[3397]),

			.SO(gen[3455]),
			.S(gen[3456]),
			.SE(gen[3457]),

			.SELF(gen[3396]),
			.cell_state(gen[3396])
		); 

/******************* CELL 3397 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3397 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3336]),
			.N(gen[3337]),
			.NE(gen[3338]),

			.O(gen[3396]),
			.E(gen[3398]),

			.SO(gen[3456]),
			.S(gen[3457]),
			.SE(gen[3458]),

			.SELF(gen[3397]),
			.cell_state(gen[3397])
		); 

/******************* CELL 3398 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3398 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3337]),
			.N(gen[3338]),
			.NE(gen[3339]),

			.O(gen[3397]),
			.E(gen[3399]),

			.SO(gen[3457]),
			.S(gen[3458]),
			.SE(gen[3459]),

			.SELF(gen[3398]),
			.cell_state(gen[3398])
		); 

/******************* CELL 3399 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3399 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3338]),
			.N(gen[3339]),
			.NE(gen[3340]),

			.O(gen[3398]),
			.E(gen[3400]),

			.SO(gen[3458]),
			.S(gen[3459]),
			.SE(gen[3460]),

			.SELF(gen[3399]),
			.cell_state(gen[3399])
		); 

/******************* CELL 3400 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3400 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3339]),
			.N(gen[3340]),
			.NE(gen[3341]),

			.O(gen[3399]),
			.E(gen[3401]),

			.SO(gen[3459]),
			.S(gen[3460]),
			.SE(gen[3461]),

			.SELF(gen[3400]),
			.cell_state(gen[3400])
		); 

/******************* CELL 3401 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3401 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3340]),
			.N(gen[3341]),
			.NE(gen[3342]),

			.O(gen[3400]),
			.E(gen[3402]),

			.SO(gen[3460]),
			.S(gen[3461]),
			.SE(gen[3462]),

			.SELF(gen[3401]),
			.cell_state(gen[3401])
		); 

/******************* CELL 3402 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3402 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3341]),
			.N(gen[3342]),
			.NE(gen[3343]),

			.O(gen[3401]),
			.E(gen[3403]),

			.SO(gen[3461]),
			.S(gen[3462]),
			.SE(gen[3463]),

			.SELF(gen[3402]),
			.cell_state(gen[3402])
		); 

/******************* CELL 3403 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3403 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3342]),
			.N(gen[3343]),
			.NE(gen[3344]),

			.O(gen[3402]),
			.E(gen[3404]),

			.SO(gen[3462]),
			.S(gen[3463]),
			.SE(gen[3464]),

			.SELF(gen[3403]),
			.cell_state(gen[3403])
		); 

/******************* CELL 3404 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3404 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3343]),
			.N(gen[3344]),
			.NE(gen[3345]),

			.O(gen[3403]),
			.E(gen[3405]),

			.SO(gen[3463]),
			.S(gen[3464]),
			.SE(gen[3465]),

			.SELF(gen[3404]),
			.cell_state(gen[3404])
		); 

/******************* CELL 3405 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3405 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3344]),
			.N(gen[3345]),
			.NE(gen[3346]),

			.O(gen[3404]),
			.E(gen[3406]),

			.SO(gen[3464]),
			.S(gen[3465]),
			.SE(gen[3466]),

			.SELF(gen[3405]),
			.cell_state(gen[3405])
		); 

/******************* CELL 3406 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3406 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3345]),
			.N(gen[3346]),
			.NE(gen[3347]),

			.O(gen[3405]),
			.E(gen[3407]),

			.SO(gen[3465]),
			.S(gen[3466]),
			.SE(gen[3467]),

			.SELF(gen[3406]),
			.cell_state(gen[3406])
		); 

/******************* CELL 3407 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3407 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3346]),
			.N(gen[3347]),
			.NE(gen[3348]),

			.O(gen[3406]),
			.E(gen[3408]),

			.SO(gen[3466]),
			.S(gen[3467]),
			.SE(gen[3468]),

			.SELF(gen[3407]),
			.cell_state(gen[3407])
		); 

/******************* CELL 3408 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3408 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3347]),
			.N(gen[3348]),
			.NE(gen[3349]),

			.O(gen[3407]),
			.E(gen[3409]),

			.SO(gen[3467]),
			.S(gen[3468]),
			.SE(gen[3469]),

			.SELF(gen[3408]),
			.cell_state(gen[3408])
		); 

/******************* CELL 3409 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3409 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3348]),
			.N(gen[3349]),
			.NE(gen[3350]),

			.O(gen[3408]),
			.E(gen[3410]),

			.SO(gen[3468]),
			.S(gen[3469]),
			.SE(gen[3470]),

			.SELF(gen[3409]),
			.cell_state(gen[3409])
		); 

/******************* CELL 3410 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3410 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3349]),
			.N(gen[3350]),
			.NE(gen[3351]),

			.O(gen[3409]),
			.E(gen[3411]),

			.SO(gen[3469]),
			.S(gen[3470]),
			.SE(gen[3471]),

			.SELF(gen[3410]),
			.cell_state(gen[3410])
		); 

/******************* CELL 3411 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3411 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3350]),
			.N(gen[3351]),
			.NE(gen[3352]),

			.O(gen[3410]),
			.E(gen[3412]),

			.SO(gen[3470]),
			.S(gen[3471]),
			.SE(gen[3472]),

			.SELF(gen[3411]),
			.cell_state(gen[3411])
		); 

/******************* CELL 3412 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3412 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3351]),
			.N(gen[3352]),
			.NE(gen[3353]),

			.O(gen[3411]),
			.E(gen[3413]),

			.SO(gen[3471]),
			.S(gen[3472]),
			.SE(gen[3473]),

			.SELF(gen[3412]),
			.cell_state(gen[3412])
		); 

/******************* CELL 3413 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3413 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3352]),
			.N(gen[3353]),
			.NE(gen[3354]),

			.O(gen[3412]),
			.E(gen[3414]),

			.SO(gen[3472]),
			.S(gen[3473]),
			.SE(gen[3474]),

			.SELF(gen[3413]),
			.cell_state(gen[3413])
		); 

/******************* CELL 3414 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3414 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3353]),
			.N(gen[3354]),
			.NE(gen[3355]),

			.O(gen[3413]),
			.E(gen[3415]),

			.SO(gen[3473]),
			.S(gen[3474]),
			.SE(gen[3475]),

			.SELF(gen[3414]),
			.cell_state(gen[3414])
		); 

/******************* CELL 3415 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3415 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3354]),
			.N(gen[3355]),
			.NE(gen[3356]),

			.O(gen[3414]),
			.E(gen[3416]),

			.SO(gen[3474]),
			.S(gen[3475]),
			.SE(gen[3476]),

			.SELF(gen[3415]),
			.cell_state(gen[3415])
		); 

/******************* CELL 3416 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3416 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3355]),
			.N(gen[3356]),
			.NE(gen[3357]),

			.O(gen[3415]),
			.E(gen[3417]),

			.SO(gen[3475]),
			.S(gen[3476]),
			.SE(gen[3477]),

			.SELF(gen[3416]),
			.cell_state(gen[3416])
		); 

/******************* CELL 3417 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3417 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3356]),
			.N(gen[3357]),
			.NE(gen[3358]),

			.O(gen[3416]),
			.E(gen[3418]),

			.SO(gen[3476]),
			.S(gen[3477]),
			.SE(gen[3478]),

			.SELF(gen[3417]),
			.cell_state(gen[3417])
		); 

/******************* CELL 3418 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3418 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3357]),
			.N(gen[3358]),
			.NE(gen[3359]),

			.O(gen[3417]),
			.E(gen[3419]),

			.SO(gen[3477]),
			.S(gen[3478]),
			.SE(gen[3479]),

			.SELF(gen[3418]),
			.cell_state(gen[3418])
		); 

/******************* CELL 3419 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3419 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3358]),
			.N(gen[3359]),
			.NE(gen[3358]),

			.O(gen[3418]),
			.E(gen[3418]),

			.SO(gen[3478]),
			.S(gen[3479]),
			.SE(gen[3478]),

			.SELF(gen[3419]),
			.cell_state(gen[3419])
		); 

/******************* CELL 3420 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3420 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3361]),
			.N(gen[3360]),
			.NE(gen[3361]),

			.O(gen[3421]),
			.E(gen[3421]),

			.SO(gen[3481]),
			.S(gen[3480]),
			.SE(gen[3481]),

			.SELF(gen[3420]),
			.cell_state(gen[3420])
		); 

/******************* CELL 3421 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3421 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3360]),
			.N(gen[3361]),
			.NE(gen[3362]),

			.O(gen[3420]),
			.E(gen[3422]),

			.SO(gen[3480]),
			.S(gen[3481]),
			.SE(gen[3482]),

			.SELF(gen[3421]),
			.cell_state(gen[3421])
		); 

/******************* CELL 3422 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3422 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3361]),
			.N(gen[3362]),
			.NE(gen[3363]),

			.O(gen[3421]),
			.E(gen[3423]),

			.SO(gen[3481]),
			.S(gen[3482]),
			.SE(gen[3483]),

			.SELF(gen[3422]),
			.cell_state(gen[3422])
		); 

/******************* CELL 3423 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3423 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3362]),
			.N(gen[3363]),
			.NE(gen[3364]),

			.O(gen[3422]),
			.E(gen[3424]),

			.SO(gen[3482]),
			.S(gen[3483]),
			.SE(gen[3484]),

			.SELF(gen[3423]),
			.cell_state(gen[3423])
		); 

/******************* CELL 3424 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3424 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3363]),
			.N(gen[3364]),
			.NE(gen[3365]),

			.O(gen[3423]),
			.E(gen[3425]),

			.SO(gen[3483]),
			.S(gen[3484]),
			.SE(gen[3485]),

			.SELF(gen[3424]),
			.cell_state(gen[3424])
		); 

/******************* CELL 3425 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3425 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3364]),
			.N(gen[3365]),
			.NE(gen[3366]),

			.O(gen[3424]),
			.E(gen[3426]),

			.SO(gen[3484]),
			.S(gen[3485]),
			.SE(gen[3486]),

			.SELF(gen[3425]),
			.cell_state(gen[3425])
		); 

/******************* CELL 3426 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3426 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3365]),
			.N(gen[3366]),
			.NE(gen[3367]),

			.O(gen[3425]),
			.E(gen[3427]),

			.SO(gen[3485]),
			.S(gen[3486]),
			.SE(gen[3487]),

			.SELF(gen[3426]),
			.cell_state(gen[3426])
		); 

/******************* CELL 3427 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3427 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3366]),
			.N(gen[3367]),
			.NE(gen[3368]),

			.O(gen[3426]),
			.E(gen[3428]),

			.SO(gen[3486]),
			.S(gen[3487]),
			.SE(gen[3488]),

			.SELF(gen[3427]),
			.cell_state(gen[3427])
		); 

/******************* CELL 3428 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3428 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3367]),
			.N(gen[3368]),
			.NE(gen[3369]),

			.O(gen[3427]),
			.E(gen[3429]),

			.SO(gen[3487]),
			.S(gen[3488]),
			.SE(gen[3489]),

			.SELF(gen[3428]),
			.cell_state(gen[3428])
		); 

/******************* CELL 3429 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3429 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3368]),
			.N(gen[3369]),
			.NE(gen[3370]),

			.O(gen[3428]),
			.E(gen[3430]),

			.SO(gen[3488]),
			.S(gen[3489]),
			.SE(gen[3490]),

			.SELF(gen[3429]),
			.cell_state(gen[3429])
		); 

/******************* CELL 3430 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3430 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3369]),
			.N(gen[3370]),
			.NE(gen[3371]),

			.O(gen[3429]),
			.E(gen[3431]),

			.SO(gen[3489]),
			.S(gen[3490]),
			.SE(gen[3491]),

			.SELF(gen[3430]),
			.cell_state(gen[3430])
		); 

/******************* CELL 3431 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3431 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3370]),
			.N(gen[3371]),
			.NE(gen[3372]),

			.O(gen[3430]),
			.E(gen[3432]),

			.SO(gen[3490]),
			.S(gen[3491]),
			.SE(gen[3492]),

			.SELF(gen[3431]),
			.cell_state(gen[3431])
		); 

/******************* CELL 3432 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3432 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3371]),
			.N(gen[3372]),
			.NE(gen[3373]),

			.O(gen[3431]),
			.E(gen[3433]),

			.SO(gen[3491]),
			.S(gen[3492]),
			.SE(gen[3493]),

			.SELF(gen[3432]),
			.cell_state(gen[3432])
		); 

/******************* CELL 3433 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3433 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3372]),
			.N(gen[3373]),
			.NE(gen[3374]),

			.O(gen[3432]),
			.E(gen[3434]),

			.SO(gen[3492]),
			.S(gen[3493]),
			.SE(gen[3494]),

			.SELF(gen[3433]),
			.cell_state(gen[3433])
		); 

/******************* CELL 3434 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3434 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3373]),
			.N(gen[3374]),
			.NE(gen[3375]),

			.O(gen[3433]),
			.E(gen[3435]),

			.SO(gen[3493]),
			.S(gen[3494]),
			.SE(gen[3495]),

			.SELF(gen[3434]),
			.cell_state(gen[3434])
		); 

/******************* CELL 3435 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3435 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3374]),
			.N(gen[3375]),
			.NE(gen[3376]),

			.O(gen[3434]),
			.E(gen[3436]),

			.SO(gen[3494]),
			.S(gen[3495]),
			.SE(gen[3496]),

			.SELF(gen[3435]),
			.cell_state(gen[3435])
		); 

/******************* CELL 3436 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3436 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3375]),
			.N(gen[3376]),
			.NE(gen[3377]),

			.O(gen[3435]),
			.E(gen[3437]),

			.SO(gen[3495]),
			.S(gen[3496]),
			.SE(gen[3497]),

			.SELF(gen[3436]),
			.cell_state(gen[3436])
		); 

/******************* CELL 3437 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3437 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3376]),
			.N(gen[3377]),
			.NE(gen[3378]),

			.O(gen[3436]),
			.E(gen[3438]),

			.SO(gen[3496]),
			.S(gen[3497]),
			.SE(gen[3498]),

			.SELF(gen[3437]),
			.cell_state(gen[3437])
		); 

/******************* CELL 3438 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3438 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3377]),
			.N(gen[3378]),
			.NE(gen[3379]),

			.O(gen[3437]),
			.E(gen[3439]),

			.SO(gen[3497]),
			.S(gen[3498]),
			.SE(gen[3499]),

			.SELF(gen[3438]),
			.cell_state(gen[3438])
		); 

/******************* CELL 3439 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3439 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3378]),
			.N(gen[3379]),
			.NE(gen[3380]),

			.O(gen[3438]),
			.E(gen[3440]),

			.SO(gen[3498]),
			.S(gen[3499]),
			.SE(gen[3500]),

			.SELF(gen[3439]),
			.cell_state(gen[3439])
		); 

/******************* CELL 3440 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3440 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3379]),
			.N(gen[3380]),
			.NE(gen[3381]),

			.O(gen[3439]),
			.E(gen[3441]),

			.SO(gen[3499]),
			.S(gen[3500]),
			.SE(gen[3501]),

			.SELF(gen[3440]),
			.cell_state(gen[3440])
		); 

/******************* CELL 3441 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3441 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3380]),
			.N(gen[3381]),
			.NE(gen[3382]),

			.O(gen[3440]),
			.E(gen[3442]),

			.SO(gen[3500]),
			.S(gen[3501]),
			.SE(gen[3502]),

			.SELF(gen[3441]),
			.cell_state(gen[3441])
		); 

/******************* CELL 3442 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3442 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3381]),
			.N(gen[3382]),
			.NE(gen[3383]),

			.O(gen[3441]),
			.E(gen[3443]),

			.SO(gen[3501]),
			.S(gen[3502]),
			.SE(gen[3503]),

			.SELF(gen[3442]),
			.cell_state(gen[3442])
		); 

/******************* CELL 3443 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3443 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3382]),
			.N(gen[3383]),
			.NE(gen[3384]),

			.O(gen[3442]),
			.E(gen[3444]),

			.SO(gen[3502]),
			.S(gen[3503]),
			.SE(gen[3504]),

			.SELF(gen[3443]),
			.cell_state(gen[3443])
		); 

/******************* CELL 3444 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3444 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3383]),
			.N(gen[3384]),
			.NE(gen[3385]),

			.O(gen[3443]),
			.E(gen[3445]),

			.SO(gen[3503]),
			.S(gen[3504]),
			.SE(gen[3505]),

			.SELF(gen[3444]),
			.cell_state(gen[3444])
		); 

/******************* CELL 3445 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3445 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3384]),
			.N(gen[3385]),
			.NE(gen[3386]),

			.O(gen[3444]),
			.E(gen[3446]),

			.SO(gen[3504]),
			.S(gen[3505]),
			.SE(gen[3506]),

			.SELF(gen[3445]),
			.cell_state(gen[3445])
		); 

/******************* CELL 3446 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3446 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3385]),
			.N(gen[3386]),
			.NE(gen[3387]),

			.O(gen[3445]),
			.E(gen[3447]),

			.SO(gen[3505]),
			.S(gen[3506]),
			.SE(gen[3507]),

			.SELF(gen[3446]),
			.cell_state(gen[3446])
		); 

/******************* CELL 3447 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3447 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3386]),
			.N(gen[3387]),
			.NE(gen[3388]),

			.O(gen[3446]),
			.E(gen[3448]),

			.SO(gen[3506]),
			.S(gen[3507]),
			.SE(gen[3508]),

			.SELF(gen[3447]),
			.cell_state(gen[3447])
		); 

/******************* CELL 3448 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3448 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3387]),
			.N(gen[3388]),
			.NE(gen[3389]),

			.O(gen[3447]),
			.E(gen[3449]),

			.SO(gen[3507]),
			.S(gen[3508]),
			.SE(gen[3509]),

			.SELF(gen[3448]),
			.cell_state(gen[3448])
		); 

/******************* CELL 3449 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3449 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3388]),
			.N(gen[3389]),
			.NE(gen[3390]),

			.O(gen[3448]),
			.E(gen[3450]),

			.SO(gen[3508]),
			.S(gen[3509]),
			.SE(gen[3510]),

			.SELF(gen[3449]),
			.cell_state(gen[3449])
		); 

/******************* CELL 3450 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3450 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3389]),
			.N(gen[3390]),
			.NE(gen[3391]),

			.O(gen[3449]),
			.E(gen[3451]),

			.SO(gen[3509]),
			.S(gen[3510]),
			.SE(gen[3511]),

			.SELF(gen[3450]),
			.cell_state(gen[3450])
		); 

/******************* CELL 3451 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3451 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3390]),
			.N(gen[3391]),
			.NE(gen[3392]),

			.O(gen[3450]),
			.E(gen[3452]),

			.SO(gen[3510]),
			.S(gen[3511]),
			.SE(gen[3512]),

			.SELF(gen[3451]),
			.cell_state(gen[3451])
		); 

/******************* CELL 3452 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3452 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3391]),
			.N(gen[3392]),
			.NE(gen[3393]),

			.O(gen[3451]),
			.E(gen[3453]),

			.SO(gen[3511]),
			.S(gen[3512]),
			.SE(gen[3513]),

			.SELF(gen[3452]),
			.cell_state(gen[3452])
		); 

/******************* CELL 3453 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3453 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3392]),
			.N(gen[3393]),
			.NE(gen[3394]),

			.O(gen[3452]),
			.E(gen[3454]),

			.SO(gen[3512]),
			.S(gen[3513]),
			.SE(gen[3514]),

			.SELF(gen[3453]),
			.cell_state(gen[3453])
		); 

/******************* CELL 3454 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3454 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3393]),
			.N(gen[3394]),
			.NE(gen[3395]),

			.O(gen[3453]),
			.E(gen[3455]),

			.SO(gen[3513]),
			.S(gen[3514]),
			.SE(gen[3515]),

			.SELF(gen[3454]),
			.cell_state(gen[3454])
		); 

/******************* CELL 3455 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3455 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3394]),
			.N(gen[3395]),
			.NE(gen[3396]),

			.O(gen[3454]),
			.E(gen[3456]),

			.SO(gen[3514]),
			.S(gen[3515]),
			.SE(gen[3516]),

			.SELF(gen[3455]),
			.cell_state(gen[3455])
		); 

/******************* CELL 3456 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3456 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3395]),
			.N(gen[3396]),
			.NE(gen[3397]),

			.O(gen[3455]),
			.E(gen[3457]),

			.SO(gen[3515]),
			.S(gen[3516]),
			.SE(gen[3517]),

			.SELF(gen[3456]),
			.cell_state(gen[3456])
		); 

/******************* CELL 3457 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3457 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3396]),
			.N(gen[3397]),
			.NE(gen[3398]),

			.O(gen[3456]),
			.E(gen[3458]),

			.SO(gen[3516]),
			.S(gen[3517]),
			.SE(gen[3518]),

			.SELF(gen[3457]),
			.cell_state(gen[3457])
		); 

/******************* CELL 3458 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3458 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3397]),
			.N(gen[3398]),
			.NE(gen[3399]),

			.O(gen[3457]),
			.E(gen[3459]),

			.SO(gen[3517]),
			.S(gen[3518]),
			.SE(gen[3519]),

			.SELF(gen[3458]),
			.cell_state(gen[3458])
		); 

/******************* CELL 3459 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3459 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3398]),
			.N(gen[3399]),
			.NE(gen[3400]),

			.O(gen[3458]),
			.E(gen[3460]),

			.SO(gen[3518]),
			.S(gen[3519]),
			.SE(gen[3520]),

			.SELF(gen[3459]),
			.cell_state(gen[3459])
		); 

/******************* CELL 3460 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3460 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3399]),
			.N(gen[3400]),
			.NE(gen[3401]),

			.O(gen[3459]),
			.E(gen[3461]),

			.SO(gen[3519]),
			.S(gen[3520]),
			.SE(gen[3521]),

			.SELF(gen[3460]),
			.cell_state(gen[3460])
		); 

/******************* CELL 3461 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3461 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3400]),
			.N(gen[3401]),
			.NE(gen[3402]),

			.O(gen[3460]),
			.E(gen[3462]),

			.SO(gen[3520]),
			.S(gen[3521]),
			.SE(gen[3522]),

			.SELF(gen[3461]),
			.cell_state(gen[3461])
		); 

/******************* CELL 3462 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3462 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3401]),
			.N(gen[3402]),
			.NE(gen[3403]),

			.O(gen[3461]),
			.E(gen[3463]),

			.SO(gen[3521]),
			.S(gen[3522]),
			.SE(gen[3523]),

			.SELF(gen[3462]),
			.cell_state(gen[3462])
		); 

/******************* CELL 3463 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3463 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3402]),
			.N(gen[3403]),
			.NE(gen[3404]),

			.O(gen[3462]),
			.E(gen[3464]),

			.SO(gen[3522]),
			.S(gen[3523]),
			.SE(gen[3524]),

			.SELF(gen[3463]),
			.cell_state(gen[3463])
		); 

/******************* CELL 3464 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3464 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3403]),
			.N(gen[3404]),
			.NE(gen[3405]),

			.O(gen[3463]),
			.E(gen[3465]),

			.SO(gen[3523]),
			.S(gen[3524]),
			.SE(gen[3525]),

			.SELF(gen[3464]),
			.cell_state(gen[3464])
		); 

/******************* CELL 3465 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3465 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3404]),
			.N(gen[3405]),
			.NE(gen[3406]),

			.O(gen[3464]),
			.E(gen[3466]),

			.SO(gen[3524]),
			.S(gen[3525]),
			.SE(gen[3526]),

			.SELF(gen[3465]),
			.cell_state(gen[3465])
		); 

/******************* CELL 3466 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3466 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3405]),
			.N(gen[3406]),
			.NE(gen[3407]),

			.O(gen[3465]),
			.E(gen[3467]),

			.SO(gen[3525]),
			.S(gen[3526]),
			.SE(gen[3527]),

			.SELF(gen[3466]),
			.cell_state(gen[3466])
		); 

/******************* CELL 3467 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3467 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3406]),
			.N(gen[3407]),
			.NE(gen[3408]),

			.O(gen[3466]),
			.E(gen[3468]),

			.SO(gen[3526]),
			.S(gen[3527]),
			.SE(gen[3528]),

			.SELF(gen[3467]),
			.cell_state(gen[3467])
		); 

/******************* CELL 3468 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3468 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3407]),
			.N(gen[3408]),
			.NE(gen[3409]),

			.O(gen[3467]),
			.E(gen[3469]),

			.SO(gen[3527]),
			.S(gen[3528]),
			.SE(gen[3529]),

			.SELF(gen[3468]),
			.cell_state(gen[3468])
		); 

/******************* CELL 3469 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3469 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3408]),
			.N(gen[3409]),
			.NE(gen[3410]),

			.O(gen[3468]),
			.E(gen[3470]),

			.SO(gen[3528]),
			.S(gen[3529]),
			.SE(gen[3530]),

			.SELF(gen[3469]),
			.cell_state(gen[3469])
		); 

/******************* CELL 3470 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3470 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3409]),
			.N(gen[3410]),
			.NE(gen[3411]),

			.O(gen[3469]),
			.E(gen[3471]),

			.SO(gen[3529]),
			.S(gen[3530]),
			.SE(gen[3531]),

			.SELF(gen[3470]),
			.cell_state(gen[3470])
		); 

/******************* CELL 3471 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3471 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3410]),
			.N(gen[3411]),
			.NE(gen[3412]),

			.O(gen[3470]),
			.E(gen[3472]),

			.SO(gen[3530]),
			.S(gen[3531]),
			.SE(gen[3532]),

			.SELF(gen[3471]),
			.cell_state(gen[3471])
		); 

/******************* CELL 3472 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3472 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3411]),
			.N(gen[3412]),
			.NE(gen[3413]),

			.O(gen[3471]),
			.E(gen[3473]),

			.SO(gen[3531]),
			.S(gen[3532]),
			.SE(gen[3533]),

			.SELF(gen[3472]),
			.cell_state(gen[3472])
		); 

/******************* CELL 3473 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3473 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3412]),
			.N(gen[3413]),
			.NE(gen[3414]),

			.O(gen[3472]),
			.E(gen[3474]),

			.SO(gen[3532]),
			.S(gen[3533]),
			.SE(gen[3534]),

			.SELF(gen[3473]),
			.cell_state(gen[3473])
		); 

/******************* CELL 3474 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3474 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3413]),
			.N(gen[3414]),
			.NE(gen[3415]),

			.O(gen[3473]),
			.E(gen[3475]),

			.SO(gen[3533]),
			.S(gen[3534]),
			.SE(gen[3535]),

			.SELF(gen[3474]),
			.cell_state(gen[3474])
		); 

/******************* CELL 3475 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3475 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3414]),
			.N(gen[3415]),
			.NE(gen[3416]),

			.O(gen[3474]),
			.E(gen[3476]),

			.SO(gen[3534]),
			.S(gen[3535]),
			.SE(gen[3536]),

			.SELF(gen[3475]),
			.cell_state(gen[3475])
		); 

/******************* CELL 3476 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3476 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3415]),
			.N(gen[3416]),
			.NE(gen[3417]),

			.O(gen[3475]),
			.E(gen[3477]),

			.SO(gen[3535]),
			.S(gen[3536]),
			.SE(gen[3537]),

			.SELF(gen[3476]),
			.cell_state(gen[3476])
		); 

/******************* CELL 3477 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3477 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3416]),
			.N(gen[3417]),
			.NE(gen[3418]),

			.O(gen[3476]),
			.E(gen[3478]),

			.SO(gen[3536]),
			.S(gen[3537]),
			.SE(gen[3538]),

			.SELF(gen[3477]),
			.cell_state(gen[3477])
		); 

/******************* CELL 3478 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3478 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3417]),
			.N(gen[3418]),
			.NE(gen[3419]),

			.O(gen[3477]),
			.E(gen[3479]),

			.SO(gen[3537]),
			.S(gen[3538]),
			.SE(gen[3539]),

			.SELF(gen[3478]),
			.cell_state(gen[3478])
		); 

/******************* CELL 3479 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3479 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3418]),
			.N(gen[3419]),
			.NE(gen[3418]),

			.O(gen[3478]),
			.E(gen[3478]),

			.SO(gen[3538]),
			.S(gen[3539]),
			.SE(gen[3538]),

			.SELF(gen[3479]),
			.cell_state(gen[3479])
		); 

/******************* CELL 3480 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3480 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3421]),
			.N(gen[3420]),
			.NE(gen[3421]),

			.O(gen[3481]),
			.E(gen[3481]),

			.SO(gen[3541]),
			.S(gen[3540]),
			.SE(gen[3541]),

			.SELF(gen[3480]),
			.cell_state(gen[3480])
		); 

/******************* CELL 3481 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3481 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3420]),
			.N(gen[3421]),
			.NE(gen[3422]),

			.O(gen[3480]),
			.E(gen[3482]),

			.SO(gen[3540]),
			.S(gen[3541]),
			.SE(gen[3542]),

			.SELF(gen[3481]),
			.cell_state(gen[3481])
		); 

/******************* CELL 3482 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3482 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3421]),
			.N(gen[3422]),
			.NE(gen[3423]),

			.O(gen[3481]),
			.E(gen[3483]),

			.SO(gen[3541]),
			.S(gen[3542]),
			.SE(gen[3543]),

			.SELF(gen[3482]),
			.cell_state(gen[3482])
		); 

/******************* CELL 3483 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3483 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3422]),
			.N(gen[3423]),
			.NE(gen[3424]),

			.O(gen[3482]),
			.E(gen[3484]),

			.SO(gen[3542]),
			.S(gen[3543]),
			.SE(gen[3544]),

			.SELF(gen[3483]),
			.cell_state(gen[3483])
		); 

/******************* CELL 3484 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3484 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3423]),
			.N(gen[3424]),
			.NE(gen[3425]),

			.O(gen[3483]),
			.E(gen[3485]),

			.SO(gen[3543]),
			.S(gen[3544]),
			.SE(gen[3545]),

			.SELF(gen[3484]),
			.cell_state(gen[3484])
		); 

/******************* CELL 3485 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3485 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3424]),
			.N(gen[3425]),
			.NE(gen[3426]),

			.O(gen[3484]),
			.E(gen[3486]),

			.SO(gen[3544]),
			.S(gen[3545]),
			.SE(gen[3546]),

			.SELF(gen[3485]),
			.cell_state(gen[3485])
		); 

/******************* CELL 3486 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3486 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3425]),
			.N(gen[3426]),
			.NE(gen[3427]),

			.O(gen[3485]),
			.E(gen[3487]),

			.SO(gen[3545]),
			.S(gen[3546]),
			.SE(gen[3547]),

			.SELF(gen[3486]),
			.cell_state(gen[3486])
		); 

/******************* CELL 3487 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3487 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3426]),
			.N(gen[3427]),
			.NE(gen[3428]),

			.O(gen[3486]),
			.E(gen[3488]),

			.SO(gen[3546]),
			.S(gen[3547]),
			.SE(gen[3548]),

			.SELF(gen[3487]),
			.cell_state(gen[3487])
		); 

/******************* CELL 3488 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3488 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3427]),
			.N(gen[3428]),
			.NE(gen[3429]),

			.O(gen[3487]),
			.E(gen[3489]),

			.SO(gen[3547]),
			.S(gen[3548]),
			.SE(gen[3549]),

			.SELF(gen[3488]),
			.cell_state(gen[3488])
		); 

/******************* CELL 3489 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3489 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3428]),
			.N(gen[3429]),
			.NE(gen[3430]),

			.O(gen[3488]),
			.E(gen[3490]),

			.SO(gen[3548]),
			.S(gen[3549]),
			.SE(gen[3550]),

			.SELF(gen[3489]),
			.cell_state(gen[3489])
		); 

/******************* CELL 3490 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3490 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3429]),
			.N(gen[3430]),
			.NE(gen[3431]),

			.O(gen[3489]),
			.E(gen[3491]),

			.SO(gen[3549]),
			.S(gen[3550]),
			.SE(gen[3551]),

			.SELF(gen[3490]),
			.cell_state(gen[3490])
		); 

/******************* CELL 3491 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3491 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3430]),
			.N(gen[3431]),
			.NE(gen[3432]),

			.O(gen[3490]),
			.E(gen[3492]),

			.SO(gen[3550]),
			.S(gen[3551]),
			.SE(gen[3552]),

			.SELF(gen[3491]),
			.cell_state(gen[3491])
		); 

/******************* CELL 3492 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3492 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3431]),
			.N(gen[3432]),
			.NE(gen[3433]),

			.O(gen[3491]),
			.E(gen[3493]),

			.SO(gen[3551]),
			.S(gen[3552]),
			.SE(gen[3553]),

			.SELF(gen[3492]),
			.cell_state(gen[3492])
		); 

/******************* CELL 3493 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3493 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3432]),
			.N(gen[3433]),
			.NE(gen[3434]),

			.O(gen[3492]),
			.E(gen[3494]),

			.SO(gen[3552]),
			.S(gen[3553]),
			.SE(gen[3554]),

			.SELF(gen[3493]),
			.cell_state(gen[3493])
		); 

/******************* CELL 3494 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3494 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3433]),
			.N(gen[3434]),
			.NE(gen[3435]),

			.O(gen[3493]),
			.E(gen[3495]),

			.SO(gen[3553]),
			.S(gen[3554]),
			.SE(gen[3555]),

			.SELF(gen[3494]),
			.cell_state(gen[3494])
		); 

/******************* CELL 3495 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3495 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3434]),
			.N(gen[3435]),
			.NE(gen[3436]),

			.O(gen[3494]),
			.E(gen[3496]),

			.SO(gen[3554]),
			.S(gen[3555]),
			.SE(gen[3556]),

			.SELF(gen[3495]),
			.cell_state(gen[3495])
		); 

/******************* CELL 3496 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3496 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3435]),
			.N(gen[3436]),
			.NE(gen[3437]),

			.O(gen[3495]),
			.E(gen[3497]),

			.SO(gen[3555]),
			.S(gen[3556]),
			.SE(gen[3557]),

			.SELF(gen[3496]),
			.cell_state(gen[3496])
		); 

/******************* CELL 3497 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3497 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3436]),
			.N(gen[3437]),
			.NE(gen[3438]),

			.O(gen[3496]),
			.E(gen[3498]),

			.SO(gen[3556]),
			.S(gen[3557]),
			.SE(gen[3558]),

			.SELF(gen[3497]),
			.cell_state(gen[3497])
		); 

/******************* CELL 3498 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3498 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3437]),
			.N(gen[3438]),
			.NE(gen[3439]),

			.O(gen[3497]),
			.E(gen[3499]),

			.SO(gen[3557]),
			.S(gen[3558]),
			.SE(gen[3559]),

			.SELF(gen[3498]),
			.cell_state(gen[3498])
		); 

/******************* CELL 3499 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3499 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3438]),
			.N(gen[3439]),
			.NE(gen[3440]),

			.O(gen[3498]),
			.E(gen[3500]),

			.SO(gen[3558]),
			.S(gen[3559]),
			.SE(gen[3560]),

			.SELF(gen[3499]),
			.cell_state(gen[3499])
		); 

/******************* CELL 3500 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3500 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3439]),
			.N(gen[3440]),
			.NE(gen[3441]),

			.O(gen[3499]),
			.E(gen[3501]),

			.SO(gen[3559]),
			.S(gen[3560]),
			.SE(gen[3561]),

			.SELF(gen[3500]),
			.cell_state(gen[3500])
		); 

/******************* CELL 3501 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3501 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3440]),
			.N(gen[3441]),
			.NE(gen[3442]),

			.O(gen[3500]),
			.E(gen[3502]),

			.SO(gen[3560]),
			.S(gen[3561]),
			.SE(gen[3562]),

			.SELF(gen[3501]),
			.cell_state(gen[3501])
		); 

/******************* CELL 3502 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3502 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3441]),
			.N(gen[3442]),
			.NE(gen[3443]),

			.O(gen[3501]),
			.E(gen[3503]),

			.SO(gen[3561]),
			.S(gen[3562]),
			.SE(gen[3563]),

			.SELF(gen[3502]),
			.cell_state(gen[3502])
		); 

/******************* CELL 3503 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3503 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3442]),
			.N(gen[3443]),
			.NE(gen[3444]),

			.O(gen[3502]),
			.E(gen[3504]),

			.SO(gen[3562]),
			.S(gen[3563]),
			.SE(gen[3564]),

			.SELF(gen[3503]),
			.cell_state(gen[3503])
		); 

/******************* CELL 3504 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3504 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3443]),
			.N(gen[3444]),
			.NE(gen[3445]),

			.O(gen[3503]),
			.E(gen[3505]),

			.SO(gen[3563]),
			.S(gen[3564]),
			.SE(gen[3565]),

			.SELF(gen[3504]),
			.cell_state(gen[3504])
		); 

/******************* CELL 3505 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3505 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3444]),
			.N(gen[3445]),
			.NE(gen[3446]),

			.O(gen[3504]),
			.E(gen[3506]),

			.SO(gen[3564]),
			.S(gen[3565]),
			.SE(gen[3566]),

			.SELF(gen[3505]),
			.cell_state(gen[3505])
		); 

/******************* CELL 3506 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3506 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3445]),
			.N(gen[3446]),
			.NE(gen[3447]),

			.O(gen[3505]),
			.E(gen[3507]),

			.SO(gen[3565]),
			.S(gen[3566]),
			.SE(gen[3567]),

			.SELF(gen[3506]),
			.cell_state(gen[3506])
		); 

/******************* CELL 3507 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3507 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3446]),
			.N(gen[3447]),
			.NE(gen[3448]),

			.O(gen[3506]),
			.E(gen[3508]),

			.SO(gen[3566]),
			.S(gen[3567]),
			.SE(gen[3568]),

			.SELF(gen[3507]),
			.cell_state(gen[3507])
		); 

/******************* CELL 3508 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3508 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3447]),
			.N(gen[3448]),
			.NE(gen[3449]),

			.O(gen[3507]),
			.E(gen[3509]),

			.SO(gen[3567]),
			.S(gen[3568]),
			.SE(gen[3569]),

			.SELF(gen[3508]),
			.cell_state(gen[3508])
		); 

/******************* CELL 3509 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3509 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3448]),
			.N(gen[3449]),
			.NE(gen[3450]),

			.O(gen[3508]),
			.E(gen[3510]),

			.SO(gen[3568]),
			.S(gen[3569]),
			.SE(gen[3570]),

			.SELF(gen[3509]),
			.cell_state(gen[3509])
		); 

/******************* CELL 3510 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3510 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3449]),
			.N(gen[3450]),
			.NE(gen[3451]),

			.O(gen[3509]),
			.E(gen[3511]),

			.SO(gen[3569]),
			.S(gen[3570]),
			.SE(gen[3571]),

			.SELF(gen[3510]),
			.cell_state(gen[3510])
		); 

/******************* CELL 3511 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3511 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3450]),
			.N(gen[3451]),
			.NE(gen[3452]),

			.O(gen[3510]),
			.E(gen[3512]),

			.SO(gen[3570]),
			.S(gen[3571]),
			.SE(gen[3572]),

			.SELF(gen[3511]),
			.cell_state(gen[3511])
		); 

/******************* CELL 3512 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3512 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3451]),
			.N(gen[3452]),
			.NE(gen[3453]),

			.O(gen[3511]),
			.E(gen[3513]),

			.SO(gen[3571]),
			.S(gen[3572]),
			.SE(gen[3573]),

			.SELF(gen[3512]),
			.cell_state(gen[3512])
		); 

/******************* CELL 3513 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3513 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3452]),
			.N(gen[3453]),
			.NE(gen[3454]),

			.O(gen[3512]),
			.E(gen[3514]),

			.SO(gen[3572]),
			.S(gen[3573]),
			.SE(gen[3574]),

			.SELF(gen[3513]),
			.cell_state(gen[3513])
		); 

/******************* CELL 3514 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3514 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3453]),
			.N(gen[3454]),
			.NE(gen[3455]),

			.O(gen[3513]),
			.E(gen[3515]),

			.SO(gen[3573]),
			.S(gen[3574]),
			.SE(gen[3575]),

			.SELF(gen[3514]),
			.cell_state(gen[3514])
		); 

/******************* CELL 3515 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3515 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3454]),
			.N(gen[3455]),
			.NE(gen[3456]),

			.O(gen[3514]),
			.E(gen[3516]),

			.SO(gen[3574]),
			.S(gen[3575]),
			.SE(gen[3576]),

			.SELF(gen[3515]),
			.cell_state(gen[3515])
		); 

/******************* CELL 3516 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3516 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3455]),
			.N(gen[3456]),
			.NE(gen[3457]),

			.O(gen[3515]),
			.E(gen[3517]),

			.SO(gen[3575]),
			.S(gen[3576]),
			.SE(gen[3577]),

			.SELF(gen[3516]),
			.cell_state(gen[3516])
		); 

/******************* CELL 3517 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3517 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3456]),
			.N(gen[3457]),
			.NE(gen[3458]),

			.O(gen[3516]),
			.E(gen[3518]),

			.SO(gen[3576]),
			.S(gen[3577]),
			.SE(gen[3578]),

			.SELF(gen[3517]),
			.cell_state(gen[3517])
		); 

/******************* CELL 3518 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3518 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3457]),
			.N(gen[3458]),
			.NE(gen[3459]),

			.O(gen[3517]),
			.E(gen[3519]),

			.SO(gen[3577]),
			.S(gen[3578]),
			.SE(gen[3579]),

			.SELF(gen[3518]),
			.cell_state(gen[3518])
		); 

/******************* CELL 3519 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3519 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3458]),
			.N(gen[3459]),
			.NE(gen[3460]),

			.O(gen[3518]),
			.E(gen[3520]),

			.SO(gen[3578]),
			.S(gen[3579]),
			.SE(gen[3580]),

			.SELF(gen[3519]),
			.cell_state(gen[3519])
		); 

/******************* CELL 3520 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3520 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3459]),
			.N(gen[3460]),
			.NE(gen[3461]),

			.O(gen[3519]),
			.E(gen[3521]),

			.SO(gen[3579]),
			.S(gen[3580]),
			.SE(gen[3581]),

			.SELF(gen[3520]),
			.cell_state(gen[3520])
		); 

/******************* CELL 3521 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3521 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3460]),
			.N(gen[3461]),
			.NE(gen[3462]),

			.O(gen[3520]),
			.E(gen[3522]),

			.SO(gen[3580]),
			.S(gen[3581]),
			.SE(gen[3582]),

			.SELF(gen[3521]),
			.cell_state(gen[3521])
		); 

/******************* CELL 3522 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3522 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3461]),
			.N(gen[3462]),
			.NE(gen[3463]),

			.O(gen[3521]),
			.E(gen[3523]),

			.SO(gen[3581]),
			.S(gen[3582]),
			.SE(gen[3583]),

			.SELF(gen[3522]),
			.cell_state(gen[3522])
		); 

/******************* CELL 3523 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3523 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3462]),
			.N(gen[3463]),
			.NE(gen[3464]),

			.O(gen[3522]),
			.E(gen[3524]),

			.SO(gen[3582]),
			.S(gen[3583]),
			.SE(gen[3584]),

			.SELF(gen[3523]),
			.cell_state(gen[3523])
		); 

/******************* CELL 3524 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3524 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3463]),
			.N(gen[3464]),
			.NE(gen[3465]),

			.O(gen[3523]),
			.E(gen[3525]),

			.SO(gen[3583]),
			.S(gen[3584]),
			.SE(gen[3585]),

			.SELF(gen[3524]),
			.cell_state(gen[3524])
		); 

/******************* CELL 3525 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3525 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3464]),
			.N(gen[3465]),
			.NE(gen[3466]),

			.O(gen[3524]),
			.E(gen[3526]),

			.SO(gen[3584]),
			.S(gen[3585]),
			.SE(gen[3586]),

			.SELF(gen[3525]),
			.cell_state(gen[3525])
		); 

/******************* CELL 3526 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3526 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3465]),
			.N(gen[3466]),
			.NE(gen[3467]),

			.O(gen[3525]),
			.E(gen[3527]),

			.SO(gen[3585]),
			.S(gen[3586]),
			.SE(gen[3587]),

			.SELF(gen[3526]),
			.cell_state(gen[3526])
		); 

/******************* CELL 3527 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3527 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3466]),
			.N(gen[3467]),
			.NE(gen[3468]),

			.O(gen[3526]),
			.E(gen[3528]),

			.SO(gen[3586]),
			.S(gen[3587]),
			.SE(gen[3588]),

			.SELF(gen[3527]),
			.cell_state(gen[3527])
		); 

/******************* CELL 3528 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3528 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3467]),
			.N(gen[3468]),
			.NE(gen[3469]),

			.O(gen[3527]),
			.E(gen[3529]),

			.SO(gen[3587]),
			.S(gen[3588]),
			.SE(gen[3589]),

			.SELF(gen[3528]),
			.cell_state(gen[3528])
		); 

/******************* CELL 3529 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3529 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3468]),
			.N(gen[3469]),
			.NE(gen[3470]),

			.O(gen[3528]),
			.E(gen[3530]),

			.SO(gen[3588]),
			.S(gen[3589]),
			.SE(gen[3590]),

			.SELF(gen[3529]),
			.cell_state(gen[3529])
		); 

/******************* CELL 3530 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3530 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3469]),
			.N(gen[3470]),
			.NE(gen[3471]),

			.O(gen[3529]),
			.E(gen[3531]),

			.SO(gen[3589]),
			.S(gen[3590]),
			.SE(gen[3591]),

			.SELF(gen[3530]),
			.cell_state(gen[3530])
		); 

/******************* CELL 3531 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3531 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3470]),
			.N(gen[3471]),
			.NE(gen[3472]),

			.O(gen[3530]),
			.E(gen[3532]),

			.SO(gen[3590]),
			.S(gen[3591]),
			.SE(gen[3592]),

			.SELF(gen[3531]),
			.cell_state(gen[3531])
		); 

/******************* CELL 3532 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3532 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3471]),
			.N(gen[3472]),
			.NE(gen[3473]),

			.O(gen[3531]),
			.E(gen[3533]),

			.SO(gen[3591]),
			.S(gen[3592]),
			.SE(gen[3593]),

			.SELF(gen[3532]),
			.cell_state(gen[3532])
		); 

/******************* CELL 3533 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3533 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3472]),
			.N(gen[3473]),
			.NE(gen[3474]),

			.O(gen[3532]),
			.E(gen[3534]),

			.SO(gen[3592]),
			.S(gen[3593]),
			.SE(gen[3594]),

			.SELF(gen[3533]),
			.cell_state(gen[3533])
		); 

/******************* CELL 3534 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3534 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3473]),
			.N(gen[3474]),
			.NE(gen[3475]),

			.O(gen[3533]),
			.E(gen[3535]),

			.SO(gen[3593]),
			.S(gen[3594]),
			.SE(gen[3595]),

			.SELF(gen[3534]),
			.cell_state(gen[3534])
		); 

/******************* CELL 3535 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3535 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3474]),
			.N(gen[3475]),
			.NE(gen[3476]),

			.O(gen[3534]),
			.E(gen[3536]),

			.SO(gen[3594]),
			.S(gen[3595]),
			.SE(gen[3596]),

			.SELF(gen[3535]),
			.cell_state(gen[3535])
		); 

/******************* CELL 3536 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3536 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3475]),
			.N(gen[3476]),
			.NE(gen[3477]),

			.O(gen[3535]),
			.E(gen[3537]),

			.SO(gen[3595]),
			.S(gen[3596]),
			.SE(gen[3597]),

			.SELF(gen[3536]),
			.cell_state(gen[3536])
		); 

/******************* CELL 3537 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3537 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3476]),
			.N(gen[3477]),
			.NE(gen[3478]),

			.O(gen[3536]),
			.E(gen[3538]),

			.SO(gen[3596]),
			.S(gen[3597]),
			.SE(gen[3598]),

			.SELF(gen[3537]),
			.cell_state(gen[3537])
		); 

/******************* CELL 3538 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3538 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3477]),
			.N(gen[3478]),
			.NE(gen[3479]),

			.O(gen[3537]),
			.E(gen[3539]),

			.SO(gen[3597]),
			.S(gen[3598]),
			.SE(gen[3599]),

			.SELF(gen[3538]),
			.cell_state(gen[3538])
		); 

/******************* CELL 3539 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(0))

		cell3539 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3478]),
			.N(gen[3479]),
			.NE(gen[3478]),

			.O(gen[3538]),
			.E(gen[3538]),

			.SO(gen[3598]),
			.S(gen[3599]),
			.SE(gen[3598]),

			.SELF(gen[3539]),
			.cell_state(gen[3539])
		); 

/******************* CELL 3540 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3540 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3481]),
			.N(gen[3480]),
			.NE(gen[3481]),

			.O(gen[3541]),
			.E(gen[3541]),

			.SO(gen[3481]),
			.S(gen[3480]),
			.SE(gen[3481]),

			.SELF(gen[3540]),
			.cell_state(gen[3540])
		); 

/******************* CELL 3541 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3541 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3480]),
			.N(gen[3481]),
			.NE(gen[3482]),

			.O(gen[3540]),
			.E(gen[3542]),

			.SO(gen[3480]),
			.S(gen[3481]),
			.SE(gen[3482]),

			.SELF(gen[3541]),
			.cell_state(gen[3541])
		); 

/******************* CELL 3542 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3542 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3481]),
			.N(gen[3482]),
			.NE(gen[3483]),

			.O(gen[3541]),
			.E(gen[3543]),

			.SO(gen[3481]),
			.S(gen[3482]),
			.SE(gen[3483]),

			.SELF(gen[3542]),
			.cell_state(gen[3542])
		); 

/******************* CELL 3543 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3543 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3482]),
			.N(gen[3483]),
			.NE(gen[3484]),

			.O(gen[3542]),
			.E(gen[3544]),

			.SO(gen[3482]),
			.S(gen[3483]),
			.SE(gen[3484]),

			.SELF(gen[3543]),
			.cell_state(gen[3543])
		); 

/******************* CELL 3544 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3544 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3483]),
			.N(gen[3484]),
			.NE(gen[3485]),

			.O(gen[3543]),
			.E(gen[3545]),

			.SO(gen[3483]),
			.S(gen[3484]),
			.SE(gen[3485]),

			.SELF(gen[3544]),
			.cell_state(gen[3544])
		); 

/******************* CELL 3545 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3545 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3484]),
			.N(gen[3485]),
			.NE(gen[3486]),

			.O(gen[3544]),
			.E(gen[3546]),

			.SO(gen[3484]),
			.S(gen[3485]),
			.SE(gen[3486]),

			.SELF(gen[3545]),
			.cell_state(gen[3545])
		); 

/******************* CELL 3546 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3546 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3485]),
			.N(gen[3486]),
			.NE(gen[3487]),

			.O(gen[3545]),
			.E(gen[3547]),

			.SO(gen[3485]),
			.S(gen[3486]),
			.SE(gen[3487]),

			.SELF(gen[3546]),
			.cell_state(gen[3546])
		); 

/******************* CELL 3547 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3547 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3486]),
			.N(gen[3487]),
			.NE(gen[3488]),

			.O(gen[3546]),
			.E(gen[3548]),

			.SO(gen[3486]),
			.S(gen[3487]),
			.SE(gen[3488]),

			.SELF(gen[3547]),
			.cell_state(gen[3547])
		); 

/******************* CELL 3548 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3548 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3487]),
			.N(gen[3488]),
			.NE(gen[3489]),

			.O(gen[3547]),
			.E(gen[3549]),

			.SO(gen[3487]),
			.S(gen[3488]),
			.SE(gen[3489]),

			.SELF(gen[3548]),
			.cell_state(gen[3548])
		); 

/******************* CELL 3549 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3549 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3488]),
			.N(gen[3489]),
			.NE(gen[3490]),

			.O(gen[3548]),
			.E(gen[3550]),

			.SO(gen[3488]),
			.S(gen[3489]),
			.SE(gen[3490]),

			.SELF(gen[3549]),
			.cell_state(gen[3549])
		); 

/******************* CELL 3550 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3550 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3489]),
			.N(gen[3490]),
			.NE(gen[3491]),

			.O(gen[3549]),
			.E(gen[3551]),

			.SO(gen[3489]),
			.S(gen[3490]),
			.SE(gen[3491]),

			.SELF(gen[3550]),
			.cell_state(gen[3550])
		); 

/******************* CELL 3551 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3551 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3490]),
			.N(gen[3491]),
			.NE(gen[3492]),

			.O(gen[3550]),
			.E(gen[3552]),

			.SO(gen[3490]),
			.S(gen[3491]),
			.SE(gen[3492]),

			.SELF(gen[3551]),
			.cell_state(gen[3551])
		); 

/******************* CELL 3552 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3552 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3491]),
			.N(gen[3492]),
			.NE(gen[3493]),

			.O(gen[3551]),
			.E(gen[3553]),

			.SO(gen[3491]),
			.S(gen[3492]),
			.SE(gen[3493]),

			.SELF(gen[3552]),
			.cell_state(gen[3552])
		); 

/******************* CELL 3553 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3553 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3492]),
			.N(gen[3493]),
			.NE(gen[3494]),

			.O(gen[3552]),
			.E(gen[3554]),

			.SO(gen[3492]),
			.S(gen[3493]),
			.SE(gen[3494]),

			.SELF(gen[3553]),
			.cell_state(gen[3553])
		); 

/******************* CELL 3554 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3554 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3493]),
			.N(gen[3494]),
			.NE(gen[3495]),

			.O(gen[3553]),
			.E(gen[3555]),

			.SO(gen[3493]),
			.S(gen[3494]),
			.SE(gen[3495]),

			.SELF(gen[3554]),
			.cell_state(gen[3554])
		); 

/******************* CELL 3555 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3555 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3494]),
			.N(gen[3495]),
			.NE(gen[3496]),

			.O(gen[3554]),
			.E(gen[3556]),

			.SO(gen[3494]),
			.S(gen[3495]),
			.SE(gen[3496]),

			.SELF(gen[3555]),
			.cell_state(gen[3555])
		); 

/******************* CELL 3556 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3556 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3495]),
			.N(gen[3496]),
			.NE(gen[3497]),

			.O(gen[3555]),
			.E(gen[3557]),

			.SO(gen[3495]),
			.S(gen[3496]),
			.SE(gen[3497]),

			.SELF(gen[3556]),
			.cell_state(gen[3556])
		); 

/******************* CELL 3557 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3557 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3496]),
			.N(gen[3497]),
			.NE(gen[3498]),

			.O(gen[3556]),
			.E(gen[3558]),

			.SO(gen[3496]),
			.S(gen[3497]),
			.SE(gen[3498]),

			.SELF(gen[3557]),
			.cell_state(gen[3557])
		); 

/******************* CELL 3558 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3558 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3497]),
			.N(gen[3498]),
			.NE(gen[3499]),

			.O(gen[3557]),
			.E(gen[3559]),

			.SO(gen[3497]),
			.S(gen[3498]),
			.SE(gen[3499]),

			.SELF(gen[3558]),
			.cell_state(gen[3558])
		); 

/******************* CELL 3559 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3559 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3498]),
			.N(gen[3499]),
			.NE(gen[3500]),

			.O(gen[3558]),
			.E(gen[3560]),

			.SO(gen[3498]),
			.S(gen[3499]),
			.SE(gen[3500]),

			.SELF(gen[3559]),
			.cell_state(gen[3559])
		); 

/******************* CELL 3560 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3560 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3499]),
			.N(gen[3500]),
			.NE(gen[3501]),

			.O(gen[3559]),
			.E(gen[3561]),

			.SO(gen[3499]),
			.S(gen[3500]),
			.SE(gen[3501]),

			.SELF(gen[3560]),
			.cell_state(gen[3560])
		); 

/******************* CELL 3561 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3561 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3500]),
			.N(gen[3501]),
			.NE(gen[3502]),

			.O(gen[3560]),
			.E(gen[3562]),

			.SO(gen[3500]),
			.S(gen[3501]),
			.SE(gen[3502]),

			.SELF(gen[3561]),
			.cell_state(gen[3561])
		); 

/******************* CELL 3562 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3562 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3501]),
			.N(gen[3502]),
			.NE(gen[3503]),

			.O(gen[3561]),
			.E(gen[3563]),

			.SO(gen[3501]),
			.S(gen[3502]),
			.SE(gen[3503]),

			.SELF(gen[3562]),
			.cell_state(gen[3562])
		); 

/******************* CELL 3563 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3563 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3502]),
			.N(gen[3503]),
			.NE(gen[3504]),

			.O(gen[3562]),
			.E(gen[3564]),

			.SO(gen[3502]),
			.S(gen[3503]),
			.SE(gen[3504]),

			.SELF(gen[3563]),
			.cell_state(gen[3563])
		); 

/******************* CELL 3564 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3564 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3503]),
			.N(gen[3504]),
			.NE(gen[3505]),

			.O(gen[3563]),
			.E(gen[3565]),

			.SO(gen[3503]),
			.S(gen[3504]),
			.SE(gen[3505]),

			.SELF(gen[3564]),
			.cell_state(gen[3564])
		); 

/******************* CELL 3565 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3565 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3504]),
			.N(gen[3505]),
			.NE(gen[3506]),

			.O(gen[3564]),
			.E(gen[3566]),

			.SO(gen[3504]),
			.S(gen[3505]),
			.SE(gen[3506]),

			.SELF(gen[3565]),
			.cell_state(gen[3565])
		); 

/******************* CELL 3566 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3566 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3505]),
			.N(gen[3506]),
			.NE(gen[3507]),

			.O(gen[3565]),
			.E(gen[3567]),

			.SO(gen[3505]),
			.S(gen[3506]),
			.SE(gen[3507]),

			.SELF(gen[3566]),
			.cell_state(gen[3566])
		); 

/******************* CELL 3567 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3567 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3506]),
			.N(gen[3507]),
			.NE(gen[3508]),

			.O(gen[3566]),
			.E(gen[3568]),

			.SO(gen[3506]),
			.S(gen[3507]),
			.SE(gen[3508]),

			.SELF(gen[3567]),
			.cell_state(gen[3567])
		); 

/******************* CELL 3568 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3568 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3507]),
			.N(gen[3508]),
			.NE(gen[3509]),

			.O(gen[3567]),
			.E(gen[3569]),

			.SO(gen[3507]),
			.S(gen[3508]),
			.SE(gen[3509]),

			.SELF(gen[3568]),
			.cell_state(gen[3568])
		); 

/******************* CELL 3569 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3569 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3508]),
			.N(gen[3509]),
			.NE(gen[3510]),

			.O(gen[3568]),
			.E(gen[3570]),

			.SO(gen[3508]),
			.S(gen[3509]),
			.SE(gen[3510]),

			.SELF(gen[3569]),
			.cell_state(gen[3569])
		); 

/******************* CELL 3570 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3570 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3509]),
			.N(gen[3510]),
			.NE(gen[3511]),

			.O(gen[3569]),
			.E(gen[3571]),

			.SO(gen[3509]),
			.S(gen[3510]),
			.SE(gen[3511]),

			.SELF(gen[3570]),
			.cell_state(gen[3570])
		); 

/******************* CELL 3571 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3571 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3510]),
			.N(gen[3511]),
			.NE(gen[3512]),

			.O(gen[3570]),
			.E(gen[3572]),

			.SO(gen[3510]),
			.S(gen[3511]),
			.SE(gen[3512]),

			.SELF(gen[3571]),
			.cell_state(gen[3571])
		); 

/******************* CELL 3572 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3572 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3511]),
			.N(gen[3512]),
			.NE(gen[3513]),

			.O(gen[3571]),
			.E(gen[3573]),

			.SO(gen[3511]),
			.S(gen[3512]),
			.SE(gen[3513]),

			.SELF(gen[3572]),
			.cell_state(gen[3572])
		); 

/******************* CELL 3573 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3573 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3512]),
			.N(gen[3513]),
			.NE(gen[3514]),

			.O(gen[3572]),
			.E(gen[3574]),

			.SO(gen[3512]),
			.S(gen[3513]),
			.SE(gen[3514]),

			.SELF(gen[3573]),
			.cell_state(gen[3573])
		); 

/******************* CELL 3574 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3574 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3513]),
			.N(gen[3514]),
			.NE(gen[3515]),

			.O(gen[3573]),
			.E(gen[3575]),

			.SO(gen[3513]),
			.S(gen[3514]),
			.SE(gen[3515]),

			.SELF(gen[3574]),
			.cell_state(gen[3574])
		); 

/******************* CELL 3575 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3575 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3514]),
			.N(gen[3515]),
			.NE(gen[3516]),

			.O(gen[3574]),
			.E(gen[3576]),

			.SO(gen[3514]),
			.S(gen[3515]),
			.SE(gen[3516]),

			.SELF(gen[3575]),
			.cell_state(gen[3575])
		); 

/******************* CELL 3576 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3576 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3515]),
			.N(gen[3516]),
			.NE(gen[3517]),

			.O(gen[3575]),
			.E(gen[3577]),

			.SO(gen[3515]),
			.S(gen[3516]),
			.SE(gen[3517]),

			.SELF(gen[3576]),
			.cell_state(gen[3576])
		); 

/******************* CELL 3577 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3577 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3516]),
			.N(gen[3517]),
			.NE(gen[3518]),

			.O(gen[3576]),
			.E(gen[3578]),

			.SO(gen[3516]),
			.S(gen[3517]),
			.SE(gen[3518]),

			.SELF(gen[3577]),
			.cell_state(gen[3577])
		); 

/******************* CELL 3578 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3578 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3517]),
			.N(gen[3518]),
			.NE(gen[3519]),

			.O(gen[3577]),
			.E(gen[3579]),

			.SO(gen[3517]),
			.S(gen[3518]),
			.SE(gen[3519]),

			.SELF(gen[3578]),
			.cell_state(gen[3578])
		); 

/******************* CELL 3579 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3579 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3518]),
			.N(gen[3519]),
			.NE(gen[3520]),

			.O(gen[3578]),
			.E(gen[3580]),

			.SO(gen[3518]),
			.S(gen[3519]),
			.SE(gen[3520]),

			.SELF(gen[3579]),
			.cell_state(gen[3579])
		); 

/******************* CELL 3580 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3580 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3519]),
			.N(gen[3520]),
			.NE(gen[3521]),

			.O(gen[3579]),
			.E(gen[3581]),

			.SO(gen[3519]),
			.S(gen[3520]),
			.SE(gen[3521]),

			.SELF(gen[3580]),
			.cell_state(gen[3580])
		); 

/******************* CELL 3581 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3581 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3520]),
			.N(gen[3521]),
			.NE(gen[3522]),

			.O(gen[3580]),
			.E(gen[3582]),

			.SO(gen[3520]),
			.S(gen[3521]),
			.SE(gen[3522]),

			.SELF(gen[3581]),
			.cell_state(gen[3581])
		); 

/******************* CELL 3582 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3582 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3521]),
			.N(gen[3522]),
			.NE(gen[3523]),

			.O(gen[3581]),
			.E(gen[3583]),

			.SO(gen[3521]),
			.S(gen[3522]),
			.SE(gen[3523]),

			.SELF(gen[3582]),
			.cell_state(gen[3582])
		); 

/******************* CELL 3583 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3583 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3522]),
			.N(gen[3523]),
			.NE(gen[3524]),

			.O(gen[3582]),
			.E(gen[3584]),

			.SO(gen[3522]),
			.S(gen[3523]),
			.SE(gen[3524]),

			.SELF(gen[3583]),
			.cell_state(gen[3583])
		); 

/******************* CELL 3584 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3584 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3523]),
			.N(gen[3524]),
			.NE(gen[3525]),

			.O(gen[3583]),
			.E(gen[3585]),

			.SO(gen[3523]),
			.S(gen[3524]),
			.SE(gen[3525]),

			.SELF(gen[3584]),
			.cell_state(gen[3584])
		); 

/******************* CELL 3585 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3585 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3524]),
			.N(gen[3525]),
			.NE(gen[3526]),

			.O(gen[3584]),
			.E(gen[3586]),

			.SO(gen[3524]),
			.S(gen[3525]),
			.SE(gen[3526]),

			.SELF(gen[3585]),
			.cell_state(gen[3585])
		); 

/******************* CELL 3586 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3586 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3525]),
			.N(gen[3526]),
			.NE(gen[3527]),

			.O(gen[3585]),
			.E(gen[3587]),

			.SO(gen[3525]),
			.S(gen[3526]),
			.SE(gen[3527]),

			.SELF(gen[3586]),
			.cell_state(gen[3586])
		); 

/******************* CELL 3587 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3587 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3526]),
			.N(gen[3527]),
			.NE(gen[3528]),

			.O(gen[3586]),
			.E(gen[3588]),

			.SO(gen[3526]),
			.S(gen[3527]),
			.SE(gen[3528]),

			.SELF(gen[3587]),
			.cell_state(gen[3587])
		); 

/******************* CELL 3588 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3588 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3527]),
			.N(gen[3528]),
			.NE(gen[3529]),

			.O(gen[3587]),
			.E(gen[3589]),

			.SO(gen[3527]),
			.S(gen[3528]),
			.SE(gen[3529]),

			.SELF(gen[3588]),
			.cell_state(gen[3588])
		); 

/******************* CELL 3589 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3589 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3528]),
			.N(gen[3529]),
			.NE(gen[3530]),

			.O(gen[3588]),
			.E(gen[3590]),

			.SO(gen[3528]),
			.S(gen[3529]),
			.SE(gen[3530]),

			.SELF(gen[3589]),
			.cell_state(gen[3589])
		); 

/******************* CELL 3590 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3590 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3529]),
			.N(gen[3530]),
			.NE(gen[3531]),

			.O(gen[3589]),
			.E(gen[3591]),

			.SO(gen[3529]),
			.S(gen[3530]),
			.SE(gen[3531]),

			.SELF(gen[3590]),
			.cell_state(gen[3590])
		); 

/******************* CELL 3591 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3591 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3530]),
			.N(gen[3531]),
			.NE(gen[3532]),

			.O(gen[3590]),
			.E(gen[3592]),

			.SO(gen[3530]),
			.S(gen[3531]),
			.SE(gen[3532]),

			.SELF(gen[3591]),
			.cell_state(gen[3591])
		); 

/******************* CELL 3592 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3592 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3531]),
			.N(gen[3532]),
			.NE(gen[3533]),

			.O(gen[3591]),
			.E(gen[3593]),

			.SO(gen[3531]),
			.S(gen[3532]),
			.SE(gen[3533]),

			.SELF(gen[3592]),
			.cell_state(gen[3592])
		); 

/******************* CELL 3593 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3593 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3532]),
			.N(gen[3533]),
			.NE(gen[3534]),

			.O(gen[3592]),
			.E(gen[3594]),

			.SO(gen[3532]),
			.S(gen[3533]),
			.SE(gen[3534]),

			.SELF(gen[3593]),
			.cell_state(gen[3593])
		); 

/******************* CELL 3594 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3594 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3533]),
			.N(gen[3534]),
			.NE(gen[3535]),

			.O(gen[3593]),
			.E(gen[3595]),

			.SO(gen[3533]),
			.S(gen[3534]),
			.SE(gen[3535]),

			.SELF(gen[3594]),
			.cell_state(gen[3594])
		); 

/******************* CELL 3595 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3595 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3534]),
			.N(gen[3535]),
			.NE(gen[3536]),

			.O(gen[3594]),
			.E(gen[3596]),

			.SO(gen[3534]),
			.S(gen[3535]),
			.SE(gen[3536]),

			.SELF(gen[3595]),
			.cell_state(gen[3595])
		); 

/******************* CELL 3596 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3596 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3535]),
			.N(gen[3536]),
			.NE(gen[3537]),

			.O(gen[3595]),
			.E(gen[3597]),

			.SO(gen[3535]),
			.S(gen[3536]),
			.SE(gen[3537]),

			.SELF(gen[3596]),
			.cell_state(gen[3596])
		); 

/******************* CELL 3597 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3597 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3536]),
			.N(gen[3537]),
			.NE(gen[3538]),

			.O(gen[3596]),
			.E(gen[3598]),

			.SO(gen[3536]),
			.S(gen[3537]),
			.SE(gen[3538]),

			.SELF(gen[3597]),
			.cell_state(gen[3597])
		); 

/******************* CELL 3598 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3598 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3537]),
			.N(gen[3538]),
			.NE(gen[3539]),

			.O(gen[3597]),
			.E(gen[3599]),

			.SO(gen[3537]),
			.S(gen[3538]),
			.SE(gen[3539]),

			.SELF(gen[3598]),
			.cell_state(gen[3598])
		); 

/******************* CELL 3599 ***************/  

	CELDA   #(.ic(0), .top_row(0), .bottom_row(1))

		cell3599 (
 			.clk(clk),
			.reset(reset),

			.operation(operation),

			.NO(gen[3538]),
			.N(gen[3539]),
			.NE(gen[3538]),

			.O(gen[3598]),
			.E(gen[3598]),

			.SO(gen[3538]),
			.S(gen[3539]),
			.SE(gen[3538]),

			.SELF(gen[3599]),
			.cell_state(gen[3599])
		); 



 assign data_out = {7'b0, gen[3599]};

endmodule